library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity LEDCUBE_8_8_8 is
	port (CLK : in std_logic;
			RST : in std_logic;
			SW1 : in std_logic;
			SW2 : in std_logic;
			SW3 : in std_logic;
			SW4 : in std_logic;
			SW5 : in std_logic;
			SW6 : in std_logic;
			SW7 : in std_logic;
			SW8 : in std_logic;
			SW9 : in std_logic;
			LED : out std_logic_vector(63 downto 0));
end LEDCUBE_8_8_8;

architecture Behavioral of LEDCUBE_8_8_8 is
	signal cnt23 : std_logic_vector(21 downto 0);
	signal cnt4 : std_logic_vector(3 downto 0);
	signal cnt7 : std_logic_vector(6 downto 0);
	

begin

process(CLK)
begin
	if(CLK'event and CLK='1')then
		if(RST='0')then
			cnt23 <= "0000000000000000000000";
		else
			cnt23 <= cnt23 + '1';
		end if;
	end if;
end process;

process(CLK)
begin
	if(CLK' event and CLK='1')then
		if(RST='0')then
			cnt4 <= "1111";
			cnt7 <= "0000000";
		elsif(cnt23="1111111111111111111111")then
			if(cnt4="1101")then
				cnt4 <= "0000";
			elsif(cnt7="1101111")then
				cnt7 <= "0000000";
			else
				cnt4 <= cnt4 + '1';
				cnt7 <= cnt7 + '1';
			end if;
		end if;
	end if;
end process;

process(cnt4,cnt7,SW1,SW2,SW3)
begin
	if(SW1='1' and SW2='0' and SW3='0' and SW4='0' and SW5='0' and SW6='0' and SW7='0' and SW8='0' and SW9='0')then
		case cnt4 is
			when "0000" => LED <= "0000000000000000000000000000000000000000000000000000000011111111";
			when "0001" => LED <= "0000000000000000000000000000000000000000000000001111111100000000";
			when "0010" => LED <= "0000000000000000000000000000000000000000111111110000000000000000";
			when "0011" => LED <= "0000000000000000000000000000000011111111000000000000000000000000";
			when "0100" => LED <= "0000000000000000000000001111111100000000000000000000000000000000";
			when "0101" => LED <= "0000000000000000111111110000000000000000000000000000000000000000";
			when "0110" => LED <= "0000000011111111000000000000000000000000000000000000000000000000";
			when "0111" => LED <= "1111111100000000000000000000000000000000000000000000000000000000";
			when "1000" => LED <= "0000000011111111000000000000000000000000000000000000000000000000";
			when "1001" => LED <= "0000000000000000111111110000000000000000000000000000000000000000";
			when "1010" => LED <= "0000000000000000000000001111111100000000000000000000000000000000";
			when "1011" => LED <= "0000000000000000000000000000000011111111000000000000000000000000";
			when "1100" => LED <= "0000000000000000000000000000000000000000111111110000000000000000";
			when "1101" => LED <= "0000000000000000000000000000000000000000000000001111111100000000";
			
			when "1111" => LED <= "0000000000000000000000000000000000000000000000000000000000000000";
			when others => null;
		end case;
		
	elsif(SW1='0' and SW2='1' and SW3='0' and SW4='0' and SW5='0' and SW6='0' and SW7='0' and SW8='0' and SW9='0')then
		case cnt4 is
			when "0000" => LED <= "0000000000000000000000000000000000000000000000000000000011111111";
			when "0001" => LED <= "0000000000000000000000000000000000000000000000001111111111111111";
			when "0010" => LED <= "0000000000000000000000000000000000000000111111111111111111111111";
			when "0011" => LED <= "0000000000000000000000000000000011111111111111111111111111111111";
			when "0100" => LED <= "0000000000000000000000001111111111111111111111111111111111111111";
			when "0101" => LED <= "0000000000000000111111111111111111111111111111111111111111111111";
			when "0110" => LED <= "0000000011111111111111111111111111111111111111111111111111111111";
			when "0111" => LED <= "1111111111111111111111111111111111111111111111111111111111111111";
			when "1000" => LED <= "0000000011111111111111111111111111111111111111111111111111111111";
			when "1001" => LED <= "0000000000000000111111111111111111111111111111111111111111111111";
			when "1010" => LED <= "0000000000000000000000001111111111111111111111111111111111111111";
			when "1011" => LED <= "0000000000000000000000000000000011111111111111111111111111111111";
			when "1100" => LED <= "0000000000000000000000000000000000000000111111111111111111111111";
			when "1101" => LED <= "0000000000000000000000000000000000000000000000001111111111111111";
			
			when "1111" => LED <= "0000000000000000000000000000000000000000000000000000000000000000";
			when others => null;
		end case;
		
		
	elsif(SW1='0' and SW2='0' and SW3='1' and SW4='0' and SW5='0' and SW6='0' and SW7='0' and SW8='0' and SW9='0')then
		case cnt4 is
			when "0000" => LED <= "0000000100000001000000010000000100000001000000010000000100000001";
			when "0001" => LED <= "0000001000000010000000100000001000000010000000100000001000000010";
			when "0010" => LED <= "0000010000000100000001000000010000000100000001000000010000000100";
			when "0011" => LED <= "0000100000001000000010000000100000001000000010000000100000001000";
			when "0100" => LED <= "0001000000010000000100000001000000010000000100000001000000010000";
			when "0101" => LED <= "0010000000100000001000000010000000100000001000000010000000100000";
			when "0110" => LED <= "0100000001000000010000000100000001000000010000000100000001000000";
			when "0111" => LED <= "1000000010000000100000001000000010000000100000001000000010000000";
			when "1000" => LED <= "0100000001000000010000000100000001000000010000000100000001000000";
			when "1001" => LED <= "0010000000100000001000000010000000100000001000000010000000100000";
			when "1010" => LED <= "0001000000010000000100000001000000010000000100000001000000010000";
			when "1011" => LED <= "0000100000001000000010000000100000001000000010000000100000001000";
			when "1100" => LED <= "0000010000000100000001000000010000000100000001000000010000000100";
			when "1101" => LED <= "0000001000000010000000100000001000000010000000100000001000000010";
			
			when "1111" => LED <= "0000000000000000000000000000000000000000000000000000000000000000";
			when others => null;
		end case;
		
	elsif(SW1='0' and SW2='0' and SW3='0' and SW4='1' and SW5='0' and SW6='0' and SW7='0' and SW8='0' and SW9='0')then
		case cnt4 is
			when "0000" => LED <= "0000000100000001000000010000000100000001000000010000000100000001";
			when "0001" => LED <= "0000001100000011000000110000001100000011000000110000001100000011";
			when "0010" => LED <= "0000011100000111000001110000011100000111000001110000011100000111";
			when "0011" => LED <= "0000111100001111000011110000111100001111000011110000111100001111";
			when "0100" => LED <= "0001111100011111000111110001111100011111000111110001111100011111";
			when "0101" => LED <= "0011111100111111001111110011111100111111001111110011111100111111";
			when "0110" => LED <= "0111111101111111011111110111111101111111011111110111111101111111";
			when "0111" => LED <= "1111111111111111111111111111111111111111111111111111111111111111";
			when "1000" => LED <= "0111111101111111011111110111111101111111011111110111111101111111";
			when "1001" => LED <= "0011111100111111001111110011111100111111001111110011111100111111";
			when "1010" => LED <= "0001111100011111000111110001111100011111000111110001111100011111";
			when "1011" => LED <= "0000111100001111000011110000111100001111000011110000111100001111";
			when "1100" => LED <= "0000011100000111000001110000011100000111000001110000011100000111";
			when "1101" => LED <= "0000001100000011000000110000001100000011000000110000001100000011";
			
			when "1111" => LED <= "0000000000000000000000000000000000000000000000000000000000000000";
			when others => null;
		end case;
		
		
	elsif(SW1='0' and SW2='0' and SW3='0' and SW4='0' and SW5='0' and SW6='1' and SW7='0' and SW8='0' and SW9='0')then
		case cnt4 is
			when "0000" => LED <= "0000000000000000000000000001100000011000000000000000000000000000";
			when "0001" => LED <= "0000000000000000001111000011110000111100001111000000000000000000";
			when "0010" => LED <= "0000000001111110011111100111111001111110011111100111111000000000";
			when "0011" => LED <= "1111111111111111111111111111111111111111111111111111111111111111";
			when "0100" => LED <= "0000000001111110011111100111111001111110011111100111111000000000";
			when "0101" => LED <= "0000000000000000001111000011110000111100001111000000000000000000";
			when "0110" => LED <= "0000000000000000000000000001100000011000000000000000000000000000";
			when "0111" => LED <= "0000000000000000001111000011110000111100001111000000000000000000";
			when "1000" => LED <= "0000000001111110011111100111111001111110011111100111111000000000";
			when "1001" => LED <= "1111111111111111111111111111111111111111111111111111111111111111";
			when "1010" => LED <= "0000000001111110011111100111111001111110011111100111111000000000";
			when "1011" => LED <= "0000000000000000001111000011110000111100001111000000000000000000";
			when "1100" => LED <= "0000000000000000000000000001100000011000000000000000000000000000";
			when "1101" => LED <= "0000000000000000000000000001100000011000000000000000000000000000";
			
			when "1111" => LED <= "0000000000000000000000000000000000000000000000000000000000000000";
			when others => null;
		end case;
		
		
	elsif(SW1='0' and SW2='0' and SW3='0' and SW4='0' and SW5='1' and SW6='0' and SW7='0' and SW8='0' and SW9='0')then
		case cnt4 is
			when "0000" => LED <= "0000000000000000000000000001100000011000000000000000000000000000";
			when "0001" => LED <= "0000000000000000001111000010010000100100001111000000000000000000";
			when "0010" => LED <= "0000000001111110010000100100001001000010010000100111111000000000";
			when "0011" => LED <= "1111111110000001100000011000000110000001100000011000000111111111";
			when "0100" => LED <= "0000000001111110010000100100001001000010010000100111111000000000";
			when "0101" => LED <= "0000000000000000001111000010010000100100001111000000000000000000";
			when "0110" => LED <= "0000000000000000000000000001100000011000000000000000000000000000";
			when "0111" => LED <= "0000000000000000001111000010010000100100001111000000000000000000";
			when "1000" => LED <= "0000000001111110010000100100001001000010010000100111111000000000";
			when "1001" => LED <= "1111111110000001100000011000000110000001100000011000000111111111";
			when "1010" => LED <= "0000000001111110010000100100001001000010010000100111111000000000";
			when "1011" => LED <= "0000000000000000001111000010010000100100001111000000000000000000";
			when "1100" => LED <= "0000000000000000000000000001100000011000000000000000000000000000";
			when "1101" => LED <= "0000000000000000000000000001100000011000000000000000000000000000";
			
			when "1111" => LED <= "0000000000000000000000000000000000000000000000000000000000000000";
			when others => null;
		end case;
		
		
	elsif(SW1='0' and SW2='0' and SW3='0' and SW4='0' and SW5='0' and SW6='0' and SW7='1' and SW8='0' and SW9='0')then
		case cnt4 is
			when "0000" => LED <= "1111111100000000000000000000000000000000000000000000000011111111";
			when "0001" => LED <= "0000000011111111000000000000000000000000000000001111111100000000";
			when "0010" => LED <= "0000000000000000111111110000000000000000111111110000000000000000";
			when "0011" => LED <= "0000000000000000000000001111111111111111000000000000000000000000";
			when "0100" => LED <= "0000000000000000000000001111111111111111000000000000000000000000";
			when "0101" => LED <= "0000000000000000111111110000000000000000111111110000000000000000";
			when "0110" => LED <= "0000000011111111000000000000000000000000000000001111111100000000";
			when "0111" => LED <= "1111111100000000000000000000000000000000000000000000000011111111";
			when "1000" => LED <= "0000000011111111000000000000000000000000000000001111111100000000";
			when "1001" => LED <= "0000000000000000111111110000000000000000111111110000000000000000";
			when "1010" => LED <= "0000000000000000000000001111111111111111000000000000000000000000";
			when "1011" => LED <= "0000000000000000000000001111111111111111000000000000000000000000";
			when "1100" => LED <= "0000000000000000111111110000000000000000111111110000000000000000";
			when "1101" => LED <= "0000000011111111000000000000000000000000000000001111111100000000";
			
			when "1111" => LED <= "0000000000000000000000000000000000000000000000000000000000000000";
			when others => null;
		end case;
	
	
	elsif(SW1='0' and SW2='0' and SW3='0' and SW4='0' and SW5='0' and SW6='0' and SW7='0' and SW8='1' and SW9='0')then
		case cnt4 is
			when "0000" => LED <= "1000000110000001100000011000000110000001100000011000000110000001";
			when "0001" => LED <= "0100001001000010010000100100001001000010010000100100001001000010";
			when "0010" => LED <= "0010010000100100001001000010010000100100001001000010010000100100";
			when "0011" => LED <= "0001100000011000000110000001100000011000000110000001100000011000";
			when "0100" => LED <= "0001100000011000000110000001100000011000000110000001100000011000";
			when "0101" => LED <= "0010010000100100001001000010010000100100001001000010010000100100";
			when "0110" => LED <= "0100001001000010010000100100001001000010010000100100001001000010";
			when "0111" => LED <= "1000000110000001100000011000000110000001100000011000000110000001";
			when "1000" => LED <= "0100001001000010010000100100001001000010010000100100001001000010";
			when "1001" => LED <= "0010010000100100001001000010010000100100001001000010010000100100";
			when "1010" => LED <= "0001100000011000000110000001100000011000000110000001100000011000";
			when "1011" => LED <= "0001100000011000000110000001100000011000000110000001100000011000";
			when "1100" => LED <= "0010010000100100001001000010010000100100001001000010010000100100";
			when "1101" => LED <= "0100001001000010010000100100001001000010010000100100001001000010";
			
			when "1111" => LED <= "0000000000000000000000000000000000000000000000000000000000000000";
			when others => null;
		end case;
	
	
	elsif(SW1='0' and SW2='0' and SW3='0' and SW4='0' and SW5='0' and SW6='0' and SW7='0' and SW8='0' and SW9='1')then
		case cnt7 is
			when "0000000" => LED <= "0000000000000000000000000000000000000000000000000000000011111111";
			when "0000001" => LED <= "0000000000000000000000000000000000000000000000001111111100000000";
			when "0000010" => LED <= "0000000000000000000000000000000000000000111111110000000000000000";
			when "0000011" => LED <= "0000000000000000000000000000000011111111000000000000000000000000";
			when "0000100" => LED <= "0000000000000000000000001111111100000000000000000000000000000000";
			when "0000101" => LED <= "0000000000000000111111110000000000000000000000000000000000000000";
			when "0000110" => LED <= "0000000011111111000000000000000000000000000000000000000000000000";
			when "0000111" => LED <= "1111111100000000000000000000000000000000000000000000000000000000";
			when "0001000" => LED <= "0000000011111111000000000000000000000000000000000000000000000000";
			when "0001001" => LED <= "0000000000000000111111110000000000000000000000000000000000000000";
			when "0001010" => LED <= "0000000000000000000000001111111100000000000000000000000000000000";
			when "0001011" => LED <= "0000000000000000000000000000000011111111000000000000000000000000";
			when "0001100" => LED <= "0000000000000000000000000000000000000000111111110000000000000000";
			when "0001101" => LED <= "0000000000000000000000000000000000000000000000001111111100000000";
			
			when "0001110" => LED <= "0000000000000000000000000000000000000000000000000000000011111111";
			when "0001111" => LED <= "0000000000000000000000000000000000000000000000001111111111111111";
			when "0010000" => LED <= "0000000000000000000000000000000000000000111111111111111111111111";
			when "0010001" => LED <= "0000000000000000000000000000000011111111111111111111111111111111";
			when "0010010" => LED <= "0000000000000000000000001111111111111111111111111111111111111111";
			when "0010011" => LED <= "0000000000000000111111111111111111111111111111111111111111111111";
			when "0010100" => LED <= "0000000011111111111111111111111111111111111111111111111111111111";
			when "0010101" => LED <= "1111111111111111111111111111111111111111111111111111111111111111";
			when "0010110" => LED <= "0000000011111111111111111111111111111111111111111111111111111111";
			when "0010111" => LED <= "0000000000000000111111111111111111111111111111111111111111111111";
			when "0011000" => LED <= "0000000000000000000000001111111111111111111111111111111111111111";
			when "0011001" => LED <= "0000000000000000000000000000000011111111111111111111111111111111";
			when "0011010" => LED <= "0000000000000000000000000000000000000000111111111111111111111111";
			when "0011011" => LED <= "0000000000000000000000000000000000000000000000001111111111111111";
			
			when "0011100" => LED <= "0000000100000001000000010000000100000001000000010000000100000001";
			when "0011101" => LED <= "0000001000000010000000100000001000000010000000100000001000000010";
			when "0011110" => LED <= "0000010000000100000001000000010000000100000001000000010000000100";
			when "0011111" => LED <= "0000100000001000000010000000100000001000000010000000100000001000";
			when "0100000" => LED <= "0001000000010000000100000001000000010000000100000001000000010000";
			when "0100001" => LED <= "0010000000100000001000000010000000100000001000000010000000100000";
			when "0100010" => LED <= "0100000001000000010000000100000001000000010000000100000001000000";
			when "0100011" => LED <= "1000000010000000100000001000000010000000100000001000000010000000";
			when "0100100" => LED <= "0100000001000000010000000100000001000000010000000100000001000000";
			when "0100101" => LED <= "0010000000100000001000000010000000100000001000000010000000100000";
			when "0100110" => LED <= "0001000000010000000100000001000000010000000100000001000000010000";
			when "0100111" => LED <= "0000100000001000000010000000100000001000000010000000100000001000";
			when "0101000" => LED <= "0000010000000100000001000000010000000100000001000000010000000100";
			when "0101001" => LED <= "0000001000000010000000100000001000000010000000100000001000000010";
			
			when "0101010" => LED <= "0000000100000001000000010000000100000001000000010000000100000001";
			when "0101011" => LED <= "0000001100000011000000110000001100000011000000110000001100000011";
			when "0101100" => LED <= "0000011100000111000001110000011100000111000001110000011100000111";
			when "0101101" => LED <= "0000111100001111000011110000111100001111000011110000111100001111";
			when "0101110" => LED <= "0001111100011111000111110001111100011111000111110001111100011111";
			when "0101111" => LED <= "0011111100111111001111110011111100111111001111110011111100111111";
			when "0110000" => LED <= "0111111101111111011111110111111101111111011111110111111101111111";
			when "0110001" => LED <= "1111111111111111111111111111111111111111111111111111111111111111";
			when "0110010" => LED <= "0111111101111111011111110111111101111111011111110111111101111111";
			when "0110011" => LED <= "0011111100111111001111110011111100111111001111110011111100111111";
			when "0110100" => LED <= "0001111100011111000111110001111100011111000111110001111100011111";
			when "0110101" => LED <= "0000111100001111000011110000111100001111000011110000111100001111";
			when "0110110" => LED <= "0000011100000111000001110000011100000111000001110000011100000111";
			when "0110111" => LED <= "0000001100000011000000110000001100000011000000110000001100000011";
			
			when "0111000" => LED <= "0000000000000000000000000001100000011000000000000000000000000000";
			when "0111001" => LED <= "0000000000000000001111000010010000100100001111000000000000000000";
			when "0111010" => LED <= "0000000001111110010000100100001001000010010000100111111000000000";
			when "0111011" => LED <= "1111111110000001100000011000000110000001100000011000000111111111";
			when "0111100" => LED <= "0000000001111110010000100100001001000010010000100111111000000000";
			when "0111101" => LED <= "0000000000000000001111000010010000100100001111000000000000000000";
			when "0111110" => LED <= "0000000000000000000000000001100000011000000000000000000000000000";
			when "0111111" => LED <= "0000000000000000001111000010010000100100001111000000000000000000";
			when "1000000" => LED <= "0000000001111110010000100100001001000010010000100111111000000000";
			when "1000001" => LED <= "1111111110000001100000011000000110000001100000011000000111111111";
			when "1000010" => LED <= "0000000001111110010000100100001001000010010000100111111000000000";
			when "1000011" => LED <= "0000000000000000001111000010010000100100001111000000000000000000";
			when "1000100" => LED <= "0000000000000000000000000001100000011000000000000000000000000000";
			when "1000101" => LED <= "0000000000000000000000000001100000011000000000000000000000000000";
			
			when "1000110" => LED <= "0000000000000000000000000001100000011000000000000000000000000000";
			when "1000111" => LED <= "0000000000000000001111000011110000111100001111000000000000000000";
			when "1001000" => LED <= "0000000001111110011111100111111001111110011111100111111000000000";
			when "1001001" => LED <= "1111111111111111111111111111111111111111111111111111111111111111";
			when "1001010" => LED <= "0000000001111110011111100111111001111110011111100111111000000000";
			when "1001011" => LED <= "0000000000000000001111000011110000111100001111000000000000000000";
			when "1001100" => LED <= "0000000000000000000000000001100000011000000000000000000000000000";
			when "1001101" => LED <= "0000000000000000001111000011110000111100001111000000000000000000";
			when "1001110" => LED <= "0000000001111110011111100111111001111110011111100111111000000000";
			when "1001111" => LED <= "1111111111111111111111111111111111111111111111111111111111111111";
			when "1010000" => LED <= "0000000001111110011111100111111001111110011111100111111000000000";
			when "1010001" => LED <= "0000000000000000001111000011110000111100001111000000000000000000";
			when "1010010" => LED <= "0000000000000000000000000001100000011000000000000000000000000000";
			when "1010011" => LED <= "0000000000000000000000000001100000011000000000000000000000000000";
			
			when "1010100" => LED <= "1111111100000000000000000000000000000000000000000000000011111111";
			when "1010101" => LED <= "0000000011111111000000000000000000000000000000001111111100000000";
			when "1010110" => LED <= "0000000000000000111111110000000000000000111111110000000000000000";
			when "1010111" => LED <= "0000000000000000000000001111111111111111000000000000000000000000";
			when "1011000" => LED <= "0000000000000000000000001111111111111111000000000000000000000000";
			when "1011001" => LED <= "0000000000000000111111110000000000000000111111110000000000000000";
			when "1011010" => LED <= "0000000011111111000000000000000000000000000000001111111100000000";
			when "1011011" => LED <= "1111111100000000000000000000000000000000000000000000000011111111";
			when "1011100" => LED <= "0000000011111111000000000000000000000000000000001111111100000000";
			when "1011101" => LED <= "0000000000000000111111110000000000000000111111110000000000000000";
			when "1011110" => LED <= "0000000000000000000000001111111111111111000000000000000000000000";
			when "1011111" => LED <= "0000000000000000000000001111111111111111000000000000000000000000";
			when "1100000" => LED <= "0000000000000000111111110000000000000000111111110000000000000000";
			when "1100001" => LED <= "0000000011111111000000000000000000000000000000001111111100000000";
			
			when "1100010" => LED <= "1000000110000001100000011000000110000001100000011000000110000001";
			when "1100011" => LED <= "0100001001000010010000100100001001000010010000100100001001000010";
			when "1100100" => LED <= "0010010000100100001001000010010000100100001001000010010000100100";
			when "1100101" => LED <= "0001100000011000000110000001100000011000000110000001100000011000";
			when "1100110" => LED <= "0001100000011000000110000001100000011000000110000001100000011000";
			when "1100111" => LED <= "0010010000100100001001000010010000100100001001000010010000100100";
			when "1101000" => LED <= "0100001001000010010000100100001001000010010000100100001001000010";
			when "1101001" => LED <= "1000000110000001100000011000000110000001100000011000000110000001";
			when "1101010" => LED <= "0100001001000010010000100100001001000010010000100100001001000010";
			when "1101011" => LED <= "0010010000100100001001000010010000100100001001000010010000100100";
			when "1101100" => LED <= "0001100000011000000110000001100000011000000110000001100000011000";
			when "1101101" => LED <= "0001100000011000000110000001100000011000000110000001100000011000";
			when "1101110" => LED <= "0010010000100100001001000010010000100100001001000010010000100100";
			when "1101111" => LED <= "0100001001000010010000100100001001000010010000100100001001000010";
			
			when "1111111" => LED <= "0000000000000000000000000000000000000000000000000000000000000000";
			when others => null;
		end case;
	
	else
		LED <= "0000000000000000000000000000000000000000000000000000000000000000";
	end if;
end process;

end Behavioral;