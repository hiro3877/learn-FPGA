`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/08/20 20:43:41
// Design Name: 
// Module Name: top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
/////////////////////////////////////////////////////////////////////////////////

`include "./nettype.h"
`include "./std_define.h"

module top_io(
input wire clk,
input wire signed [`InBus]		in_r,
input wire signed [`InBus]		in_i,
output wire signed [`OutBus]		out_r,
output wire signed [`OutBus]		out_i

);

wire signed [`InBus]		in_1_1_r;
wire signed [`InBus]		in_1_1_i;
wire signed [`InBus]		in_1_2_r;
wire signed [`InBus]		in_1_2_i;
wire signed [`InBus]		in_1_3_r;
wire signed [`InBus]		in_1_3_i;
wire signed [`InBus]		in_1_4_r;
wire signed [`InBus]		in_1_4_i;
wire signed [`InBus]		in_1_5_r;
wire signed [`InBus]		in_1_5_i;
wire signed [`InBus]		in_1_6_r;
wire signed [`InBus]		in_1_6_i;
wire signed [`InBus]		in_1_7_r;
wire signed [`InBus]		in_1_7_i;
wire signed [`InBus]		in_1_8_r;
wire signed [`InBus]		in_1_8_i;
wire signed [`InBus]		in_1_9_r;
wire signed [`InBus]		in_1_9_i;
wire signed [`InBus]		in_1_10_r;
wire signed [`InBus]		in_1_10_i;
wire signed [`InBus]		in_1_11_r;
wire signed [`InBus]		in_1_11_i;
wire signed [`InBus]		in_1_12_r;
wire signed [`InBus]		in_1_12_i;
wire signed [`InBus]		in_1_13_r;
wire signed [`InBus]		in_1_13_i;
wire signed [`InBus]		in_1_14_r;
wire signed [`InBus]		in_1_14_i;
wire signed [`InBus]		in_1_15_r;
wire signed [`InBus]		in_1_15_i;
wire signed [`InBus]		in_1_16_r;
wire signed [`InBus]		in_1_16_i;
wire signed [`InBus]		in_1_17_r;
wire signed [`InBus]		in_1_17_i;
wire signed [`InBus]		in_1_18_r;
wire signed [`InBus]		in_1_18_i;
wire signed [`InBus]		in_1_19_r;
wire signed [`InBus]		in_1_19_i;
wire signed [`InBus]		in_1_20_r;
wire signed [`InBus]		in_1_20_i;
wire signed [`InBus]		in_1_21_r;
wire signed [`InBus]		in_1_21_i;
wire signed [`InBus]		in_1_22_r;
wire signed [`InBus]		in_1_22_i;
wire signed [`InBus]		in_1_23_r;
wire signed [`InBus]		in_1_23_i;
wire signed [`InBus]		in_1_24_r;
wire signed [`InBus]		in_1_24_i;
wire signed [`InBus]		in_1_25_r;
wire signed [`InBus]		in_1_25_i;
wire signed [`InBus]		in_1_26_r;
wire signed [`InBus]		in_1_26_i;
wire signed [`InBus]		in_1_27_r;
wire signed [`InBus]		in_1_27_i;
wire signed [`InBus]		in_1_28_r;
wire signed [`InBus]		in_1_28_i;
wire signed [`InBus]		in_1_29_r;
wire signed [`InBus]		in_1_29_i;
wire signed [`InBus]		in_1_30_r;
wire signed [`InBus]		in_1_30_i;
wire signed [`InBus]		in_1_31_r;
wire signed [`InBus]		in_1_31_i;
wire signed [`InBus]		in_1_32_r;
wire signed [`InBus]		in_1_32_i;
wire signed [`InBus]		in_2_1_r;
wire signed [`InBus]		in_2_1_i;
wire signed [`InBus]		in_2_2_r;
wire signed [`InBus]		in_2_2_i;
wire signed [`InBus]		in_2_3_r;
wire signed [`InBus]		in_2_3_i;
wire signed [`InBus]		in_2_4_r;
wire signed [`InBus]		in_2_4_i;
wire signed [`InBus]		in_2_5_r;
wire signed [`InBus]		in_2_5_i;
wire signed [`InBus]		in_2_6_r;
wire signed [`InBus]		in_2_6_i;
wire signed [`InBus]		in_2_7_r;
wire signed [`InBus]		in_2_7_i;
wire signed [`InBus]		in_2_8_r;
wire signed [`InBus]		in_2_8_i;
wire signed [`InBus]		in_2_9_r;
wire signed [`InBus]		in_2_9_i;
wire signed [`InBus]		in_2_10_r;
wire signed [`InBus]		in_2_10_i;
wire signed [`InBus]		in_2_11_r;
wire signed [`InBus]		in_2_11_i;
wire signed [`InBus]		in_2_12_r;
wire signed [`InBus]		in_2_12_i;
wire signed [`InBus]		in_2_13_r;
wire signed [`InBus]		in_2_13_i;
wire signed [`InBus]		in_2_14_r;
wire signed [`InBus]		in_2_14_i;
wire signed [`InBus]		in_2_15_r;
wire signed [`InBus]		in_2_15_i;
wire signed [`InBus]		in_2_16_r;
wire signed [`InBus]		in_2_16_i;
wire signed [`InBus]		in_2_17_r;
wire signed [`InBus]		in_2_17_i;
wire signed [`InBus]		in_2_18_r;
wire signed [`InBus]		in_2_18_i;
wire signed [`InBus]		in_2_19_r;
wire signed [`InBus]		in_2_19_i;
wire signed [`InBus]		in_2_20_r;
wire signed [`InBus]		in_2_20_i;
wire signed [`InBus]		in_2_21_r;
wire signed [`InBus]		in_2_21_i;
wire signed [`InBus]		in_2_22_r;
wire signed [`InBus]		in_2_22_i;
wire signed [`InBus]		in_2_23_r;
wire signed [`InBus]		in_2_23_i;
wire signed [`InBus]		in_2_24_r;
wire signed [`InBus]		in_2_24_i;
wire signed [`InBus]		in_2_25_r;
wire signed [`InBus]		in_2_25_i;
wire signed [`InBus]		in_2_26_r;
wire signed [`InBus]		in_2_26_i;
wire signed [`InBus]		in_2_27_r;
wire signed [`InBus]		in_2_27_i;
wire signed [`InBus]		in_2_28_r;
wire signed [`InBus]		in_2_28_i;
wire signed [`InBus]		in_2_29_r;
wire signed [`InBus]		in_2_29_i;
wire signed [`InBus]		in_2_30_r;
wire signed [`InBus]		in_2_30_i;
wire signed [`InBus]		in_2_31_r;
wire signed [`InBus]		in_2_31_i;
wire signed [`InBus]		in_2_32_r;
wire signed [`InBus]		in_2_32_i;
wire signed [`InBus]		in_3_1_r;
wire signed [`InBus]		in_3_1_i;
wire signed [`InBus]		in_3_2_r;
wire signed [`InBus]		in_3_2_i;
wire signed [`InBus]		in_3_3_r;
wire signed [`InBus]		in_3_3_i;
wire signed [`InBus]		in_3_4_r;
wire signed [`InBus]		in_3_4_i;
wire signed [`InBus]		in_3_5_r;
wire signed [`InBus]		in_3_5_i;
wire signed [`InBus]		in_3_6_r;
wire signed [`InBus]		in_3_6_i;
wire signed [`InBus]		in_3_7_r;
wire signed [`InBus]		in_3_7_i;
wire signed [`InBus]		in_3_8_r;
wire signed [`InBus]		in_3_8_i;
wire signed [`InBus]		in_3_9_r;
wire signed [`InBus]		in_3_9_i;
wire signed [`InBus]		in_3_10_r;
wire signed [`InBus]		in_3_10_i;
wire signed [`InBus]		in_3_11_r;
wire signed [`InBus]		in_3_11_i;
wire signed [`InBus]		in_3_12_r;
wire signed [`InBus]		in_3_12_i;
wire signed [`InBus]		in_3_13_r;
wire signed [`InBus]		in_3_13_i;
wire signed [`InBus]		in_3_14_r;
wire signed [`InBus]		in_3_14_i;
wire signed [`InBus]		in_3_15_r;
wire signed [`InBus]		in_3_15_i;
wire signed [`InBus]		in_3_16_r;
wire signed [`InBus]		in_3_16_i;
wire signed [`InBus]		in_3_17_r;
wire signed [`InBus]		in_3_17_i;
wire signed [`InBus]		in_3_18_r;
wire signed [`InBus]		in_3_18_i;
wire signed [`InBus]		in_3_19_r;
wire signed [`InBus]		in_3_19_i;
wire signed [`InBus]		in_3_20_r;
wire signed [`InBus]		in_3_20_i;
wire signed [`InBus]		in_3_21_r;
wire signed [`InBus]		in_3_21_i;
wire signed [`InBus]		in_3_22_r;
wire signed [`InBus]		in_3_22_i;
wire signed [`InBus]		in_3_23_r;
wire signed [`InBus]		in_3_23_i;
wire signed [`InBus]		in_3_24_r;
wire signed [`InBus]		in_3_24_i;
wire signed [`InBus]		in_3_25_r;
wire signed [`InBus]		in_3_25_i;
wire signed [`InBus]		in_3_26_r;
wire signed [`InBus]		in_3_26_i;
wire signed [`InBus]		in_3_27_r;
wire signed [`InBus]		in_3_27_i;
wire signed [`InBus]		in_3_28_r;
wire signed [`InBus]		in_3_28_i;
wire signed [`InBus]		in_3_29_r;
wire signed [`InBus]		in_3_29_i;
wire signed [`InBus]		in_3_30_r;
wire signed [`InBus]		in_3_30_i;
wire signed [`InBus]		in_3_31_r;
wire signed [`InBus]		in_3_31_i;
wire signed [`InBus]		in_3_32_r;
wire signed [`InBus]		in_3_32_i;
wire signed [`InBus]		in_4_1_r;
wire signed [`InBus]		in_4_1_i;
wire signed [`InBus]		in_4_2_r;
wire signed [`InBus]		in_4_2_i;
wire signed [`InBus]		in_4_3_r;
wire signed [`InBus]		in_4_3_i;
wire signed [`InBus]		in_4_4_r;
wire signed [`InBus]		in_4_4_i;
wire signed [`InBus]		in_4_5_r;
wire signed [`InBus]		in_4_5_i;
wire signed [`InBus]		in_4_6_r;
wire signed [`InBus]		in_4_6_i;
wire signed [`InBus]		in_4_7_r;
wire signed [`InBus]		in_4_7_i;
wire signed [`InBus]		in_4_8_r;
wire signed [`InBus]		in_4_8_i;
wire signed [`InBus]		in_4_9_r;
wire signed [`InBus]		in_4_9_i;
wire signed [`InBus]		in_4_10_r;
wire signed [`InBus]		in_4_10_i;
wire signed [`InBus]		in_4_11_r;
wire signed [`InBus]		in_4_11_i;
wire signed [`InBus]		in_4_12_r;
wire signed [`InBus]		in_4_12_i;
wire signed [`InBus]		in_4_13_r;
wire signed [`InBus]		in_4_13_i;
wire signed [`InBus]		in_4_14_r;
wire signed [`InBus]		in_4_14_i;
wire signed [`InBus]		in_4_15_r;
wire signed [`InBus]		in_4_15_i;
wire signed [`InBus]		in_4_16_r;
wire signed [`InBus]		in_4_16_i;
wire signed [`InBus]		in_4_17_r;
wire signed [`InBus]		in_4_17_i;
wire signed [`InBus]		in_4_18_r;
wire signed [`InBus]		in_4_18_i;
wire signed [`InBus]		in_4_19_r;
wire signed [`InBus]		in_4_19_i;
wire signed [`InBus]		in_4_20_r;
wire signed [`InBus]		in_4_20_i;
wire signed [`InBus]		in_4_21_r;
wire signed [`InBus]		in_4_21_i;
wire signed [`InBus]		in_4_22_r;
wire signed [`InBus]		in_4_22_i;
wire signed [`InBus]		in_4_23_r;
wire signed [`InBus]		in_4_23_i;
wire signed [`InBus]		in_4_24_r;
wire signed [`InBus]		in_4_24_i;
wire signed [`InBus]		in_4_25_r;
wire signed [`InBus]		in_4_25_i;
wire signed [`InBus]		in_4_26_r;
wire signed [`InBus]		in_4_26_i;
wire signed [`InBus]		in_4_27_r;
wire signed [`InBus]		in_4_27_i;
wire signed [`InBus]		in_4_28_r;
wire signed [`InBus]		in_4_28_i;
wire signed [`InBus]		in_4_29_r;
wire signed [`InBus]		in_4_29_i;
wire signed [`InBus]		in_4_30_r;
wire signed [`InBus]		in_4_30_i;
wire signed [`InBus]		in_4_31_r;
wire signed [`InBus]		in_4_31_i;
wire signed [`InBus]		in_4_32_r;
wire signed [`InBus]		in_4_32_i;
wire signed [`InBus]		in_5_1_r;
wire signed [`InBus]		in_5_1_i;
wire signed [`InBus]		in_5_2_r;
wire signed [`InBus]		in_5_2_i;
wire signed [`InBus]		in_5_3_r;
wire signed [`InBus]		in_5_3_i;
wire signed [`InBus]		in_5_4_r;
wire signed [`InBus]		in_5_4_i;
wire signed [`InBus]		in_5_5_r;
wire signed [`InBus]		in_5_5_i;
wire signed [`InBus]		in_5_6_r;
wire signed [`InBus]		in_5_6_i;
wire signed [`InBus]		in_5_7_r;
wire signed [`InBus]		in_5_7_i;
wire signed [`InBus]		in_5_8_r;
wire signed [`InBus]		in_5_8_i;
wire signed [`InBus]		in_5_9_r;
wire signed [`InBus]		in_5_9_i;
wire signed [`InBus]		in_5_10_r;
wire signed [`InBus]		in_5_10_i;
wire signed [`InBus]		in_5_11_r;
wire signed [`InBus]		in_5_11_i;
wire signed [`InBus]		in_5_12_r;
wire signed [`InBus]		in_5_12_i;
wire signed [`InBus]		in_5_13_r;
wire signed [`InBus]		in_5_13_i;
wire signed [`InBus]		in_5_14_r;
wire signed [`InBus]		in_5_14_i;
wire signed [`InBus]		in_5_15_r;
wire signed [`InBus]		in_5_15_i;
wire signed [`InBus]		in_5_16_r;
wire signed [`InBus]		in_5_16_i;
wire signed [`InBus]		in_5_17_r;
wire signed [`InBus]		in_5_17_i;
wire signed [`InBus]		in_5_18_r;
wire signed [`InBus]		in_5_18_i;
wire signed [`InBus]		in_5_19_r;
wire signed [`InBus]		in_5_19_i;
wire signed [`InBus]		in_5_20_r;
wire signed [`InBus]		in_5_20_i;
wire signed [`InBus]		in_5_21_r;
wire signed [`InBus]		in_5_21_i;
wire signed [`InBus]		in_5_22_r;
wire signed [`InBus]		in_5_22_i;
wire signed [`InBus]		in_5_23_r;
wire signed [`InBus]		in_5_23_i;
wire signed [`InBus]		in_5_24_r;
wire signed [`InBus]		in_5_24_i;
wire signed [`InBus]		in_5_25_r;
wire signed [`InBus]		in_5_25_i;
wire signed [`InBus]		in_5_26_r;
wire signed [`InBus]		in_5_26_i;
wire signed [`InBus]		in_5_27_r;
wire signed [`InBus]		in_5_27_i;
wire signed [`InBus]		in_5_28_r;
wire signed [`InBus]		in_5_28_i;
wire signed [`InBus]		in_5_29_r;
wire signed [`InBus]		in_5_29_i;
wire signed [`InBus]		in_5_30_r;
wire signed [`InBus]		in_5_30_i;
wire signed [`InBus]		in_5_31_r;
wire signed [`InBus]		in_5_31_i;
wire signed [`InBus]		in_5_32_r;
wire signed [`InBus]		in_5_32_i;
wire signed [`InBus]		in_6_1_r;
wire signed [`InBus]		in_6_1_i;
wire signed [`InBus]		in_6_2_r;
wire signed [`InBus]		in_6_2_i;
wire signed [`InBus]		in_6_3_r;
wire signed [`InBus]		in_6_3_i;
wire signed [`InBus]		in_6_4_r;
wire signed [`InBus]		in_6_4_i;
wire signed [`InBus]		in_6_5_r;
wire signed [`InBus]		in_6_5_i;
wire signed [`InBus]		in_6_6_r;
wire signed [`InBus]		in_6_6_i;
wire signed [`InBus]		in_6_7_r;
wire signed [`InBus]		in_6_7_i;
wire signed [`InBus]		in_6_8_r;
wire signed [`InBus]		in_6_8_i;
wire signed [`InBus]		in_6_9_r;
wire signed [`InBus]		in_6_9_i;
wire signed [`InBus]		in_6_10_r;
wire signed [`InBus]		in_6_10_i;
wire signed [`InBus]		in_6_11_r;
wire signed [`InBus]		in_6_11_i;
wire signed [`InBus]		in_6_12_r;
wire signed [`InBus]		in_6_12_i;
wire signed [`InBus]		in_6_13_r;
wire signed [`InBus]		in_6_13_i;
wire signed [`InBus]		in_6_14_r;
wire signed [`InBus]		in_6_14_i;
wire signed [`InBus]		in_6_15_r;
wire signed [`InBus]		in_6_15_i;
wire signed [`InBus]		in_6_16_r;
wire signed [`InBus]		in_6_16_i;
wire signed [`InBus]		in_6_17_r;
wire signed [`InBus]		in_6_17_i;
wire signed [`InBus]		in_6_18_r;
wire signed [`InBus]		in_6_18_i;
wire signed [`InBus]		in_6_19_r;
wire signed [`InBus]		in_6_19_i;
wire signed [`InBus]		in_6_20_r;
wire signed [`InBus]		in_6_20_i;
wire signed [`InBus]		in_6_21_r;
wire signed [`InBus]		in_6_21_i;
wire signed [`InBus]		in_6_22_r;
wire signed [`InBus]		in_6_22_i;
wire signed [`InBus]		in_6_23_r;
wire signed [`InBus]		in_6_23_i;
wire signed [`InBus]		in_6_24_r;
wire signed [`InBus]		in_6_24_i;
wire signed [`InBus]		in_6_25_r;
wire signed [`InBus]		in_6_25_i;
wire signed [`InBus]		in_6_26_r;
wire signed [`InBus]		in_6_26_i;
wire signed [`InBus]		in_6_27_r;
wire signed [`InBus]		in_6_27_i;
wire signed [`InBus]		in_6_28_r;
wire signed [`InBus]		in_6_28_i;
wire signed [`InBus]		in_6_29_r;
wire signed [`InBus]		in_6_29_i;
wire signed [`InBus]		in_6_30_r;
wire signed [`InBus]		in_6_30_i;
wire signed [`InBus]		in_6_31_r;
wire signed [`InBus]		in_6_31_i;
wire signed [`InBus]		in_6_32_r;
wire signed [`InBus]		in_6_32_i;
wire signed [`InBus]		in_7_1_r;
wire signed [`InBus]		in_7_1_i;
wire signed [`InBus]		in_7_2_r;
wire signed [`InBus]		in_7_2_i;
wire signed [`InBus]		in_7_3_r;
wire signed [`InBus]		in_7_3_i;
wire signed [`InBus]		in_7_4_r;
wire signed [`InBus]		in_7_4_i;
wire signed [`InBus]		in_7_5_r;
wire signed [`InBus]		in_7_5_i;
wire signed [`InBus]		in_7_6_r;
wire signed [`InBus]		in_7_6_i;
wire signed [`InBus]		in_7_7_r;
wire signed [`InBus]		in_7_7_i;
wire signed [`InBus]		in_7_8_r;
wire signed [`InBus]		in_7_8_i;
wire signed [`InBus]		in_7_9_r;
wire signed [`InBus]		in_7_9_i;
wire signed [`InBus]		in_7_10_r;
wire signed [`InBus]		in_7_10_i;
wire signed [`InBus]		in_7_11_r;
wire signed [`InBus]		in_7_11_i;
wire signed [`InBus]		in_7_12_r;
wire signed [`InBus]		in_7_12_i;
wire signed [`InBus]		in_7_13_r;
wire signed [`InBus]		in_7_13_i;
wire signed [`InBus]		in_7_14_r;
wire signed [`InBus]		in_7_14_i;
wire signed [`InBus]		in_7_15_r;
wire signed [`InBus]		in_7_15_i;
wire signed [`InBus]		in_7_16_r;
wire signed [`InBus]		in_7_16_i;
wire signed [`InBus]		in_7_17_r;
wire signed [`InBus]		in_7_17_i;
wire signed [`InBus]		in_7_18_r;
wire signed [`InBus]		in_7_18_i;
wire signed [`InBus]		in_7_19_r;
wire signed [`InBus]		in_7_19_i;
wire signed [`InBus]		in_7_20_r;
wire signed [`InBus]		in_7_20_i;
wire signed [`InBus]		in_7_21_r;
wire signed [`InBus]		in_7_21_i;
wire signed [`InBus]		in_7_22_r;
wire signed [`InBus]		in_7_22_i;
wire signed [`InBus]		in_7_23_r;
wire signed [`InBus]		in_7_23_i;
wire signed [`InBus]		in_7_24_r;
wire signed [`InBus]		in_7_24_i;
wire signed [`InBus]		in_7_25_r;
wire signed [`InBus]		in_7_25_i;
wire signed [`InBus]		in_7_26_r;
wire signed [`InBus]		in_7_26_i;
wire signed [`InBus]		in_7_27_r;
wire signed [`InBus]		in_7_27_i;
wire signed [`InBus]		in_7_28_r;
wire signed [`InBus]		in_7_28_i;
wire signed [`InBus]		in_7_29_r;
wire signed [`InBus]		in_7_29_i;
wire signed [`InBus]		in_7_30_r;
wire signed [`InBus]		in_7_30_i;
wire signed [`InBus]		in_7_31_r;
wire signed [`InBus]		in_7_31_i;
wire signed [`InBus]		in_7_32_r;
wire signed [`InBus]		in_7_32_i;
wire signed [`InBus]		in_8_1_r;
wire signed [`InBus]		in_8_1_i;
wire signed [`InBus]		in_8_2_r;
wire signed [`InBus]		in_8_2_i;
wire signed [`InBus]		in_8_3_r;
wire signed [`InBus]		in_8_3_i;
wire signed [`InBus]		in_8_4_r;
wire signed [`InBus]		in_8_4_i;
wire signed [`InBus]		in_8_5_r;
wire signed [`InBus]		in_8_5_i;
wire signed [`InBus]		in_8_6_r;
wire signed [`InBus]		in_8_6_i;
wire signed [`InBus]		in_8_7_r;
wire signed [`InBus]		in_8_7_i;
wire signed [`InBus]		in_8_8_r;
wire signed [`InBus]		in_8_8_i;
wire signed [`InBus]		in_8_9_r;
wire signed [`InBus]		in_8_9_i;
wire signed [`InBus]		in_8_10_r;
wire signed [`InBus]		in_8_10_i;
wire signed [`InBus]		in_8_11_r;
wire signed [`InBus]		in_8_11_i;
wire signed [`InBus]		in_8_12_r;
wire signed [`InBus]		in_8_12_i;
wire signed [`InBus]		in_8_13_r;
wire signed [`InBus]		in_8_13_i;
wire signed [`InBus]		in_8_14_r;
wire signed [`InBus]		in_8_14_i;
wire signed [`InBus]		in_8_15_r;
wire signed [`InBus]		in_8_15_i;
wire signed [`InBus]		in_8_16_r;
wire signed [`InBus]		in_8_16_i;
wire signed [`InBus]		in_8_17_r;
wire signed [`InBus]		in_8_17_i;
wire signed [`InBus]		in_8_18_r;
wire signed [`InBus]		in_8_18_i;
wire signed [`InBus]		in_8_19_r;
wire signed [`InBus]		in_8_19_i;
wire signed [`InBus]		in_8_20_r;
wire signed [`InBus]		in_8_20_i;
wire signed [`InBus]		in_8_21_r;
wire signed [`InBus]		in_8_21_i;
wire signed [`InBus]		in_8_22_r;
wire signed [`InBus]		in_8_22_i;
wire signed [`InBus]		in_8_23_r;
wire signed [`InBus]		in_8_23_i;
wire signed [`InBus]		in_8_24_r;
wire signed [`InBus]		in_8_24_i;
wire signed [`InBus]		in_8_25_r;
wire signed [`InBus]		in_8_25_i;
wire signed [`InBus]		in_8_26_r;
wire signed [`InBus]		in_8_26_i;
wire signed [`InBus]		in_8_27_r;
wire signed [`InBus]		in_8_27_i;
wire signed [`InBus]		in_8_28_r;
wire signed [`InBus]		in_8_28_i;
wire signed [`InBus]		in_8_29_r;
wire signed [`InBus]		in_8_29_i;
wire signed [`InBus]		in_8_30_r;
wire signed [`InBus]		in_8_30_i;
wire signed [`InBus]		in_8_31_r;
wire signed [`InBus]		in_8_31_i;
wire signed [`InBus]		in_8_32_r;
wire signed [`InBus]		in_8_32_i;
wire signed [`InBus]		in_9_1_r;
wire signed [`InBus]		in_9_1_i;
wire signed [`InBus]		in_9_2_r;
wire signed [`InBus]		in_9_2_i;
wire signed [`InBus]		in_9_3_r;
wire signed [`InBus]		in_9_3_i;
wire signed [`InBus]		in_9_4_r;
wire signed [`InBus]		in_9_4_i;
wire signed [`InBus]		in_9_5_r;
wire signed [`InBus]		in_9_5_i;
wire signed [`InBus]		in_9_6_r;
wire signed [`InBus]		in_9_6_i;
wire signed [`InBus]		in_9_7_r;
wire signed [`InBus]		in_9_7_i;
wire signed [`InBus]		in_9_8_r;
wire signed [`InBus]		in_9_8_i;
wire signed [`InBus]		in_9_9_r;
wire signed [`InBus]		in_9_9_i;
wire signed [`InBus]		in_9_10_r;
wire signed [`InBus]		in_9_10_i;
wire signed [`InBus]		in_9_11_r;
wire signed [`InBus]		in_9_11_i;
wire signed [`InBus]		in_9_12_r;
wire signed [`InBus]		in_9_12_i;
wire signed [`InBus]		in_9_13_r;
wire signed [`InBus]		in_9_13_i;
wire signed [`InBus]		in_9_14_r;
wire signed [`InBus]		in_9_14_i;
wire signed [`InBus]		in_9_15_r;
wire signed [`InBus]		in_9_15_i;
wire signed [`InBus]		in_9_16_r;
wire signed [`InBus]		in_9_16_i;
wire signed [`InBus]		in_9_17_r;
wire signed [`InBus]		in_9_17_i;
wire signed [`InBus]		in_9_18_r;
wire signed [`InBus]		in_9_18_i;
wire signed [`InBus]		in_9_19_r;
wire signed [`InBus]		in_9_19_i;
wire signed [`InBus]		in_9_20_r;
wire signed [`InBus]		in_9_20_i;
wire signed [`InBus]		in_9_21_r;
wire signed [`InBus]		in_9_21_i;
wire signed [`InBus]		in_9_22_r;
wire signed [`InBus]		in_9_22_i;
wire signed [`InBus]		in_9_23_r;
wire signed [`InBus]		in_9_23_i;
wire signed [`InBus]		in_9_24_r;
wire signed [`InBus]		in_9_24_i;
wire signed [`InBus]		in_9_25_r;
wire signed [`InBus]		in_9_25_i;
wire signed [`InBus]		in_9_26_r;
wire signed [`InBus]		in_9_26_i;
wire signed [`InBus]		in_9_27_r;
wire signed [`InBus]		in_9_27_i;
wire signed [`InBus]		in_9_28_r;
wire signed [`InBus]		in_9_28_i;
wire signed [`InBus]		in_9_29_r;
wire signed [`InBus]		in_9_29_i;
wire signed [`InBus]		in_9_30_r;
wire signed [`InBus]		in_9_30_i;
wire signed [`InBus]		in_9_31_r;
wire signed [`InBus]		in_9_31_i;
wire signed [`InBus]		in_9_32_r;
wire signed [`InBus]		in_9_32_i;
wire signed [`InBus]		in_10_1_r;
wire signed [`InBus]		in_10_1_i;
wire signed [`InBus]		in_10_2_r;
wire signed [`InBus]		in_10_2_i;
wire signed [`InBus]		in_10_3_r;
wire signed [`InBus]		in_10_3_i;
wire signed [`InBus]		in_10_4_r;
wire signed [`InBus]		in_10_4_i;
wire signed [`InBus]		in_10_5_r;
wire signed [`InBus]		in_10_5_i;
wire signed [`InBus]		in_10_6_r;
wire signed [`InBus]		in_10_6_i;
wire signed [`InBus]		in_10_7_r;
wire signed [`InBus]		in_10_7_i;
wire signed [`InBus]		in_10_8_r;
wire signed [`InBus]		in_10_8_i;
wire signed [`InBus]		in_10_9_r;
wire signed [`InBus]		in_10_9_i;
wire signed [`InBus]		in_10_10_r;
wire signed [`InBus]		in_10_10_i;
wire signed [`InBus]		in_10_11_r;
wire signed [`InBus]		in_10_11_i;
wire signed [`InBus]		in_10_12_r;
wire signed [`InBus]		in_10_12_i;
wire signed [`InBus]		in_10_13_r;
wire signed [`InBus]		in_10_13_i;
wire signed [`InBus]		in_10_14_r;
wire signed [`InBus]		in_10_14_i;
wire signed [`InBus]		in_10_15_r;
wire signed [`InBus]		in_10_15_i;
wire signed [`InBus]		in_10_16_r;
wire signed [`InBus]		in_10_16_i;
wire signed [`InBus]		in_10_17_r;
wire signed [`InBus]		in_10_17_i;
wire signed [`InBus]		in_10_18_r;
wire signed [`InBus]		in_10_18_i;
wire signed [`InBus]		in_10_19_r;
wire signed [`InBus]		in_10_19_i;
wire signed [`InBus]		in_10_20_r;
wire signed [`InBus]		in_10_20_i;
wire signed [`InBus]		in_10_21_r;
wire signed [`InBus]		in_10_21_i;
wire signed [`InBus]		in_10_22_r;
wire signed [`InBus]		in_10_22_i;
wire signed [`InBus]		in_10_23_r;
wire signed [`InBus]		in_10_23_i;
wire signed [`InBus]		in_10_24_r;
wire signed [`InBus]		in_10_24_i;
wire signed [`InBus]		in_10_25_r;
wire signed [`InBus]		in_10_25_i;
wire signed [`InBus]		in_10_26_r;
wire signed [`InBus]		in_10_26_i;
wire signed [`InBus]		in_10_27_r;
wire signed [`InBus]		in_10_27_i;
wire signed [`InBus]		in_10_28_r;
wire signed [`InBus]		in_10_28_i;
wire signed [`InBus]		in_10_29_r;
wire signed [`InBus]		in_10_29_i;
wire signed [`InBus]		in_10_30_r;
wire signed [`InBus]		in_10_30_i;
wire signed [`InBus]		in_10_31_r;
wire signed [`InBus]		in_10_31_i;
wire signed [`InBus]		in_10_32_r;
wire signed [`InBus]		in_10_32_i;
wire signed [`InBus]		in_11_1_r;
wire signed [`InBus]		in_11_1_i;
wire signed [`InBus]		in_11_2_r;
wire signed [`InBus]		in_11_2_i;
wire signed [`InBus]		in_11_3_r;
wire signed [`InBus]		in_11_3_i;
wire signed [`InBus]		in_11_4_r;
wire signed [`InBus]		in_11_4_i;
wire signed [`InBus]		in_11_5_r;
wire signed [`InBus]		in_11_5_i;
wire signed [`InBus]		in_11_6_r;
wire signed [`InBus]		in_11_6_i;
wire signed [`InBus]		in_11_7_r;
wire signed [`InBus]		in_11_7_i;
wire signed [`InBus]		in_11_8_r;
wire signed [`InBus]		in_11_8_i;
wire signed [`InBus]		in_11_9_r;
wire signed [`InBus]		in_11_9_i;
wire signed [`InBus]		in_11_10_r;
wire signed [`InBus]		in_11_10_i;
wire signed [`InBus]		in_11_11_r;
wire signed [`InBus]		in_11_11_i;
wire signed [`InBus]		in_11_12_r;
wire signed [`InBus]		in_11_12_i;
wire signed [`InBus]		in_11_13_r;
wire signed [`InBus]		in_11_13_i;
wire signed [`InBus]		in_11_14_r;
wire signed [`InBus]		in_11_14_i;
wire signed [`InBus]		in_11_15_r;
wire signed [`InBus]		in_11_15_i;
wire signed [`InBus]		in_11_16_r;
wire signed [`InBus]		in_11_16_i;
wire signed [`InBus]		in_11_17_r;
wire signed [`InBus]		in_11_17_i;
wire signed [`InBus]		in_11_18_r;
wire signed [`InBus]		in_11_18_i;
wire signed [`InBus]		in_11_19_r;
wire signed [`InBus]		in_11_19_i;
wire signed [`InBus]		in_11_20_r;
wire signed [`InBus]		in_11_20_i;
wire signed [`InBus]		in_11_21_r;
wire signed [`InBus]		in_11_21_i;
wire signed [`InBus]		in_11_22_r;
wire signed [`InBus]		in_11_22_i;
wire signed [`InBus]		in_11_23_r;
wire signed [`InBus]		in_11_23_i;
wire signed [`InBus]		in_11_24_r;
wire signed [`InBus]		in_11_24_i;
wire signed [`InBus]		in_11_25_r;
wire signed [`InBus]		in_11_25_i;
wire signed [`InBus]		in_11_26_r;
wire signed [`InBus]		in_11_26_i;
wire signed [`InBus]		in_11_27_r;
wire signed [`InBus]		in_11_27_i;
wire signed [`InBus]		in_11_28_r;
wire signed [`InBus]		in_11_28_i;
wire signed [`InBus]		in_11_29_r;
wire signed [`InBus]		in_11_29_i;
wire signed [`InBus]		in_11_30_r;
wire signed [`InBus]		in_11_30_i;
wire signed [`InBus]		in_11_31_r;
wire signed [`InBus]		in_11_31_i;
wire signed [`InBus]		in_11_32_r;
wire signed [`InBus]		in_11_32_i;
wire signed [`InBus]		in_12_1_r;
wire signed [`InBus]		in_12_1_i;
wire signed [`InBus]		in_12_2_r;
wire signed [`InBus]		in_12_2_i;
wire signed [`InBus]		in_12_3_r;
wire signed [`InBus]		in_12_3_i;
wire signed [`InBus]		in_12_4_r;
wire signed [`InBus]		in_12_4_i;
wire signed [`InBus]		in_12_5_r;
wire signed [`InBus]		in_12_5_i;
wire signed [`InBus]		in_12_6_r;
wire signed [`InBus]		in_12_6_i;
wire signed [`InBus]		in_12_7_r;
wire signed [`InBus]		in_12_7_i;
wire signed [`InBus]		in_12_8_r;
wire signed [`InBus]		in_12_8_i;
wire signed [`InBus]		in_12_9_r;
wire signed [`InBus]		in_12_9_i;
wire signed [`InBus]		in_12_10_r;
wire signed [`InBus]		in_12_10_i;
wire signed [`InBus]		in_12_11_r;
wire signed [`InBus]		in_12_11_i;
wire signed [`InBus]		in_12_12_r;
wire signed [`InBus]		in_12_12_i;
wire signed [`InBus]		in_12_13_r;
wire signed [`InBus]		in_12_13_i;
wire signed [`InBus]		in_12_14_r;
wire signed [`InBus]		in_12_14_i;
wire signed [`InBus]		in_12_15_r;
wire signed [`InBus]		in_12_15_i;
wire signed [`InBus]		in_12_16_r;
wire signed [`InBus]		in_12_16_i;
wire signed [`InBus]		in_12_17_r;
wire signed [`InBus]		in_12_17_i;
wire signed [`InBus]		in_12_18_r;
wire signed [`InBus]		in_12_18_i;
wire signed [`InBus]		in_12_19_r;
wire signed [`InBus]		in_12_19_i;
wire signed [`InBus]		in_12_20_r;
wire signed [`InBus]		in_12_20_i;
wire signed [`InBus]		in_12_21_r;
wire signed [`InBus]		in_12_21_i;
wire signed [`InBus]		in_12_22_r;
wire signed [`InBus]		in_12_22_i;
wire signed [`InBus]		in_12_23_r;
wire signed [`InBus]		in_12_23_i;
wire signed [`InBus]		in_12_24_r;
wire signed [`InBus]		in_12_24_i;
wire signed [`InBus]		in_12_25_r;
wire signed [`InBus]		in_12_25_i;
wire signed [`InBus]		in_12_26_r;
wire signed [`InBus]		in_12_26_i;
wire signed [`InBus]		in_12_27_r;
wire signed [`InBus]		in_12_27_i;
wire signed [`InBus]		in_12_28_r;
wire signed [`InBus]		in_12_28_i;
wire signed [`InBus]		in_12_29_r;
wire signed [`InBus]		in_12_29_i;
wire signed [`InBus]		in_12_30_r;
wire signed [`InBus]		in_12_30_i;
wire signed [`InBus]		in_12_31_r;
wire signed [`InBus]		in_12_31_i;
wire signed [`InBus]		in_12_32_r;
wire signed [`InBus]		in_12_32_i;
wire signed [`InBus]		in_13_1_r;
wire signed [`InBus]		in_13_1_i;
wire signed [`InBus]		in_13_2_r;
wire signed [`InBus]		in_13_2_i;
wire signed [`InBus]		in_13_3_r;
wire signed [`InBus]		in_13_3_i;
wire signed [`InBus]		in_13_4_r;
wire signed [`InBus]		in_13_4_i;
wire signed [`InBus]		in_13_5_r;
wire signed [`InBus]		in_13_5_i;
wire signed [`InBus]		in_13_6_r;
wire signed [`InBus]		in_13_6_i;
wire signed [`InBus]		in_13_7_r;
wire signed [`InBus]		in_13_7_i;
wire signed [`InBus]		in_13_8_r;
wire signed [`InBus]		in_13_8_i;
wire signed [`InBus]		in_13_9_r;
wire signed [`InBus]		in_13_9_i;
wire signed [`InBus]		in_13_10_r;
wire signed [`InBus]		in_13_10_i;
wire signed [`InBus]		in_13_11_r;
wire signed [`InBus]		in_13_11_i;
wire signed [`InBus]		in_13_12_r;
wire signed [`InBus]		in_13_12_i;
wire signed [`InBus]		in_13_13_r;
wire signed [`InBus]		in_13_13_i;
wire signed [`InBus]		in_13_14_r;
wire signed [`InBus]		in_13_14_i;
wire signed [`InBus]		in_13_15_r;
wire signed [`InBus]		in_13_15_i;
wire signed [`InBus]		in_13_16_r;
wire signed [`InBus]		in_13_16_i;
wire signed [`InBus]		in_13_17_r;
wire signed [`InBus]		in_13_17_i;
wire signed [`InBus]		in_13_18_r;
wire signed [`InBus]		in_13_18_i;
wire signed [`InBus]		in_13_19_r;
wire signed [`InBus]		in_13_19_i;
wire signed [`InBus]		in_13_20_r;
wire signed [`InBus]		in_13_20_i;
wire signed [`InBus]		in_13_21_r;
wire signed [`InBus]		in_13_21_i;
wire signed [`InBus]		in_13_22_r;
wire signed [`InBus]		in_13_22_i;
wire signed [`InBus]		in_13_23_r;
wire signed [`InBus]		in_13_23_i;
wire signed [`InBus]		in_13_24_r;
wire signed [`InBus]		in_13_24_i;
wire signed [`InBus]		in_13_25_r;
wire signed [`InBus]		in_13_25_i;
wire signed [`InBus]		in_13_26_r;
wire signed [`InBus]		in_13_26_i;
wire signed [`InBus]		in_13_27_r;
wire signed [`InBus]		in_13_27_i;
wire signed [`InBus]		in_13_28_r;
wire signed [`InBus]		in_13_28_i;
wire signed [`InBus]		in_13_29_r;
wire signed [`InBus]		in_13_29_i;
wire signed [`InBus]		in_13_30_r;
wire signed [`InBus]		in_13_30_i;
wire signed [`InBus]		in_13_31_r;
wire signed [`InBus]		in_13_31_i;
wire signed [`InBus]		in_13_32_r;
wire signed [`InBus]		in_13_32_i;
wire signed [`InBus]		in_14_1_r;
wire signed [`InBus]		in_14_1_i;
wire signed [`InBus]		in_14_2_r;
wire signed [`InBus]		in_14_2_i;
wire signed [`InBus]		in_14_3_r;
wire signed [`InBus]		in_14_3_i;
wire signed [`InBus]		in_14_4_r;
wire signed [`InBus]		in_14_4_i;
wire signed [`InBus]		in_14_5_r;
wire signed [`InBus]		in_14_5_i;
wire signed [`InBus]		in_14_6_r;
wire signed [`InBus]		in_14_6_i;
wire signed [`InBus]		in_14_7_r;
wire signed [`InBus]		in_14_7_i;
wire signed [`InBus]		in_14_8_r;
wire signed [`InBus]		in_14_8_i;
wire signed [`InBus]		in_14_9_r;
wire signed [`InBus]		in_14_9_i;
wire signed [`InBus]		in_14_10_r;
wire signed [`InBus]		in_14_10_i;
wire signed [`InBus]		in_14_11_r;
wire signed [`InBus]		in_14_11_i;
wire signed [`InBus]		in_14_12_r;
wire signed [`InBus]		in_14_12_i;
wire signed [`InBus]		in_14_13_r;
wire signed [`InBus]		in_14_13_i;
wire signed [`InBus]		in_14_14_r;
wire signed [`InBus]		in_14_14_i;
wire signed [`InBus]		in_14_15_r;
wire signed [`InBus]		in_14_15_i;
wire signed [`InBus]		in_14_16_r;
wire signed [`InBus]		in_14_16_i;
wire signed [`InBus]		in_14_17_r;
wire signed [`InBus]		in_14_17_i;
wire signed [`InBus]		in_14_18_r;
wire signed [`InBus]		in_14_18_i;
wire signed [`InBus]		in_14_19_r;
wire signed [`InBus]		in_14_19_i;
wire signed [`InBus]		in_14_20_r;
wire signed [`InBus]		in_14_20_i;
wire signed [`InBus]		in_14_21_r;
wire signed [`InBus]		in_14_21_i;
wire signed [`InBus]		in_14_22_r;
wire signed [`InBus]		in_14_22_i;
wire signed [`InBus]		in_14_23_r;
wire signed [`InBus]		in_14_23_i;
wire signed [`InBus]		in_14_24_r;
wire signed [`InBus]		in_14_24_i;
wire signed [`InBus]		in_14_25_r;
wire signed [`InBus]		in_14_25_i;
wire signed [`InBus]		in_14_26_r;
wire signed [`InBus]		in_14_26_i;
wire signed [`InBus]		in_14_27_r;
wire signed [`InBus]		in_14_27_i;
wire signed [`InBus]		in_14_28_r;
wire signed [`InBus]		in_14_28_i;
wire signed [`InBus]		in_14_29_r;
wire signed [`InBus]		in_14_29_i;
wire signed [`InBus]		in_14_30_r;
wire signed [`InBus]		in_14_30_i;
wire signed [`InBus]		in_14_31_r;
wire signed [`InBus]		in_14_31_i;
wire signed [`InBus]		in_14_32_r;
wire signed [`InBus]		in_14_32_i;
wire signed [`InBus]		in_15_1_r;
wire signed [`InBus]		in_15_1_i;
wire signed [`InBus]		in_15_2_r;
wire signed [`InBus]		in_15_2_i;
wire signed [`InBus]		in_15_3_r;
wire signed [`InBus]		in_15_3_i;
wire signed [`InBus]		in_15_4_r;
wire signed [`InBus]		in_15_4_i;
wire signed [`InBus]		in_15_5_r;
wire signed [`InBus]		in_15_5_i;
wire signed [`InBus]		in_15_6_r;
wire signed [`InBus]		in_15_6_i;
wire signed [`InBus]		in_15_7_r;
wire signed [`InBus]		in_15_7_i;
wire signed [`InBus]		in_15_8_r;
wire signed [`InBus]		in_15_8_i;
wire signed [`InBus]		in_15_9_r;
wire signed [`InBus]		in_15_9_i;
wire signed [`InBus]		in_15_10_r;
wire signed [`InBus]		in_15_10_i;
wire signed [`InBus]		in_15_11_r;
wire signed [`InBus]		in_15_11_i;
wire signed [`InBus]		in_15_12_r;
wire signed [`InBus]		in_15_12_i;
wire signed [`InBus]		in_15_13_r;
wire signed [`InBus]		in_15_13_i;
wire signed [`InBus]		in_15_14_r;
wire signed [`InBus]		in_15_14_i;
wire signed [`InBus]		in_15_15_r;
wire signed [`InBus]		in_15_15_i;
wire signed [`InBus]		in_15_16_r;
wire signed [`InBus]		in_15_16_i;
wire signed [`InBus]		in_15_17_r;
wire signed [`InBus]		in_15_17_i;
wire signed [`InBus]		in_15_18_r;
wire signed [`InBus]		in_15_18_i;
wire signed [`InBus]		in_15_19_r;
wire signed [`InBus]		in_15_19_i;
wire signed [`InBus]		in_15_20_r;
wire signed [`InBus]		in_15_20_i;
wire signed [`InBus]		in_15_21_r;
wire signed [`InBus]		in_15_21_i;
wire signed [`InBus]		in_15_22_r;
wire signed [`InBus]		in_15_22_i;
wire signed [`InBus]		in_15_23_r;
wire signed [`InBus]		in_15_23_i;
wire signed [`InBus]		in_15_24_r;
wire signed [`InBus]		in_15_24_i;
wire signed [`InBus]		in_15_25_r;
wire signed [`InBus]		in_15_25_i;
wire signed [`InBus]		in_15_26_r;
wire signed [`InBus]		in_15_26_i;
wire signed [`InBus]		in_15_27_r;
wire signed [`InBus]		in_15_27_i;
wire signed [`InBus]		in_15_28_r;
wire signed [`InBus]		in_15_28_i;
wire signed [`InBus]		in_15_29_r;
wire signed [`InBus]		in_15_29_i;
wire signed [`InBus]		in_15_30_r;
wire signed [`InBus]		in_15_30_i;
wire signed [`InBus]		in_15_31_r;
wire signed [`InBus]		in_15_31_i;
wire signed [`InBus]		in_15_32_r;
wire signed [`InBus]		in_15_32_i;
wire signed [`InBus]		in_16_1_r;
wire signed [`InBus]		in_16_1_i;
wire signed [`InBus]		in_16_2_r;
wire signed [`InBus]		in_16_2_i;
wire signed [`InBus]		in_16_3_r;
wire signed [`InBus]		in_16_3_i;
wire signed [`InBus]		in_16_4_r;
wire signed [`InBus]		in_16_4_i;
wire signed [`InBus]		in_16_5_r;
wire signed [`InBus]		in_16_5_i;
wire signed [`InBus]		in_16_6_r;
wire signed [`InBus]		in_16_6_i;
wire signed [`InBus]		in_16_7_r;
wire signed [`InBus]		in_16_7_i;
wire signed [`InBus]		in_16_8_r;
wire signed [`InBus]		in_16_8_i;
wire signed [`InBus]		in_16_9_r;
wire signed [`InBus]		in_16_9_i;
wire signed [`InBus]		in_16_10_r;
wire signed [`InBus]		in_16_10_i;
wire signed [`InBus]		in_16_11_r;
wire signed [`InBus]		in_16_11_i;
wire signed [`InBus]		in_16_12_r;
wire signed [`InBus]		in_16_12_i;
wire signed [`InBus]		in_16_13_r;
wire signed [`InBus]		in_16_13_i;
wire signed [`InBus]		in_16_14_r;
wire signed [`InBus]		in_16_14_i;
wire signed [`InBus]		in_16_15_r;
wire signed [`InBus]		in_16_15_i;
wire signed [`InBus]		in_16_16_r;
wire signed [`InBus]		in_16_16_i;
wire signed [`InBus]		in_16_17_r;
wire signed [`InBus]		in_16_17_i;
wire signed [`InBus]		in_16_18_r;
wire signed [`InBus]		in_16_18_i;
wire signed [`InBus]		in_16_19_r;
wire signed [`InBus]		in_16_19_i;
wire signed [`InBus]		in_16_20_r;
wire signed [`InBus]		in_16_20_i;
wire signed [`InBus]		in_16_21_r;
wire signed [`InBus]		in_16_21_i;
wire signed [`InBus]		in_16_22_r;
wire signed [`InBus]		in_16_22_i;
wire signed [`InBus]		in_16_23_r;
wire signed [`InBus]		in_16_23_i;
wire signed [`InBus]		in_16_24_r;
wire signed [`InBus]		in_16_24_i;
wire signed [`InBus]		in_16_25_r;
wire signed [`InBus]		in_16_25_i;
wire signed [`InBus]		in_16_26_r;
wire signed [`InBus]		in_16_26_i;
wire signed [`InBus]		in_16_27_r;
wire signed [`InBus]		in_16_27_i;
wire signed [`InBus]		in_16_28_r;
wire signed [`InBus]		in_16_28_i;
wire signed [`InBus]		in_16_29_r;
wire signed [`InBus]		in_16_29_i;
wire signed [`InBus]		in_16_30_r;
wire signed [`InBus]		in_16_30_i;
wire signed [`InBus]		in_16_31_r;
wire signed [`InBus]		in_16_31_i;
wire signed [`InBus]		in_16_32_r;
wire signed [`InBus]		in_16_32_i;
wire signed [`InBus]		in_17_1_r;
wire signed [`InBus]		in_17_1_i;
wire signed [`InBus]		in_17_2_r;
wire signed [`InBus]		in_17_2_i;
wire signed [`InBus]		in_17_3_r;
wire signed [`InBus]		in_17_3_i;
wire signed [`InBus]		in_17_4_r;
wire signed [`InBus]		in_17_4_i;
wire signed [`InBus]		in_17_5_r;
wire signed [`InBus]		in_17_5_i;
wire signed [`InBus]		in_17_6_r;
wire signed [`InBus]		in_17_6_i;
wire signed [`InBus]		in_17_7_r;
wire signed [`InBus]		in_17_7_i;
wire signed [`InBus]		in_17_8_r;
wire signed [`InBus]		in_17_8_i;
wire signed [`InBus]		in_17_9_r;
wire signed [`InBus]		in_17_9_i;
wire signed [`InBus]		in_17_10_r;
wire signed [`InBus]		in_17_10_i;
wire signed [`InBus]		in_17_11_r;
wire signed [`InBus]		in_17_11_i;
wire signed [`InBus]		in_17_12_r;
wire signed [`InBus]		in_17_12_i;
wire signed [`InBus]		in_17_13_r;
wire signed [`InBus]		in_17_13_i;
wire signed [`InBus]		in_17_14_r;
wire signed [`InBus]		in_17_14_i;
wire signed [`InBus]		in_17_15_r;
wire signed [`InBus]		in_17_15_i;
wire signed [`InBus]		in_17_16_r;
wire signed [`InBus]		in_17_16_i;
wire signed [`InBus]		in_17_17_r;
wire signed [`InBus]		in_17_17_i;
wire signed [`InBus]		in_17_18_r;
wire signed [`InBus]		in_17_18_i;
wire signed [`InBus]		in_17_19_r;
wire signed [`InBus]		in_17_19_i;
wire signed [`InBus]		in_17_20_r;
wire signed [`InBus]		in_17_20_i;
wire signed [`InBus]		in_17_21_r;
wire signed [`InBus]		in_17_21_i;
wire signed [`InBus]		in_17_22_r;
wire signed [`InBus]		in_17_22_i;
wire signed [`InBus]		in_17_23_r;
wire signed [`InBus]		in_17_23_i;
wire signed [`InBus]		in_17_24_r;
wire signed [`InBus]		in_17_24_i;
wire signed [`InBus]		in_17_25_r;
wire signed [`InBus]		in_17_25_i;
wire signed [`InBus]		in_17_26_r;
wire signed [`InBus]		in_17_26_i;
wire signed [`InBus]		in_17_27_r;
wire signed [`InBus]		in_17_27_i;
wire signed [`InBus]		in_17_28_r;
wire signed [`InBus]		in_17_28_i;
wire signed [`InBus]		in_17_29_r;
wire signed [`InBus]		in_17_29_i;
wire signed [`InBus]		in_17_30_r;
wire signed [`InBus]		in_17_30_i;
wire signed [`InBus]		in_17_31_r;
wire signed [`InBus]		in_17_31_i;
wire signed [`InBus]		in_17_32_r;
wire signed [`InBus]		in_17_32_i;
wire signed [`InBus]		in_18_1_r;
wire signed [`InBus]		in_18_1_i;
wire signed [`InBus]		in_18_2_r;
wire signed [`InBus]		in_18_2_i;
wire signed [`InBus]		in_18_3_r;
wire signed [`InBus]		in_18_3_i;
wire signed [`InBus]		in_18_4_r;
wire signed [`InBus]		in_18_4_i;
wire signed [`InBus]		in_18_5_r;
wire signed [`InBus]		in_18_5_i;
wire signed [`InBus]		in_18_6_r;
wire signed [`InBus]		in_18_6_i;
wire signed [`InBus]		in_18_7_r;
wire signed [`InBus]		in_18_7_i;
wire signed [`InBus]		in_18_8_r;
wire signed [`InBus]		in_18_8_i;
wire signed [`InBus]		in_18_9_r;
wire signed [`InBus]		in_18_9_i;
wire signed [`InBus]		in_18_10_r;
wire signed [`InBus]		in_18_10_i;
wire signed [`InBus]		in_18_11_r;
wire signed [`InBus]		in_18_11_i;
wire signed [`InBus]		in_18_12_r;
wire signed [`InBus]		in_18_12_i;
wire signed [`InBus]		in_18_13_r;
wire signed [`InBus]		in_18_13_i;
wire signed [`InBus]		in_18_14_r;
wire signed [`InBus]		in_18_14_i;
wire signed [`InBus]		in_18_15_r;
wire signed [`InBus]		in_18_15_i;
wire signed [`InBus]		in_18_16_r;
wire signed [`InBus]		in_18_16_i;
wire signed [`InBus]		in_18_17_r;
wire signed [`InBus]		in_18_17_i;
wire signed [`InBus]		in_18_18_r;
wire signed [`InBus]		in_18_18_i;
wire signed [`InBus]		in_18_19_r;
wire signed [`InBus]		in_18_19_i;
wire signed [`InBus]		in_18_20_r;
wire signed [`InBus]		in_18_20_i;
wire signed [`InBus]		in_18_21_r;
wire signed [`InBus]		in_18_21_i;
wire signed [`InBus]		in_18_22_r;
wire signed [`InBus]		in_18_22_i;
wire signed [`InBus]		in_18_23_r;
wire signed [`InBus]		in_18_23_i;
wire signed [`InBus]		in_18_24_r;
wire signed [`InBus]		in_18_24_i;
wire signed [`InBus]		in_18_25_r;
wire signed [`InBus]		in_18_25_i;
wire signed [`InBus]		in_18_26_r;
wire signed [`InBus]		in_18_26_i;
wire signed [`InBus]		in_18_27_r;
wire signed [`InBus]		in_18_27_i;
wire signed [`InBus]		in_18_28_r;
wire signed [`InBus]		in_18_28_i;
wire signed [`InBus]		in_18_29_r;
wire signed [`InBus]		in_18_29_i;
wire signed [`InBus]		in_18_30_r;
wire signed [`InBus]		in_18_30_i;
wire signed [`InBus]		in_18_31_r;
wire signed [`InBus]		in_18_31_i;
wire signed [`InBus]		in_18_32_r;
wire signed [`InBus]		in_18_32_i;
wire signed [`InBus]		in_19_1_r;
wire signed [`InBus]		in_19_1_i;
wire signed [`InBus]		in_19_2_r;
wire signed [`InBus]		in_19_2_i;
wire signed [`InBus]		in_19_3_r;
wire signed [`InBus]		in_19_3_i;
wire signed [`InBus]		in_19_4_r;
wire signed [`InBus]		in_19_4_i;
wire signed [`InBus]		in_19_5_r;
wire signed [`InBus]		in_19_5_i;
wire signed [`InBus]		in_19_6_r;
wire signed [`InBus]		in_19_6_i;
wire signed [`InBus]		in_19_7_r;
wire signed [`InBus]		in_19_7_i;
wire signed [`InBus]		in_19_8_r;
wire signed [`InBus]		in_19_8_i;
wire signed [`InBus]		in_19_9_r;
wire signed [`InBus]		in_19_9_i;
wire signed [`InBus]		in_19_10_r;
wire signed [`InBus]		in_19_10_i;
wire signed [`InBus]		in_19_11_r;
wire signed [`InBus]		in_19_11_i;
wire signed [`InBus]		in_19_12_r;
wire signed [`InBus]		in_19_12_i;
wire signed [`InBus]		in_19_13_r;
wire signed [`InBus]		in_19_13_i;
wire signed [`InBus]		in_19_14_r;
wire signed [`InBus]		in_19_14_i;
wire signed [`InBus]		in_19_15_r;
wire signed [`InBus]		in_19_15_i;
wire signed [`InBus]		in_19_16_r;
wire signed [`InBus]		in_19_16_i;
wire signed [`InBus]		in_19_17_r;
wire signed [`InBus]		in_19_17_i;
wire signed [`InBus]		in_19_18_r;
wire signed [`InBus]		in_19_18_i;
wire signed [`InBus]		in_19_19_r;
wire signed [`InBus]		in_19_19_i;
wire signed [`InBus]		in_19_20_r;
wire signed [`InBus]		in_19_20_i;
wire signed [`InBus]		in_19_21_r;
wire signed [`InBus]		in_19_21_i;
wire signed [`InBus]		in_19_22_r;
wire signed [`InBus]		in_19_22_i;
wire signed [`InBus]		in_19_23_r;
wire signed [`InBus]		in_19_23_i;
wire signed [`InBus]		in_19_24_r;
wire signed [`InBus]		in_19_24_i;
wire signed [`InBus]		in_19_25_r;
wire signed [`InBus]		in_19_25_i;
wire signed [`InBus]		in_19_26_r;
wire signed [`InBus]		in_19_26_i;
wire signed [`InBus]		in_19_27_r;
wire signed [`InBus]		in_19_27_i;
wire signed [`InBus]		in_19_28_r;
wire signed [`InBus]		in_19_28_i;
wire signed [`InBus]		in_19_29_r;
wire signed [`InBus]		in_19_29_i;
wire signed [`InBus]		in_19_30_r;
wire signed [`InBus]		in_19_30_i;
wire signed [`InBus]		in_19_31_r;
wire signed [`InBus]		in_19_31_i;
wire signed [`InBus]		in_19_32_r;
wire signed [`InBus]		in_19_32_i;
wire signed [`InBus]		in_20_1_r;
wire signed [`InBus]		in_20_1_i;
wire signed [`InBus]		in_20_2_r;
wire signed [`InBus]		in_20_2_i;
wire signed [`InBus]		in_20_3_r;
wire signed [`InBus]		in_20_3_i;
wire signed [`InBus]		in_20_4_r;
wire signed [`InBus]		in_20_4_i;
wire signed [`InBus]		in_20_5_r;
wire signed [`InBus]		in_20_5_i;
wire signed [`InBus]		in_20_6_r;
wire signed [`InBus]		in_20_6_i;
wire signed [`InBus]		in_20_7_r;
wire signed [`InBus]		in_20_7_i;
wire signed [`InBus]		in_20_8_r;
wire signed [`InBus]		in_20_8_i;
wire signed [`InBus]		in_20_9_r;
wire signed [`InBus]		in_20_9_i;
wire signed [`InBus]		in_20_10_r;
wire signed [`InBus]		in_20_10_i;
wire signed [`InBus]		in_20_11_r;
wire signed [`InBus]		in_20_11_i;
wire signed [`InBus]		in_20_12_r;
wire signed [`InBus]		in_20_12_i;
wire signed [`InBus]		in_20_13_r;
wire signed [`InBus]		in_20_13_i;
wire signed [`InBus]		in_20_14_r;
wire signed [`InBus]		in_20_14_i;
wire signed [`InBus]		in_20_15_r;
wire signed [`InBus]		in_20_15_i;
wire signed [`InBus]		in_20_16_r;
wire signed [`InBus]		in_20_16_i;
wire signed [`InBus]		in_20_17_r;
wire signed [`InBus]		in_20_17_i;
wire signed [`InBus]		in_20_18_r;
wire signed [`InBus]		in_20_18_i;
wire signed [`InBus]		in_20_19_r;
wire signed [`InBus]		in_20_19_i;
wire signed [`InBus]		in_20_20_r;
wire signed [`InBus]		in_20_20_i;
wire signed [`InBus]		in_20_21_r;
wire signed [`InBus]		in_20_21_i;
wire signed [`InBus]		in_20_22_r;
wire signed [`InBus]		in_20_22_i;
wire signed [`InBus]		in_20_23_r;
wire signed [`InBus]		in_20_23_i;
wire signed [`InBus]		in_20_24_r;
wire signed [`InBus]		in_20_24_i;
wire signed [`InBus]		in_20_25_r;
wire signed [`InBus]		in_20_25_i;
wire signed [`InBus]		in_20_26_r;
wire signed [`InBus]		in_20_26_i;
wire signed [`InBus]		in_20_27_r;
wire signed [`InBus]		in_20_27_i;
wire signed [`InBus]		in_20_28_r;
wire signed [`InBus]		in_20_28_i;
wire signed [`InBus]		in_20_29_r;
wire signed [`InBus]		in_20_29_i;
wire signed [`InBus]		in_20_30_r;
wire signed [`InBus]		in_20_30_i;
wire signed [`InBus]		in_20_31_r;
wire signed [`InBus]		in_20_31_i;
wire signed [`InBus]		in_20_32_r;
wire signed [`InBus]		in_20_32_i;
wire signed [`InBus]		in_21_1_r;
wire signed [`InBus]		in_21_1_i;
wire signed [`InBus]		in_21_2_r;
wire signed [`InBus]		in_21_2_i;
wire signed [`InBus]		in_21_3_r;
wire signed [`InBus]		in_21_3_i;
wire signed [`InBus]		in_21_4_r;
wire signed [`InBus]		in_21_4_i;
wire signed [`InBus]		in_21_5_r;
wire signed [`InBus]		in_21_5_i;
wire signed [`InBus]		in_21_6_r;
wire signed [`InBus]		in_21_6_i;
wire signed [`InBus]		in_21_7_r;
wire signed [`InBus]		in_21_7_i;
wire signed [`InBus]		in_21_8_r;
wire signed [`InBus]		in_21_8_i;
wire signed [`InBus]		in_21_9_r;
wire signed [`InBus]		in_21_9_i;
wire signed [`InBus]		in_21_10_r;
wire signed [`InBus]		in_21_10_i;
wire signed [`InBus]		in_21_11_r;
wire signed [`InBus]		in_21_11_i;
wire signed [`InBus]		in_21_12_r;
wire signed [`InBus]		in_21_12_i;
wire signed [`InBus]		in_21_13_r;
wire signed [`InBus]		in_21_13_i;
wire signed [`InBus]		in_21_14_r;
wire signed [`InBus]		in_21_14_i;
wire signed [`InBus]		in_21_15_r;
wire signed [`InBus]		in_21_15_i;
wire signed [`InBus]		in_21_16_r;
wire signed [`InBus]		in_21_16_i;
wire signed [`InBus]		in_21_17_r;
wire signed [`InBus]		in_21_17_i;
wire signed [`InBus]		in_21_18_r;
wire signed [`InBus]		in_21_18_i;
wire signed [`InBus]		in_21_19_r;
wire signed [`InBus]		in_21_19_i;
wire signed [`InBus]		in_21_20_r;
wire signed [`InBus]		in_21_20_i;
wire signed [`InBus]		in_21_21_r;
wire signed [`InBus]		in_21_21_i;
wire signed [`InBus]		in_21_22_r;
wire signed [`InBus]		in_21_22_i;
wire signed [`InBus]		in_21_23_r;
wire signed [`InBus]		in_21_23_i;
wire signed [`InBus]		in_21_24_r;
wire signed [`InBus]		in_21_24_i;
wire signed [`InBus]		in_21_25_r;
wire signed [`InBus]		in_21_25_i;
wire signed [`InBus]		in_21_26_r;
wire signed [`InBus]		in_21_26_i;
wire signed [`InBus]		in_21_27_r;
wire signed [`InBus]		in_21_27_i;
wire signed [`InBus]		in_21_28_r;
wire signed [`InBus]		in_21_28_i;
wire signed [`InBus]		in_21_29_r;
wire signed [`InBus]		in_21_29_i;
wire signed [`InBus]		in_21_30_r;
wire signed [`InBus]		in_21_30_i;
wire signed [`InBus]		in_21_31_r;
wire signed [`InBus]		in_21_31_i;
wire signed [`InBus]		in_21_32_r;
wire signed [`InBus]		in_21_32_i;
wire signed [`InBus]		in_22_1_r;
wire signed [`InBus]		in_22_1_i;
wire signed [`InBus]		in_22_2_r;
wire signed [`InBus]		in_22_2_i;
wire signed [`InBus]		in_22_3_r;
wire signed [`InBus]		in_22_3_i;
wire signed [`InBus]		in_22_4_r;
wire signed [`InBus]		in_22_4_i;
wire signed [`InBus]		in_22_5_r;
wire signed [`InBus]		in_22_5_i;
wire signed [`InBus]		in_22_6_r;
wire signed [`InBus]		in_22_6_i;
wire signed [`InBus]		in_22_7_r;
wire signed [`InBus]		in_22_7_i;
wire signed [`InBus]		in_22_8_r;
wire signed [`InBus]		in_22_8_i;
wire signed [`InBus]		in_22_9_r;
wire signed [`InBus]		in_22_9_i;
wire signed [`InBus]		in_22_10_r;
wire signed [`InBus]		in_22_10_i;
wire signed [`InBus]		in_22_11_r;
wire signed [`InBus]		in_22_11_i;
wire signed [`InBus]		in_22_12_r;
wire signed [`InBus]		in_22_12_i;
wire signed [`InBus]		in_22_13_r;
wire signed [`InBus]		in_22_13_i;
wire signed [`InBus]		in_22_14_r;
wire signed [`InBus]		in_22_14_i;
wire signed [`InBus]		in_22_15_r;
wire signed [`InBus]		in_22_15_i;
wire signed [`InBus]		in_22_16_r;
wire signed [`InBus]		in_22_16_i;
wire signed [`InBus]		in_22_17_r;
wire signed [`InBus]		in_22_17_i;
wire signed [`InBus]		in_22_18_r;
wire signed [`InBus]		in_22_18_i;
wire signed [`InBus]		in_22_19_r;
wire signed [`InBus]		in_22_19_i;
wire signed [`InBus]		in_22_20_r;
wire signed [`InBus]		in_22_20_i;
wire signed [`InBus]		in_22_21_r;
wire signed [`InBus]		in_22_21_i;
wire signed [`InBus]		in_22_22_r;
wire signed [`InBus]		in_22_22_i;
wire signed [`InBus]		in_22_23_r;
wire signed [`InBus]		in_22_23_i;
wire signed [`InBus]		in_22_24_r;
wire signed [`InBus]		in_22_24_i;
wire signed [`InBus]		in_22_25_r;
wire signed [`InBus]		in_22_25_i;
wire signed [`InBus]		in_22_26_r;
wire signed [`InBus]		in_22_26_i;
wire signed [`InBus]		in_22_27_r;
wire signed [`InBus]		in_22_27_i;
wire signed [`InBus]		in_22_28_r;
wire signed [`InBus]		in_22_28_i;
wire signed [`InBus]		in_22_29_r;
wire signed [`InBus]		in_22_29_i;
wire signed [`InBus]		in_22_30_r;
wire signed [`InBus]		in_22_30_i;
wire signed [`InBus]		in_22_31_r;
wire signed [`InBus]		in_22_31_i;
wire signed [`InBus]		in_22_32_r;
wire signed [`InBus]		in_22_32_i;
wire signed [`InBus]		in_23_1_r;
wire signed [`InBus]		in_23_1_i;
wire signed [`InBus]		in_23_2_r;
wire signed [`InBus]		in_23_2_i;
wire signed [`InBus]		in_23_3_r;
wire signed [`InBus]		in_23_3_i;
wire signed [`InBus]		in_23_4_r;
wire signed [`InBus]		in_23_4_i;
wire signed [`InBus]		in_23_5_r;
wire signed [`InBus]		in_23_5_i;
wire signed [`InBus]		in_23_6_r;
wire signed [`InBus]		in_23_6_i;
wire signed [`InBus]		in_23_7_r;
wire signed [`InBus]		in_23_7_i;
wire signed [`InBus]		in_23_8_r;
wire signed [`InBus]		in_23_8_i;
wire signed [`InBus]		in_23_9_r;
wire signed [`InBus]		in_23_9_i;
wire signed [`InBus]		in_23_10_r;
wire signed [`InBus]		in_23_10_i;
wire signed [`InBus]		in_23_11_r;
wire signed [`InBus]		in_23_11_i;
wire signed [`InBus]		in_23_12_r;
wire signed [`InBus]		in_23_12_i;
wire signed [`InBus]		in_23_13_r;
wire signed [`InBus]		in_23_13_i;
wire signed [`InBus]		in_23_14_r;
wire signed [`InBus]		in_23_14_i;
wire signed [`InBus]		in_23_15_r;
wire signed [`InBus]		in_23_15_i;
wire signed [`InBus]		in_23_16_r;
wire signed [`InBus]		in_23_16_i;
wire signed [`InBus]		in_23_17_r;
wire signed [`InBus]		in_23_17_i;
wire signed [`InBus]		in_23_18_r;
wire signed [`InBus]		in_23_18_i;
wire signed [`InBus]		in_23_19_r;
wire signed [`InBus]		in_23_19_i;
wire signed [`InBus]		in_23_20_r;
wire signed [`InBus]		in_23_20_i;
wire signed [`InBus]		in_23_21_r;
wire signed [`InBus]		in_23_21_i;
wire signed [`InBus]		in_23_22_r;
wire signed [`InBus]		in_23_22_i;
wire signed [`InBus]		in_23_23_r;
wire signed [`InBus]		in_23_23_i;
wire signed [`InBus]		in_23_24_r;
wire signed [`InBus]		in_23_24_i;
wire signed [`InBus]		in_23_25_r;
wire signed [`InBus]		in_23_25_i;
wire signed [`InBus]		in_23_26_r;
wire signed [`InBus]		in_23_26_i;
wire signed [`InBus]		in_23_27_r;
wire signed [`InBus]		in_23_27_i;
wire signed [`InBus]		in_23_28_r;
wire signed [`InBus]		in_23_28_i;
wire signed [`InBus]		in_23_29_r;
wire signed [`InBus]		in_23_29_i;
wire signed [`InBus]		in_23_30_r;
wire signed [`InBus]		in_23_30_i;
wire signed [`InBus]		in_23_31_r;
wire signed [`InBus]		in_23_31_i;
wire signed [`InBus]		in_23_32_r;
wire signed [`InBus]		in_23_32_i;
wire signed [`InBus]		in_24_1_r;
wire signed [`InBus]		in_24_1_i;
wire signed [`InBus]		in_24_2_r;
wire signed [`InBus]		in_24_2_i;
wire signed [`InBus]		in_24_3_r;
wire signed [`InBus]		in_24_3_i;
wire signed [`InBus]		in_24_4_r;
wire signed [`InBus]		in_24_4_i;
wire signed [`InBus]		in_24_5_r;
wire signed [`InBus]		in_24_5_i;
wire signed [`InBus]		in_24_6_r;
wire signed [`InBus]		in_24_6_i;
wire signed [`InBus]		in_24_7_r;
wire signed [`InBus]		in_24_7_i;
wire signed [`InBus]		in_24_8_r;
wire signed [`InBus]		in_24_8_i;
wire signed [`InBus]		in_24_9_r;
wire signed [`InBus]		in_24_9_i;
wire signed [`InBus]		in_24_10_r;
wire signed [`InBus]		in_24_10_i;
wire signed [`InBus]		in_24_11_r;
wire signed [`InBus]		in_24_11_i;
wire signed [`InBus]		in_24_12_r;
wire signed [`InBus]		in_24_12_i;
wire signed [`InBus]		in_24_13_r;
wire signed [`InBus]		in_24_13_i;
wire signed [`InBus]		in_24_14_r;
wire signed [`InBus]		in_24_14_i;
wire signed [`InBus]		in_24_15_r;
wire signed [`InBus]		in_24_15_i;
wire signed [`InBus]		in_24_16_r;
wire signed [`InBus]		in_24_16_i;
wire signed [`InBus]		in_24_17_r;
wire signed [`InBus]		in_24_17_i;
wire signed [`InBus]		in_24_18_r;
wire signed [`InBus]		in_24_18_i;
wire signed [`InBus]		in_24_19_r;
wire signed [`InBus]		in_24_19_i;
wire signed [`InBus]		in_24_20_r;
wire signed [`InBus]		in_24_20_i;
wire signed [`InBus]		in_24_21_r;
wire signed [`InBus]		in_24_21_i;
wire signed [`InBus]		in_24_22_r;
wire signed [`InBus]		in_24_22_i;
wire signed [`InBus]		in_24_23_r;
wire signed [`InBus]		in_24_23_i;
wire signed [`InBus]		in_24_24_r;
wire signed [`InBus]		in_24_24_i;
wire signed [`InBus]		in_24_25_r;
wire signed [`InBus]		in_24_25_i;
wire signed [`InBus]		in_24_26_r;
wire signed [`InBus]		in_24_26_i;
wire signed [`InBus]		in_24_27_r;
wire signed [`InBus]		in_24_27_i;
wire signed [`InBus]		in_24_28_r;
wire signed [`InBus]		in_24_28_i;
wire signed [`InBus]		in_24_29_r;
wire signed [`InBus]		in_24_29_i;
wire signed [`InBus]		in_24_30_r;
wire signed [`InBus]		in_24_30_i;
wire signed [`InBus]		in_24_31_r;
wire signed [`InBus]		in_24_31_i;
wire signed [`InBus]		in_24_32_r;
wire signed [`InBus]		in_24_32_i;
wire signed [`InBus]		in_25_1_r;
wire signed [`InBus]		in_25_1_i;
wire signed [`InBus]		in_25_2_r;
wire signed [`InBus]		in_25_2_i;
wire signed [`InBus]		in_25_3_r;
wire signed [`InBus]		in_25_3_i;
wire signed [`InBus]		in_25_4_r;
wire signed [`InBus]		in_25_4_i;
wire signed [`InBus]		in_25_5_r;
wire signed [`InBus]		in_25_5_i;
wire signed [`InBus]		in_25_6_r;
wire signed [`InBus]		in_25_6_i;
wire signed [`InBus]		in_25_7_r;
wire signed [`InBus]		in_25_7_i;
wire signed [`InBus]		in_25_8_r;
wire signed [`InBus]		in_25_8_i;
wire signed [`InBus]		in_25_9_r;
wire signed [`InBus]		in_25_9_i;
wire signed [`InBus]		in_25_10_r;
wire signed [`InBus]		in_25_10_i;
wire signed [`InBus]		in_25_11_r;
wire signed [`InBus]		in_25_11_i;
wire signed [`InBus]		in_25_12_r;
wire signed [`InBus]		in_25_12_i;
wire signed [`InBus]		in_25_13_r;
wire signed [`InBus]		in_25_13_i;
wire signed [`InBus]		in_25_14_r;
wire signed [`InBus]		in_25_14_i;
wire signed [`InBus]		in_25_15_r;
wire signed [`InBus]		in_25_15_i;
wire signed [`InBus]		in_25_16_r;
wire signed [`InBus]		in_25_16_i;
wire signed [`InBus]		in_25_17_r;
wire signed [`InBus]		in_25_17_i;
wire signed [`InBus]		in_25_18_r;
wire signed [`InBus]		in_25_18_i;
wire signed [`InBus]		in_25_19_r;
wire signed [`InBus]		in_25_19_i;
wire signed [`InBus]		in_25_20_r;
wire signed [`InBus]		in_25_20_i;
wire signed [`InBus]		in_25_21_r;
wire signed [`InBus]		in_25_21_i;
wire signed [`InBus]		in_25_22_r;
wire signed [`InBus]		in_25_22_i;
wire signed [`InBus]		in_25_23_r;
wire signed [`InBus]		in_25_23_i;
wire signed [`InBus]		in_25_24_r;
wire signed [`InBus]		in_25_24_i;
wire signed [`InBus]		in_25_25_r;
wire signed [`InBus]		in_25_25_i;
wire signed [`InBus]		in_25_26_r;
wire signed [`InBus]		in_25_26_i;
wire signed [`InBus]		in_25_27_r;
wire signed [`InBus]		in_25_27_i;
wire signed [`InBus]		in_25_28_r;
wire signed [`InBus]		in_25_28_i;
wire signed [`InBus]		in_25_29_r;
wire signed [`InBus]		in_25_29_i;
wire signed [`InBus]		in_25_30_r;
wire signed [`InBus]		in_25_30_i;
wire signed [`InBus]		in_25_31_r;
wire signed [`InBus]		in_25_31_i;
wire signed [`InBus]		in_25_32_r;
wire signed [`InBus]		in_25_32_i;
wire signed [`InBus]		in_26_1_r;
wire signed [`InBus]		in_26_1_i;
wire signed [`InBus]		in_26_2_r;
wire signed [`InBus]		in_26_2_i;
wire signed [`InBus]		in_26_3_r;
wire signed [`InBus]		in_26_3_i;
wire signed [`InBus]		in_26_4_r;
wire signed [`InBus]		in_26_4_i;
wire signed [`InBus]		in_26_5_r;
wire signed [`InBus]		in_26_5_i;
wire signed [`InBus]		in_26_6_r;
wire signed [`InBus]		in_26_6_i;
wire signed [`InBus]		in_26_7_r;
wire signed [`InBus]		in_26_7_i;
wire signed [`InBus]		in_26_8_r;
wire signed [`InBus]		in_26_8_i;
wire signed [`InBus]		in_26_9_r;
wire signed [`InBus]		in_26_9_i;
wire signed [`InBus]		in_26_10_r;
wire signed [`InBus]		in_26_10_i;
wire signed [`InBus]		in_26_11_r;
wire signed [`InBus]		in_26_11_i;
wire signed [`InBus]		in_26_12_r;
wire signed [`InBus]		in_26_12_i;
wire signed [`InBus]		in_26_13_r;
wire signed [`InBus]		in_26_13_i;
wire signed [`InBus]		in_26_14_r;
wire signed [`InBus]		in_26_14_i;
wire signed [`InBus]		in_26_15_r;
wire signed [`InBus]		in_26_15_i;
wire signed [`InBus]		in_26_16_r;
wire signed [`InBus]		in_26_16_i;
wire signed [`InBus]		in_26_17_r;
wire signed [`InBus]		in_26_17_i;
wire signed [`InBus]		in_26_18_r;
wire signed [`InBus]		in_26_18_i;
wire signed [`InBus]		in_26_19_r;
wire signed [`InBus]		in_26_19_i;
wire signed [`InBus]		in_26_20_r;
wire signed [`InBus]		in_26_20_i;
wire signed [`InBus]		in_26_21_r;
wire signed [`InBus]		in_26_21_i;
wire signed [`InBus]		in_26_22_r;
wire signed [`InBus]		in_26_22_i;
wire signed [`InBus]		in_26_23_r;
wire signed [`InBus]		in_26_23_i;
wire signed [`InBus]		in_26_24_r;
wire signed [`InBus]		in_26_24_i;
wire signed [`InBus]		in_26_25_r;
wire signed [`InBus]		in_26_25_i;
wire signed [`InBus]		in_26_26_r;
wire signed [`InBus]		in_26_26_i;
wire signed [`InBus]		in_26_27_r;
wire signed [`InBus]		in_26_27_i;
wire signed [`InBus]		in_26_28_r;
wire signed [`InBus]		in_26_28_i;
wire signed [`InBus]		in_26_29_r;
wire signed [`InBus]		in_26_29_i;
wire signed [`InBus]		in_26_30_r;
wire signed [`InBus]		in_26_30_i;
wire signed [`InBus]		in_26_31_r;
wire signed [`InBus]		in_26_31_i;
wire signed [`InBus]		in_26_32_r;
wire signed [`InBus]		in_26_32_i;
wire signed [`InBus]		in_27_1_r;
wire signed [`InBus]		in_27_1_i;
wire signed [`InBus]		in_27_2_r;
wire signed [`InBus]		in_27_2_i;
wire signed [`InBus]		in_27_3_r;
wire signed [`InBus]		in_27_3_i;
wire signed [`InBus]		in_27_4_r;
wire signed [`InBus]		in_27_4_i;
wire signed [`InBus]		in_27_5_r;
wire signed [`InBus]		in_27_5_i;
wire signed [`InBus]		in_27_6_r;
wire signed [`InBus]		in_27_6_i;
wire signed [`InBus]		in_27_7_r;
wire signed [`InBus]		in_27_7_i;
wire signed [`InBus]		in_27_8_r;
wire signed [`InBus]		in_27_8_i;
wire signed [`InBus]		in_27_9_r;
wire signed [`InBus]		in_27_9_i;
wire signed [`InBus]		in_27_10_r;
wire signed [`InBus]		in_27_10_i;
wire signed [`InBus]		in_27_11_r;
wire signed [`InBus]		in_27_11_i;
wire signed [`InBus]		in_27_12_r;
wire signed [`InBus]		in_27_12_i;
wire signed [`InBus]		in_27_13_r;
wire signed [`InBus]		in_27_13_i;
wire signed [`InBus]		in_27_14_r;
wire signed [`InBus]		in_27_14_i;
wire signed [`InBus]		in_27_15_r;
wire signed [`InBus]		in_27_15_i;
wire signed [`InBus]		in_27_16_r;
wire signed [`InBus]		in_27_16_i;
wire signed [`InBus]		in_27_17_r;
wire signed [`InBus]		in_27_17_i;
wire signed [`InBus]		in_27_18_r;
wire signed [`InBus]		in_27_18_i;
wire signed [`InBus]		in_27_19_r;
wire signed [`InBus]		in_27_19_i;
wire signed [`InBus]		in_27_20_r;
wire signed [`InBus]		in_27_20_i;
wire signed [`InBus]		in_27_21_r;
wire signed [`InBus]		in_27_21_i;
wire signed [`InBus]		in_27_22_r;
wire signed [`InBus]		in_27_22_i;
wire signed [`InBus]		in_27_23_r;
wire signed [`InBus]		in_27_23_i;
wire signed [`InBus]		in_27_24_r;
wire signed [`InBus]		in_27_24_i;
wire signed [`InBus]		in_27_25_r;
wire signed [`InBus]		in_27_25_i;
wire signed [`InBus]		in_27_26_r;
wire signed [`InBus]		in_27_26_i;
wire signed [`InBus]		in_27_27_r;
wire signed [`InBus]		in_27_27_i;
wire signed [`InBus]		in_27_28_r;
wire signed [`InBus]		in_27_28_i;
wire signed [`InBus]		in_27_29_r;
wire signed [`InBus]		in_27_29_i;
wire signed [`InBus]		in_27_30_r;
wire signed [`InBus]		in_27_30_i;
wire signed [`InBus]		in_27_31_r;
wire signed [`InBus]		in_27_31_i;
wire signed [`InBus]		in_27_32_r;
wire signed [`InBus]		in_27_32_i;
wire signed [`InBus]		in_28_1_r;
wire signed [`InBus]		in_28_1_i;
wire signed [`InBus]		in_28_2_r;
wire signed [`InBus]		in_28_2_i;
wire signed [`InBus]		in_28_3_r;
wire signed [`InBus]		in_28_3_i;
wire signed [`InBus]		in_28_4_r;
wire signed [`InBus]		in_28_4_i;
wire signed [`InBus]		in_28_5_r;
wire signed [`InBus]		in_28_5_i;
wire signed [`InBus]		in_28_6_r;
wire signed [`InBus]		in_28_6_i;
wire signed [`InBus]		in_28_7_r;
wire signed [`InBus]		in_28_7_i;
wire signed [`InBus]		in_28_8_r;
wire signed [`InBus]		in_28_8_i;
wire signed [`InBus]		in_28_9_r;
wire signed [`InBus]		in_28_9_i;
wire signed [`InBus]		in_28_10_r;
wire signed [`InBus]		in_28_10_i;
wire signed [`InBus]		in_28_11_r;
wire signed [`InBus]		in_28_11_i;
wire signed [`InBus]		in_28_12_r;
wire signed [`InBus]		in_28_12_i;
wire signed [`InBus]		in_28_13_r;
wire signed [`InBus]		in_28_13_i;
wire signed [`InBus]		in_28_14_r;
wire signed [`InBus]		in_28_14_i;
wire signed [`InBus]		in_28_15_r;
wire signed [`InBus]		in_28_15_i;
wire signed [`InBus]		in_28_16_r;
wire signed [`InBus]		in_28_16_i;
wire signed [`InBus]		in_28_17_r;
wire signed [`InBus]		in_28_17_i;
wire signed [`InBus]		in_28_18_r;
wire signed [`InBus]		in_28_18_i;
wire signed [`InBus]		in_28_19_r;
wire signed [`InBus]		in_28_19_i;
wire signed [`InBus]		in_28_20_r;
wire signed [`InBus]		in_28_20_i;
wire signed [`InBus]		in_28_21_r;
wire signed [`InBus]		in_28_21_i;
wire signed [`InBus]		in_28_22_r;
wire signed [`InBus]		in_28_22_i;
wire signed [`InBus]		in_28_23_r;
wire signed [`InBus]		in_28_23_i;
wire signed [`InBus]		in_28_24_r;
wire signed [`InBus]		in_28_24_i;
wire signed [`InBus]		in_28_25_r;
wire signed [`InBus]		in_28_25_i;
wire signed [`InBus]		in_28_26_r;
wire signed [`InBus]		in_28_26_i;
wire signed [`InBus]		in_28_27_r;
wire signed [`InBus]		in_28_27_i;
wire signed [`InBus]		in_28_28_r;
wire signed [`InBus]		in_28_28_i;
wire signed [`InBus]		in_28_29_r;
wire signed [`InBus]		in_28_29_i;
wire signed [`InBus]		in_28_30_r;
wire signed [`InBus]		in_28_30_i;
wire signed [`InBus]		in_28_31_r;
wire signed [`InBus]		in_28_31_i;
wire signed [`InBus]		in_28_32_r;
wire signed [`InBus]		in_28_32_i;
wire signed [`InBus]		in_29_1_r;
wire signed [`InBus]		in_29_1_i;
wire signed [`InBus]		in_29_2_r;
wire signed [`InBus]		in_29_2_i;
wire signed [`InBus]		in_29_3_r;
wire signed [`InBus]		in_29_3_i;
wire signed [`InBus]		in_29_4_r;
wire signed [`InBus]		in_29_4_i;
wire signed [`InBus]		in_29_5_r;
wire signed [`InBus]		in_29_5_i;
wire signed [`InBus]		in_29_6_r;
wire signed [`InBus]		in_29_6_i;
wire signed [`InBus]		in_29_7_r;
wire signed [`InBus]		in_29_7_i;
wire signed [`InBus]		in_29_8_r;
wire signed [`InBus]		in_29_8_i;
wire signed [`InBus]		in_29_9_r;
wire signed [`InBus]		in_29_9_i;
wire signed [`InBus]		in_29_10_r;
wire signed [`InBus]		in_29_10_i;
wire signed [`InBus]		in_29_11_r;
wire signed [`InBus]		in_29_11_i;
wire signed [`InBus]		in_29_12_r;
wire signed [`InBus]		in_29_12_i;
wire signed [`InBus]		in_29_13_r;
wire signed [`InBus]		in_29_13_i;
wire signed [`InBus]		in_29_14_r;
wire signed [`InBus]		in_29_14_i;
wire signed [`InBus]		in_29_15_r;
wire signed [`InBus]		in_29_15_i;
wire signed [`InBus]		in_29_16_r;
wire signed [`InBus]		in_29_16_i;
wire signed [`InBus]		in_29_17_r;
wire signed [`InBus]		in_29_17_i;
wire signed [`InBus]		in_29_18_r;
wire signed [`InBus]		in_29_18_i;
wire signed [`InBus]		in_29_19_r;
wire signed [`InBus]		in_29_19_i;
wire signed [`InBus]		in_29_20_r;
wire signed [`InBus]		in_29_20_i;
wire signed [`InBus]		in_29_21_r;
wire signed [`InBus]		in_29_21_i;
wire signed [`InBus]		in_29_22_r;
wire signed [`InBus]		in_29_22_i;
wire signed [`InBus]		in_29_23_r;
wire signed [`InBus]		in_29_23_i;
wire signed [`InBus]		in_29_24_r;
wire signed [`InBus]		in_29_24_i;
wire signed [`InBus]		in_29_25_r;
wire signed [`InBus]		in_29_25_i;
wire signed [`InBus]		in_29_26_r;
wire signed [`InBus]		in_29_26_i;
wire signed [`InBus]		in_29_27_r;
wire signed [`InBus]		in_29_27_i;
wire signed [`InBus]		in_29_28_r;
wire signed [`InBus]		in_29_28_i;
wire signed [`InBus]		in_29_29_r;
wire signed [`InBus]		in_29_29_i;
wire signed [`InBus]		in_29_30_r;
wire signed [`InBus]		in_29_30_i;
wire signed [`InBus]		in_29_31_r;
wire signed [`InBus]		in_29_31_i;
wire signed [`InBus]		in_29_32_r;
wire signed [`InBus]		in_29_32_i;
wire signed [`InBus]		in_30_1_r;
wire signed [`InBus]		in_30_1_i;
wire signed [`InBus]		in_30_2_r;
wire signed [`InBus]		in_30_2_i;
wire signed [`InBus]		in_30_3_r;
wire signed [`InBus]		in_30_3_i;
wire signed [`InBus]		in_30_4_r;
wire signed [`InBus]		in_30_4_i;
wire signed [`InBus]		in_30_5_r;
wire signed [`InBus]		in_30_5_i;
wire signed [`InBus]		in_30_6_r;
wire signed [`InBus]		in_30_6_i;
wire signed [`InBus]		in_30_7_r;
wire signed [`InBus]		in_30_7_i;
wire signed [`InBus]		in_30_8_r;
wire signed [`InBus]		in_30_8_i;
wire signed [`InBus]		in_30_9_r;
wire signed [`InBus]		in_30_9_i;
wire signed [`InBus]		in_30_10_r;
wire signed [`InBus]		in_30_10_i;
wire signed [`InBus]		in_30_11_r;
wire signed [`InBus]		in_30_11_i;
wire signed [`InBus]		in_30_12_r;
wire signed [`InBus]		in_30_12_i;
wire signed [`InBus]		in_30_13_r;
wire signed [`InBus]		in_30_13_i;
wire signed [`InBus]		in_30_14_r;
wire signed [`InBus]		in_30_14_i;
wire signed [`InBus]		in_30_15_r;
wire signed [`InBus]		in_30_15_i;
wire signed [`InBus]		in_30_16_r;
wire signed [`InBus]		in_30_16_i;
wire signed [`InBus]		in_30_17_r;
wire signed [`InBus]		in_30_17_i;
wire signed [`InBus]		in_30_18_r;
wire signed [`InBus]		in_30_18_i;
wire signed [`InBus]		in_30_19_r;
wire signed [`InBus]		in_30_19_i;
wire signed [`InBus]		in_30_20_r;
wire signed [`InBus]		in_30_20_i;
wire signed [`InBus]		in_30_21_r;
wire signed [`InBus]		in_30_21_i;
wire signed [`InBus]		in_30_22_r;
wire signed [`InBus]		in_30_22_i;
wire signed [`InBus]		in_30_23_r;
wire signed [`InBus]		in_30_23_i;
wire signed [`InBus]		in_30_24_r;
wire signed [`InBus]		in_30_24_i;
wire signed [`InBus]		in_30_25_r;
wire signed [`InBus]		in_30_25_i;
wire signed [`InBus]		in_30_26_r;
wire signed [`InBus]		in_30_26_i;
wire signed [`InBus]		in_30_27_r;
wire signed [`InBus]		in_30_27_i;
wire signed [`InBus]		in_30_28_r;
wire signed [`InBus]		in_30_28_i;
wire signed [`InBus]		in_30_29_r;
wire signed [`InBus]		in_30_29_i;
wire signed [`InBus]		in_30_30_r;
wire signed [`InBus]		in_30_30_i;
wire signed [`InBus]		in_30_31_r;
wire signed [`InBus]		in_30_31_i;
wire signed [`InBus]		in_30_32_r;
wire signed [`InBus]		in_30_32_i;
wire signed [`InBus]		in_31_1_r;
wire signed [`InBus]		in_31_1_i;
wire signed [`InBus]		in_31_2_r;
wire signed [`InBus]		in_31_2_i;
wire signed [`InBus]		in_31_3_r;
wire signed [`InBus]		in_31_3_i;
wire signed [`InBus]		in_31_4_r;
wire signed [`InBus]		in_31_4_i;
wire signed [`InBus]		in_31_5_r;
wire signed [`InBus]		in_31_5_i;
wire signed [`InBus]		in_31_6_r;
wire signed [`InBus]		in_31_6_i;
wire signed [`InBus]		in_31_7_r;
wire signed [`InBus]		in_31_7_i;
wire signed [`InBus]		in_31_8_r;
wire signed [`InBus]		in_31_8_i;
wire signed [`InBus]		in_31_9_r;
wire signed [`InBus]		in_31_9_i;
wire signed [`InBus]		in_31_10_r;
wire signed [`InBus]		in_31_10_i;
wire signed [`InBus]		in_31_11_r;
wire signed [`InBus]		in_31_11_i;
wire signed [`InBus]		in_31_12_r;
wire signed [`InBus]		in_31_12_i;
wire signed [`InBus]		in_31_13_r;
wire signed [`InBus]		in_31_13_i;
wire signed [`InBus]		in_31_14_r;
wire signed [`InBus]		in_31_14_i;
wire signed [`InBus]		in_31_15_r;
wire signed [`InBus]		in_31_15_i;
wire signed [`InBus]		in_31_16_r;
wire signed [`InBus]		in_31_16_i;
wire signed [`InBus]		in_31_17_r;
wire signed [`InBus]		in_31_17_i;
wire signed [`InBus]		in_31_18_r;
wire signed [`InBus]		in_31_18_i;
wire signed [`InBus]		in_31_19_r;
wire signed [`InBus]		in_31_19_i;
wire signed [`InBus]		in_31_20_r;
wire signed [`InBus]		in_31_20_i;
wire signed [`InBus]		in_31_21_r;
wire signed [`InBus]		in_31_21_i;
wire signed [`InBus]		in_31_22_r;
wire signed [`InBus]		in_31_22_i;
wire signed [`InBus]		in_31_23_r;
wire signed [`InBus]		in_31_23_i;
wire signed [`InBus]		in_31_24_r;
wire signed [`InBus]		in_31_24_i;
wire signed [`InBus]		in_31_25_r;
wire signed [`InBus]		in_31_25_i;
wire signed [`InBus]		in_31_26_r;
wire signed [`InBus]		in_31_26_i;
wire signed [`InBus]		in_31_27_r;
wire signed [`InBus]		in_31_27_i;
wire signed [`InBus]		in_31_28_r;
wire signed [`InBus]		in_31_28_i;
wire signed [`InBus]		in_31_29_r;
wire signed [`InBus]		in_31_29_i;
wire signed [`InBus]		in_31_30_r;
wire signed [`InBus]		in_31_30_i;
wire signed [`InBus]		in_31_31_r;
wire signed [`InBus]		in_31_31_i;
wire signed [`InBus]		in_31_32_r;
wire signed [`InBus]		in_31_32_i;
wire signed [`InBus]		in_32_1_r;
wire signed [`InBus]		in_32_1_i;
wire signed [`InBus]		in_32_2_r;
wire signed [`InBus]		in_32_2_i;
wire signed [`InBus]		in_32_3_r;
wire signed [`InBus]		in_32_3_i;
wire signed [`InBus]		in_32_4_r;
wire signed [`InBus]		in_32_4_i;
wire signed [`InBus]		in_32_5_r;
wire signed [`InBus]		in_32_5_i;
wire signed [`InBus]		in_32_6_r;
wire signed [`InBus]		in_32_6_i;
wire signed [`InBus]		in_32_7_r;
wire signed [`InBus]		in_32_7_i;
wire signed [`InBus]		in_32_8_r;
wire signed [`InBus]		in_32_8_i;
wire signed [`InBus]		in_32_9_r;
wire signed [`InBus]		in_32_9_i;
wire signed [`InBus]		in_32_10_r;
wire signed [`InBus]		in_32_10_i;
wire signed [`InBus]		in_32_11_r;
wire signed [`InBus]		in_32_11_i;
wire signed [`InBus]		in_32_12_r;
wire signed [`InBus]		in_32_12_i;
wire signed [`InBus]		in_32_13_r;
wire signed [`InBus]		in_32_13_i;
wire signed [`InBus]		in_32_14_r;
wire signed [`InBus]		in_32_14_i;
wire signed [`InBus]		in_32_15_r;
wire signed [`InBus]		in_32_15_i;
wire signed [`InBus]		in_32_16_r;
wire signed [`InBus]		in_32_16_i;
wire signed [`InBus]		in_32_17_r;
wire signed [`InBus]		in_32_17_i;
wire signed [`InBus]		in_32_18_r;
wire signed [`InBus]		in_32_18_i;
wire signed [`InBus]		in_32_19_r;
wire signed [`InBus]		in_32_19_i;
wire signed [`InBus]		in_32_20_r;
wire signed [`InBus]		in_32_20_i;
wire signed [`InBus]		in_32_21_r;
wire signed [`InBus]		in_32_21_i;
wire signed [`InBus]		in_32_22_r;
wire signed [`InBus]		in_32_22_i;
wire signed [`InBus]		in_32_23_r;
wire signed [`InBus]		in_32_23_i;
wire signed [`InBus]		in_32_24_r;
wire signed [`InBus]		in_32_24_i;
wire signed [`InBus]		in_32_25_r;
wire signed [`InBus]		in_32_25_i;
wire signed [`InBus]		in_32_26_r;
wire signed [`InBus]		in_32_26_i;
wire signed [`InBus]		in_32_27_r;
wire signed [`InBus]		in_32_27_i;
wire signed [`InBus]		in_32_28_r;
wire signed [`InBus]		in_32_28_i;
wire signed [`InBus]		in_32_29_r;
wire signed [`InBus]		in_32_29_i;
wire signed [`InBus]		in_32_30_r;
wire signed [`InBus]		in_32_30_i;
wire signed [`InBus]		in_32_31_r;
wire signed [`InBus]		in_32_31_i;
wire signed [`InBus]		in_32_32_r;
wire signed [`InBus]		in_32_32_i;

wire signed [`OutBus]		out_1_1_r;
wire signed [`OutBus]		out_1_1_i;
wire signed [`OutBus]		out_1_2_r;
wire signed [`OutBus]		out_1_2_i;
wire signed [`OutBus]		out_1_3_r;
wire signed [`OutBus]		out_1_3_i;
wire signed [`OutBus]		out_1_4_r;
wire signed [`OutBus]		out_1_4_i;
wire signed [`OutBus]		out_1_5_r;
wire signed [`OutBus]		out_1_5_i;
wire signed [`OutBus]		out_1_6_r;
wire signed [`OutBus]		out_1_6_i;
wire signed [`OutBus]		out_1_7_r;
wire signed [`OutBus]		out_1_7_i;
wire signed [`OutBus]		out_1_8_r;
wire signed [`OutBus]		out_1_8_i;
wire signed [`OutBus]		out_1_9_r;
wire signed [`OutBus]		out_1_9_i;
wire signed [`OutBus]		out_1_10_r;
wire signed [`OutBus]		out_1_10_i;
wire signed [`OutBus]		out_1_11_r;
wire signed [`OutBus]		out_1_11_i;
wire signed [`OutBus]		out_1_12_r;
wire signed [`OutBus]		out_1_12_i;
wire signed [`OutBus]		out_1_13_r;
wire signed [`OutBus]		out_1_13_i;
wire signed [`OutBus]		out_1_14_r;
wire signed [`OutBus]		out_1_14_i;
wire signed [`OutBus]		out_1_15_r;
wire signed [`OutBus]		out_1_15_i;
wire signed [`OutBus]		out_1_16_r;
wire signed [`OutBus]		out_1_16_i;
wire signed [`OutBus]		out_1_17_r;
wire signed [`OutBus]		out_1_17_i;
wire signed [`OutBus]		out_1_18_r;
wire signed [`OutBus]		out_1_18_i;
wire signed [`OutBus]		out_1_19_r;
wire signed [`OutBus]		out_1_19_i;
wire signed [`OutBus]		out_1_20_r;
wire signed [`OutBus]		out_1_20_i;
wire signed [`OutBus]		out_1_21_r;
wire signed [`OutBus]		out_1_21_i;
wire signed [`OutBus]		out_1_22_r;
wire signed [`OutBus]		out_1_22_i;
wire signed [`OutBus]		out_1_23_r;
wire signed [`OutBus]		out_1_23_i;
wire signed [`OutBus]		out_1_24_r;
wire signed [`OutBus]		out_1_24_i;
wire signed [`OutBus]		out_1_25_r;
wire signed [`OutBus]		out_1_25_i;
wire signed [`OutBus]		out_1_26_r;
wire signed [`OutBus]		out_1_26_i;
wire signed [`OutBus]		out_1_27_r;
wire signed [`OutBus]		out_1_27_i;
wire signed [`OutBus]		out_1_28_r;
wire signed [`OutBus]		out_1_28_i;
wire signed [`OutBus]		out_1_29_r;
wire signed [`OutBus]		out_1_29_i;
wire signed [`OutBus]		out_1_30_r;
wire signed [`OutBus]		out_1_30_i;
wire signed [`OutBus]		out_1_31_r;
wire signed [`OutBus]		out_1_31_i;
wire signed [`OutBus]		out_1_32_r;
wire signed [`OutBus]		out_1_32_i;
wire signed [`OutBus]		out_2_1_r;
wire signed [`OutBus]		out_2_1_i;
wire signed [`OutBus]		out_2_2_r;
wire signed [`OutBus]		out_2_2_i;
wire signed [`OutBus]		out_2_3_r;
wire signed [`OutBus]		out_2_3_i;
wire signed [`OutBus]		out_2_4_r;
wire signed [`OutBus]		out_2_4_i;
wire signed [`OutBus]		out_2_5_r;
wire signed [`OutBus]		out_2_5_i;
wire signed [`OutBus]		out_2_6_r;
wire signed [`OutBus]		out_2_6_i;
wire signed [`OutBus]		out_2_7_r;
wire signed [`OutBus]		out_2_7_i;
wire signed [`OutBus]		out_2_8_r;
wire signed [`OutBus]		out_2_8_i;
wire signed [`OutBus]		out_2_9_r;
wire signed [`OutBus]		out_2_9_i;
wire signed [`OutBus]		out_2_10_r;
wire signed [`OutBus]		out_2_10_i;
wire signed [`OutBus]		out_2_11_r;
wire signed [`OutBus]		out_2_11_i;
wire signed [`OutBus]		out_2_12_r;
wire signed [`OutBus]		out_2_12_i;
wire signed [`OutBus]		out_2_13_r;
wire signed [`OutBus]		out_2_13_i;
wire signed [`OutBus]		out_2_14_r;
wire signed [`OutBus]		out_2_14_i;
wire signed [`OutBus]		out_2_15_r;
wire signed [`OutBus]		out_2_15_i;
wire signed [`OutBus]		out_2_16_r;
wire signed [`OutBus]		out_2_16_i;
wire signed [`OutBus]		out_2_17_r;
wire signed [`OutBus]		out_2_17_i;
wire signed [`OutBus]		out_2_18_r;
wire signed [`OutBus]		out_2_18_i;
wire signed [`OutBus]		out_2_19_r;
wire signed [`OutBus]		out_2_19_i;
wire signed [`OutBus]		out_2_20_r;
wire signed [`OutBus]		out_2_20_i;
wire signed [`OutBus]		out_2_21_r;
wire signed [`OutBus]		out_2_21_i;
wire signed [`OutBus]		out_2_22_r;
wire signed [`OutBus]		out_2_22_i;
wire signed [`OutBus]		out_2_23_r;
wire signed [`OutBus]		out_2_23_i;
wire signed [`OutBus]		out_2_24_r;
wire signed [`OutBus]		out_2_24_i;
wire signed [`OutBus]		out_2_25_r;
wire signed [`OutBus]		out_2_25_i;
wire signed [`OutBus]		out_2_26_r;
wire signed [`OutBus]		out_2_26_i;
wire signed [`OutBus]		out_2_27_r;
wire signed [`OutBus]		out_2_27_i;
wire signed [`OutBus]		out_2_28_r;
wire signed [`OutBus]		out_2_28_i;
wire signed [`OutBus]		out_2_29_r;
wire signed [`OutBus]		out_2_29_i;
wire signed [`OutBus]		out_2_30_r;
wire signed [`OutBus]		out_2_30_i;
wire signed [`OutBus]		out_2_31_r;
wire signed [`OutBus]		out_2_31_i;
wire signed [`OutBus]		out_2_32_r;
wire signed [`OutBus]		out_2_32_i;
wire signed [`OutBus]		out_3_1_r;
wire signed [`OutBus]		out_3_1_i;
wire signed [`OutBus]		out_3_2_r;
wire signed [`OutBus]		out_3_2_i;
wire signed [`OutBus]		out_3_3_r;
wire signed [`OutBus]		out_3_3_i;
wire signed [`OutBus]		out_3_4_r;
wire signed [`OutBus]		out_3_4_i;
wire signed [`OutBus]		out_3_5_r;
wire signed [`OutBus]		out_3_5_i;
wire signed [`OutBus]		out_3_6_r;
wire signed [`OutBus]		out_3_6_i;
wire signed [`OutBus]		out_3_7_r;
wire signed [`OutBus]		out_3_7_i;
wire signed [`OutBus]		out_3_8_r;
wire signed [`OutBus]		out_3_8_i;
wire signed [`OutBus]		out_3_9_r;
wire signed [`OutBus]		out_3_9_i;
wire signed [`OutBus]		out_3_10_r;
wire signed [`OutBus]		out_3_10_i;
wire signed [`OutBus]		out_3_11_r;
wire signed [`OutBus]		out_3_11_i;
wire signed [`OutBus]		out_3_12_r;
wire signed [`OutBus]		out_3_12_i;
wire signed [`OutBus]		out_3_13_r;
wire signed [`OutBus]		out_3_13_i;
wire signed [`OutBus]		out_3_14_r;
wire signed [`OutBus]		out_3_14_i;
wire signed [`OutBus]		out_3_15_r;
wire signed [`OutBus]		out_3_15_i;
wire signed [`OutBus]		out_3_16_r;
wire signed [`OutBus]		out_3_16_i;
wire signed [`OutBus]		out_3_17_r;
wire signed [`OutBus]		out_3_17_i;
wire signed [`OutBus]		out_3_18_r;
wire signed [`OutBus]		out_3_18_i;
wire signed [`OutBus]		out_3_19_r;
wire signed [`OutBus]		out_3_19_i;
wire signed [`OutBus]		out_3_20_r;
wire signed [`OutBus]		out_3_20_i;
wire signed [`OutBus]		out_3_21_r;
wire signed [`OutBus]		out_3_21_i;
wire signed [`OutBus]		out_3_22_r;
wire signed [`OutBus]		out_3_22_i;
wire signed [`OutBus]		out_3_23_r;
wire signed [`OutBus]		out_3_23_i;
wire signed [`OutBus]		out_3_24_r;
wire signed [`OutBus]		out_3_24_i;
wire signed [`OutBus]		out_3_25_r;
wire signed [`OutBus]		out_3_25_i;
wire signed [`OutBus]		out_3_26_r;
wire signed [`OutBus]		out_3_26_i;
wire signed [`OutBus]		out_3_27_r;
wire signed [`OutBus]		out_3_27_i;
wire signed [`OutBus]		out_3_28_r;
wire signed [`OutBus]		out_3_28_i;
wire signed [`OutBus]		out_3_29_r;
wire signed [`OutBus]		out_3_29_i;
wire signed [`OutBus]		out_3_30_r;
wire signed [`OutBus]		out_3_30_i;
wire signed [`OutBus]		out_3_31_r;
wire signed [`OutBus]		out_3_31_i;
wire signed [`OutBus]		out_3_32_r;
wire signed [`OutBus]		out_3_32_i;
wire signed [`OutBus]		out_4_1_r;
wire signed [`OutBus]		out_4_1_i;
wire signed [`OutBus]		out_4_2_r;
wire signed [`OutBus]		out_4_2_i;
wire signed [`OutBus]		out_4_3_r;
wire signed [`OutBus]		out_4_3_i;
wire signed [`OutBus]		out_4_4_r;
wire signed [`OutBus]		out_4_4_i;
wire signed [`OutBus]		out_4_5_r;
wire signed [`OutBus]		out_4_5_i;
wire signed [`OutBus]		out_4_6_r;
wire signed [`OutBus]		out_4_6_i;
wire signed [`OutBus]		out_4_7_r;
wire signed [`OutBus]		out_4_7_i;
wire signed [`OutBus]		out_4_8_r;
wire signed [`OutBus]		out_4_8_i;
wire signed [`OutBus]		out_4_9_r;
wire signed [`OutBus]		out_4_9_i;
wire signed [`OutBus]		out_4_10_r;
wire signed [`OutBus]		out_4_10_i;
wire signed [`OutBus]		out_4_11_r;
wire signed [`OutBus]		out_4_11_i;
wire signed [`OutBus]		out_4_12_r;
wire signed [`OutBus]		out_4_12_i;
wire signed [`OutBus]		out_4_13_r;
wire signed [`OutBus]		out_4_13_i;
wire signed [`OutBus]		out_4_14_r;
wire signed [`OutBus]		out_4_14_i;
wire signed [`OutBus]		out_4_15_r;
wire signed [`OutBus]		out_4_15_i;
wire signed [`OutBus]		out_4_16_r;
wire signed [`OutBus]		out_4_16_i;
wire signed [`OutBus]		out_4_17_r;
wire signed [`OutBus]		out_4_17_i;
wire signed [`OutBus]		out_4_18_r;
wire signed [`OutBus]		out_4_18_i;
wire signed [`OutBus]		out_4_19_r;
wire signed [`OutBus]		out_4_19_i;
wire signed [`OutBus]		out_4_20_r;
wire signed [`OutBus]		out_4_20_i;
wire signed [`OutBus]		out_4_21_r;
wire signed [`OutBus]		out_4_21_i;
wire signed [`OutBus]		out_4_22_r;
wire signed [`OutBus]		out_4_22_i;
wire signed [`OutBus]		out_4_23_r;
wire signed [`OutBus]		out_4_23_i;
wire signed [`OutBus]		out_4_24_r;
wire signed [`OutBus]		out_4_24_i;
wire signed [`OutBus]		out_4_25_r;
wire signed [`OutBus]		out_4_25_i;
wire signed [`OutBus]		out_4_26_r;
wire signed [`OutBus]		out_4_26_i;
wire signed [`OutBus]		out_4_27_r;
wire signed [`OutBus]		out_4_27_i;
wire signed [`OutBus]		out_4_28_r;
wire signed [`OutBus]		out_4_28_i;
wire signed [`OutBus]		out_4_29_r;
wire signed [`OutBus]		out_4_29_i;
wire signed [`OutBus]		out_4_30_r;
wire signed [`OutBus]		out_4_30_i;
wire signed [`OutBus]		out_4_31_r;
wire signed [`OutBus]		out_4_31_i;
wire signed [`OutBus]		out_4_32_r;
wire signed [`OutBus]		out_4_32_i;
wire signed [`OutBus]		out_5_1_r;
wire signed [`OutBus]		out_5_1_i;
wire signed [`OutBus]		out_5_2_r;
wire signed [`OutBus]		out_5_2_i;
wire signed [`OutBus]		out_5_3_r;
wire signed [`OutBus]		out_5_3_i;
wire signed [`OutBus]		out_5_4_r;
wire signed [`OutBus]		out_5_4_i;
wire signed [`OutBus]		out_5_5_r;
wire signed [`OutBus]		out_5_5_i;
wire signed [`OutBus]		out_5_6_r;
wire signed [`OutBus]		out_5_6_i;
wire signed [`OutBus]		out_5_7_r;
wire signed [`OutBus]		out_5_7_i;
wire signed [`OutBus]		out_5_8_r;
wire signed [`OutBus]		out_5_8_i;
wire signed [`OutBus]		out_5_9_r;
wire signed [`OutBus]		out_5_9_i;
wire signed [`OutBus]		out_5_10_r;
wire signed [`OutBus]		out_5_10_i;
wire signed [`OutBus]		out_5_11_r;
wire signed [`OutBus]		out_5_11_i;
wire signed [`OutBus]		out_5_12_r;
wire signed [`OutBus]		out_5_12_i;
wire signed [`OutBus]		out_5_13_r;
wire signed [`OutBus]		out_5_13_i;
wire signed [`OutBus]		out_5_14_r;
wire signed [`OutBus]		out_5_14_i;
wire signed [`OutBus]		out_5_15_r;
wire signed [`OutBus]		out_5_15_i;
wire signed [`OutBus]		out_5_16_r;
wire signed [`OutBus]		out_5_16_i;
wire signed [`OutBus]		out_5_17_r;
wire signed [`OutBus]		out_5_17_i;
wire signed [`OutBus]		out_5_18_r;
wire signed [`OutBus]		out_5_18_i;
wire signed [`OutBus]		out_5_19_r;
wire signed [`OutBus]		out_5_19_i;
wire signed [`OutBus]		out_5_20_r;
wire signed [`OutBus]		out_5_20_i;
wire signed [`OutBus]		out_5_21_r;
wire signed [`OutBus]		out_5_21_i;
wire signed [`OutBus]		out_5_22_r;
wire signed [`OutBus]		out_5_22_i;
wire signed [`OutBus]		out_5_23_r;
wire signed [`OutBus]		out_5_23_i;
wire signed [`OutBus]		out_5_24_r;
wire signed [`OutBus]		out_5_24_i;
wire signed [`OutBus]		out_5_25_r;
wire signed [`OutBus]		out_5_25_i;
wire signed [`OutBus]		out_5_26_r;
wire signed [`OutBus]		out_5_26_i;
wire signed [`OutBus]		out_5_27_r;
wire signed [`OutBus]		out_5_27_i;
wire signed [`OutBus]		out_5_28_r;
wire signed [`OutBus]		out_5_28_i;
wire signed [`OutBus]		out_5_29_r;
wire signed [`OutBus]		out_5_29_i;
wire signed [`OutBus]		out_5_30_r;
wire signed [`OutBus]		out_5_30_i;
wire signed [`OutBus]		out_5_31_r;
wire signed [`OutBus]		out_5_31_i;
wire signed [`OutBus]		out_5_32_r;
wire signed [`OutBus]		out_5_32_i;
wire signed [`OutBus]		out_6_1_r;
wire signed [`OutBus]		out_6_1_i;
wire signed [`OutBus]		out_6_2_r;
wire signed [`OutBus]		out_6_2_i;
wire signed [`OutBus]		out_6_3_r;
wire signed [`OutBus]		out_6_3_i;
wire signed [`OutBus]		out_6_4_r;
wire signed [`OutBus]		out_6_4_i;
wire signed [`OutBus]		out_6_5_r;
wire signed [`OutBus]		out_6_5_i;
wire signed [`OutBus]		out_6_6_r;
wire signed [`OutBus]		out_6_6_i;
wire signed [`OutBus]		out_6_7_r;
wire signed [`OutBus]		out_6_7_i;
wire signed [`OutBus]		out_6_8_r;
wire signed [`OutBus]		out_6_8_i;
wire signed [`OutBus]		out_6_9_r;
wire signed [`OutBus]		out_6_9_i;
wire signed [`OutBus]		out_6_10_r;
wire signed [`OutBus]		out_6_10_i;
wire signed [`OutBus]		out_6_11_r;
wire signed [`OutBus]		out_6_11_i;
wire signed [`OutBus]		out_6_12_r;
wire signed [`OutBus]		out_6_12_i;
wire signed [`OutBus]		out_6_13_r;
wire signed [`OutBus]		out_6_13_i;
wire signed [`OutBus]		out_6_14_r;
wire signed [`OutBus]		out_6_14_i;
wire signed [`OutBus]		out_6_15_r;
wire signed [`OutBus]		out_6_15_i;
wire signed [`OutBus]		out_6_16_r;
wire signed [`OutBus]		out_6_16_i;
wire signed [`OutBus]		out_6_17_r;
wire signed [`OutBus]		out_6_17_i;
wire signed [`OutBus]		out_6_18_r;
wire signed [`OutBus]		out_6_18_i;
wire signed [`OutBus]		out_6_19_r;
wire signed [`OutBus]		out_6_19_i;
wire signed [`OutBus]		out_6_20_r;
wire signed [`OutBus]		out_6_20_i;
wire signed [`OutBus]		out_6_21_r;
wire signed [`OutBus]		out_6_21_i;
wire signed [`OutBus]		out_6_22_r;
wire signed [`OutBus]		out_6_22_i;
wire signed [`OutBus]		out_6_23_r;
wire signed [`OutBus]		out_6_23_i;
wire signed [`OutBus]		out_6_24_r;
wire signed [`OutBus]		out_6_24_i;
wire signed [`OutBus]		out_6_25_r;
wire signed [`OutBus]		out_6_25_i;
wire signed [`OutBus]		out_6_26_r;
wire signed [`OutBus]		out_6_26_i;
wire signed [`OutBus]		out_6_27_r;
wire signed [`OutBus]		out_6_27_i;
wire signed [`OutBus]		out_6_28_r;
wire signed [`OutBus]		out_6_28_i;
wire signed [`OutBus]		out_6_29_r;
wire signed [`OutBus]		out_6_29_i;
wire signed [`OutBus]		out_6_30_r;
wire signed [`OutBus]		out_6_30_i;
wire signed [`OutBus]		out_6_31_r;
wire signed [`OutBus]		out_6_31_i;
wire signed [`OutBus]		out_6_32_r;
wire signed [`OutBus]		out_6_32_i;
wire signed [`OutBus]		out_7_1_r;
wire signed [`OutBus]		out_7_1_i;
wire signed [`OutBus]		out_7_2_r;
wire signed [`OutBus]		out_7_2_i;
wire signed [`OutBus]		out_7_3_r;
wire signed [`OutBus]		out_7_3_i;
wire signed [`OutBus]		out_7_4_r;
wire signed [`OutBus]		out_7_4_i;
wire signed [`OutBus]		out_7_5_r;
wire signed [`OutBus]		out_7_5_i;
wire signed [`OutBus]		out_7_6_r;
wire signed [`OutBus]		out_7_6_i;
wire signed [`OutBus]		out_7_7_r;
wire signed [`OutBus]		out_7_7_i;
wire signed [`OutBus]		out_7_8_r;
wire signed [`OutBus]		out_7_8_i;
wire signed [`OutBus]		out_7_9_r;
wire signed [`OutBus]		out_7_9_i;
wire signed [`OutBus]		out_7_10_r;
wire signed [`OutBus]		out_7_10_i;
wire signed [`OutBus]		out_7_11_r;
wire signed [`OutBus]		out_7_11_i;
wire signed [`OutBus]		out_7_12_r;
wire signed [`OutBus]		out_7_12_i;
wire signed [`OutBus]		out_7_13_r;
wire signed [`OutBus]		out_7_13_i;
wire signed [`OutBus]		out_7_14_r;
wire signed [`OutBus]		out_7_14_i;
wire signed [`OutBus]		out_7_15_r;
wire signed [`OutBus]		out_7_15_i;
wire signed [`OutBus]		out_7_16_r;
wire signed [`OutBus]		out_7_16_i;
wire signed [`OutBus]		out_7_17_r;
wire signed [`OutBus]		out_7_17_i;
wire signed [`OutBus]		out_7_18_r;
wire signed [`OutBus]		out_7_18_i;
wire signed [`OutBus]		out_7_19_r;
wire signed [`OutBus]		out_7_19_i;
wire signed [`OutBus]		out_7_20_r;
wire signed [`OutBus]		out_7_20_i;
wire signed [`OutBus]		out_7_21_r;
wire signed [`OutBus]		out_7_21_i;
wire signed [`OutBus]		out_7_22_r;
wire signed [`OutBus]		out_7_22_i;
wire signed [`OutBus]		out_7_23_r;
wire signed [`OutBus]		out_7_23_i;
wire signed [`OutBus]		out_7_24_r;
wire signed [`OutBus]		out_7_24_i;
wire signed [`OutBus]		out_7_25_r;
wire signed [`OutBus]		out_7_25_i;
wire signed [`OutBus]		out_7_26_r;
wire signed [`OutBus]		out_7_26_i;
wire signed [`OutBus]		out_7_27_r;
wire signed [`OutBus]		out_7_27_i;
wire signed [`OutBus]		out_7_28_r;
wire signed [`OutBus]		out_7_28_i;
wire signed [`OutBus]		out_7_29_r;
wire signed [`OutBus]		out_7_29_i;
wire signed [`OutBus]		out_7_30_r;
wire signed [`OutBus]		out_7_30_i;
wire signed [`OutBus]		out_7_31_r;
wire signed [`OutBus]		out_7_31_i;
wire signed [`OutBus]		out_7_32_r;
wire signed [`OutBus]		out_7_32_i;
wire signed [`OutBus]		out_8_1_r;
wire signed [`OutBus]		out_8_1_i;
wire signed [`OutBus]		out_8_2_r;
wire signed [`OutBus]		out_8_2_i;
wire signed [`OutBus]		out_8_3_r;
wire signed [`OutBus]		out_8_3_i;
wire signed [`OutBus]		out_8_4_r;
wire signed [`OutBus]		out_8_4_i;
wire signed [`OutBus]		out_8_5_r;
wire signed [`OutBus]		out_8_5_i;
wire signed [`OutBus]		out_8_6_r;
wire signed [`OutBus]		out_8_6_i;
wire signed [`OutBus]		out_8_7_r;
wire signed [`OutBus]		out_8_7_i;
wire signed [`OutBus]		out_8_8_r;
wire signed [`OutBus]		out_8_8_i;
wire signed [`OutBus]		out_8_9_r;
wire signed [`OutBus]		out_8_9_i;
wire signed [`OutBus]		out_8_10_r;
wire signed [`OutBus]		out_8_10_i;
wire signed [`OutBus]		out_8_11_r;
wire signed [`OutBus]		out_8_11_i;
wire signed [`OutBus]		out_8_12_r;
wire signed [`OutBus]		out_8_12_i;
wire signed [`OutBus]		out_8_13_r;
wire signed [`OutBus]		out_8_13_i;
wire signed [`OutBus]		out_8_14_r;
wire signed [`OutBus]		out_8_14_i;
wire signed [`OutBus]		out_8_15_r;
wire signed [`OutBus]		out_8_15_i;
wire signed [`OutBus]		out_8_16_r;
wire signed [`OutBus]		out_8_16_i;
wire signed [`OutBus]		out_8_17_r;
wire signed [`OutBus]		out_8_17_i;
wire signed [`OutBus]		out_8_18_r;
wire signed [`OutBus]		out_8_18_i;
wire signed [`OutBus]		out_8_19_r;
wire signed [`OutBus]		out_8_19_i;
wire signed [`OutBus]		out_8_20_r;
wire signed [`OutBus]		out_8_20_i;
wire signed [`OutBus]		out_8_21_r;
wire signed [`OutBus]		out_8_21_i;
wire signed [`OutBus]		out_8_22_r;
wire signed [`OutBus]		out_8_22_i;
wire signed [`OutBus]		out_8_23_r;
wire signed [`OutBus]		out_8_23_i;
wire signed [`OutBus]		out_8_24_r;
wire signed [`OutBus]		out_8_24_i;
wire signed [`OutBus]		out_8_25_r;
wire signed [`OutBus]		out_8_25_i;
wire signed [`OutBus]		out_8_26_r;
wire signed [`OutBus]		out_8_26_i;
wire signed [`OutBus]		out_8_27_r;
wire signed [`OutBus]		out_8_27_i;
wire signed [`OutBus]		out_8_28_r;
wire signed [`OutBus]		out_8_28_i;
wire signed [`OutBus]		out_8_29_r;
wire signed [`OutBus]		out_8_29_i;
wire signed [`OutBus]		out_8_30_r;
wire signed [`OutBus]		out_8_30_i;
wire signed [`OutBus]		out_8_31_r;
wire signed [`OutBus]		out_8_31_i;
wire signed [`OutBus]		out_8_32_r;
wire signed [`OutBus]		out_8_32_i;
wire signed [`OutBus]		out_9_1_r;
wire signed [`OutBus]		out_9_1_i;
wire signed [`OutBus]		out_9_2_r;
wire signed [`OutBus]		out_9_2_i;
wire signed [`OutBus]		out_9_3_r;
wire signed [`OutBus]		out_9_3_i;
wire signed [`OutBus]		out_9_4_r;
wire signed [`OutBus]		out_9_4_i;
wire signed [`OutBus]		out_9_5_r;
wire signed [`OutBus]		out_9_5_i;
wire signed [`OutBus]		out_9_6_r;
wire signed [`OutBus]		out_9_6_i;
wire signed [`OutBus]		out_9_7_r;
wire signed [`OutBus]		out_9_7_i;
wire signed [`OutBus]		out_9_8_r;
wire signed [`OutBus]		out_9_8_i;
wire signed [`OutBus]		out_9_9_r;
wire signed [`OutBus]		out_9_9_i;
wire signed [`OutBus]		out_9_10_r;
wire signed [`OutBus]		out_9_10_i;
wire signed [`OutBus]		out_9_11_r;
wire signed [`OutBus]		out_9_11_i;
wire signed [`OutBus]		out_9_12_r;
wire signed [`OutBus]		out_9_12_i;
wire signed [`OutBus]		out_9_13_r;
wire signed [`OutBus]		out_9_13_i;
wire signed [`OutBus]		out_9_14_r;
wire signed [`OutBus]		out_9_14_i;
wire signed [`OutBus]		out_9_15_r;
wire signed [`OutBus]		out_9_15_i;
wire signed [`OutBus]		out_9_16_r;
wire signed [`OutBus]		out_9_16_i;
wire signed [`OutBus]		out_9_17_r;
wire signed [`OutBus]		out_9_17_i;
wire signed [`OutBus]		out_9_18_r;
wire signed [`OutBus]		out_9_18_i;
wire signed [`OutBus]		out_9_19_r;
wire signed [`OutBus]		out_9_19_i;
wire signed [`OutBus]		out_9_20_r;
wire signed [`OutBus]		out_9_20_i;
wire signed [`OutBus]		out_9_21_r;
wire signed [`OutBus]		out_9_21_i;
wire signed [`OutBus]		out_9_22_r;
wire signed [`OutBus]		out_9_22_i;
wire signed [`OutBus]		out_9_23_r;
wire signed [`OutBus]		out_9_23_i;
wire signed [`OutBus]		out_9_24_r;
wire signed [`OutBus]		out_9_24_i;
wire signed [`OutBus]		out_9_25_r;
wire signed [`OutBus]		out_9_25_i;
wire signed [`OutBus]		out_9_26_r;
wire signed [`OutBus]		out_9_26_i;
wire signed [`OutBus]		out_9_27_r;
wire signed [`OutBus]		out_9_27_i;
wire signed [`OutBus]		out_9_28_r;
wire signed [`OutBus]		out_9_28_i;
wire signed [`OutBus]		out_9_29_r;
wire signed [`OutBus]		out_9_29_i;
wire signed [`OutBus]		out_9_30_r;
wire signed [`OutBus]		out_9_30_i;
wire signed [`OutBus]		out_9_31_r;
wire signed [`OutBus]		out_9_31_i;
wire signed [`OutBus]		out_9_32_r;
wire signed [`OutBus]		out_9_32_i;
wire signed [`OutBus]		out_10_1_r;
wire signed [`OutBus]		out_10_1_i;
wire signed [`OutBus]		out_10_2_r;
wire signed [`OutBus]		out_10_2_i;
wire signed [`OutBus]		out_10_3_r;
wire signed [`OutBus]		out_10_3_i;
wire signed [`OutBus]		out_10_4_r;
wire signed [`OutBus]		out_10_4_i;
wire signed [`OutBus]		out_10_5_r;
wire signed [`OutBus]		out_10_5_i;
wire signed [`OutBus]		out_10_6_r;
wire signed [`OutBus]		out_10_6_i;
wire signed [`OutBus]		out_10_7_r;
wire signed [`OutBus]		out_10_7_i;
wire signed [`OutBus]		out_10_8_r;
wire signed [`OutBus]		out_10_8_i;
wire signed [`OutBus]		out_10_9_r;
wire signed [`OutBus]		out_10_9_i;
wire signed [`OutBus]		out_10_10_r;
wire signed [`OutBus]		out_10_10_i;
wire signed [`OutBus]		out_10_11_r;
wire signed [`OutBus]		out_10_11_i;
wire signed [`OutBus]		out_10_12_r;
wire signed [`OutBus]		out_10_12_i;
wire signed [`OutBus]		out_10_13_r;
wire signed [`OutBus]		out_10_13_i;
wire signed [`OutBus]		out_10_14_r;
wire signed [`OutBus]		out_10_14_i;
wire signed [`OutBus]		out_10_15_r;
wire signed [`OutBus]		out_10_15_i;
wire signed [`OutBus]		out_10_16_r;
wire signed [`OutBus]		out_10_16_i;
wire signed [`OutBus]		out_10_17_r;
wire signed [`OutBus]		out_10_17_i;
wire signed [`OutBus]		out_10_18_r;
wire signed [`OutBus]		out_10_18_i;
wire signed [`OutBus]		out_10_19_r;
wire signed [`OutBus]		out_10_19_i;
wire signed [`OutBus]		out_10_20_r;
wire signed [`OutBus]		out_10_20_i;
wire signed [`OutBus]		out_10_21_r;
wire signed [`OutBus]		out_10_21_i;
wire signed [`OutBus]		out_10_22_r;
wire signed [`OutBus]		out_10_22_i;
wire signed [`OutBus]		out_10_23_r;
wire signed [`OutBus]		out_10_23_i;
wire signed [`OutBus]		out_10_24_r;
wire signed [`OutBus]		out_10_24_i;
wire signed [`OutBus]		out_10_25_r;
wire signed [`OutBus]		out_10_25_i;
wire signed [`OutBus]		out_10_26_r;
wire signed [`OutBus]		out_10_26_i;
wire signed [`OutBus]		out_10_27_r;
wire signed [`OutBus]		out_10_27_i;
wire signed [`OutBus]		out_10_28_r;
wire signed [`OutBus]		out_10_28_i;
wire signed [`OutBus]		out_10_29_r;
wire signed [`OutBus]		out_10_29_i;
wire signed [`OutBus]		out_10_30_r;
wire signed [`OutBus]		out_10_30_i;
wire signed [`OutBus]		out_10_31_r;
wire signed [`OutBus]		out_10_31_i;
wire signed [`OutBus]		out_10_32_r;
wire signed [`OutBus]		out_10_32_i;
wire signed [`OutBus]		out_11_1_r;
wire signed [`OutBus]		out_11_1_i;
wire signed [`OutBus]		out_11_2_r;
wire signed [`OutBus]		out_11_2_i;
wire signed [`OutBus]		out_11_3_r;
wire signed [`OutBus]		out_11_3_i;
wire signed [`OutBus]		out_11_4_r;
wire signed [`OutBus]		out_11_4_i;
wire signed [`OutBus]		out_11_5_r;
wire signed [`OutBus]		out_11_5_i;
wire signed [`OutBus]		out_11_6_r;
wire signed [`OutBus]		out_11_6_i;
wire signed [`OutBus]		out_11_7_r;
wire signed [`OutBus]		out_11_7_i;
wire signed [`OutBus]		out_11_8_r;
wire signed [`OutBus]		out_11_8_i;
wire signed [`OutBus]		out_11_9_r;
wire signed [`OutBus]		out_11_9_i;
wire signed [`OutBus]		out_11_10_r;
wire signed [`OutBus]		out_11_10_i;
wire signed [`OutBus]		out_11_11_r;
wire signed [`OutBus]		out_11_11_i;
wire signed [`OutBus]		out_11_12_r;
wire signed [`OutBus]		out_11_12_i;
wire signed [`OutBus]		out_11_13_r;
wire signed [`OutBus]		out_11_13_i;
wire signed [`OutBus]		out_11_14_r;
wire signed [`OutBus]		out_11_14_i;
wire signed [`OutBus]		out_11_15_r;
wire signed [`OutBus]		out_11_15_i;
wire signed [`OutBus]		out_11_16_r;
wire signed [`OutBus]		out_11_16_i;
wire signed [`OutBus]		out_11_17_r;
wire signed [`OutBus]		out_11_17_i;
wire signed [`OutBus]		out_11_18_r;
wire signed [`OutBus]		out_11_18_i;
wire signed [`OutBus]		out_11_19_r;
wire signed [`OutBus]		out_11_19_i;
wire signed [`OutBus]		out_11_20_r;
wire signed [`OutBus]		out_11_20_i;
wire signed [`OutBus]		out_11_21_r;
wire signed [`OutBus]		out_11_21_i;
wire signed [`OutBus]		out_11_22_r;
wire signed [`OutBus]		out_11_22_i;
wire signed [`OutBus]		out_11_23_r;
wire signed [`OutBus]		out_11_23_i;
wire signed [`OutBus]		out_11_24_r;
wire signed [`OutBus]		out_11_24_i;
wire signed [`OutBus]		out_11_25_r;
wire signed [`OutBus]		out_11_25_i;
wire signed [`OutBus]		out_11_26_r;
wire signed [`OutBus]		out_11_26_i;
wire signed [`OutBus]		out_11_27_r;
wire signed [`OutBus]		out_11_27_i;
wire signed [`OutBus]		out_11_28_r;
wire signed [`OutBus]		out_11_28_i;
wire signed [`OutBus]		out_11_29_r;
wire signed [`OutBus]		out_11_29_i;
wire signed [`OutBus]		out_11_30_r;
wire signed [`OutBus]		out_11_30_i;
wire signed [`OutBus]		out_11_31_r;
wire signed [`OutBus]		out_11_31_i;
wire signed [`OutBus]		out_11_32_r;
wire signed [`OutBus]		out_11_32_i;
wire signed [`OutBus]		out_12_1_r;
wire signed [`OutBus]		out_12_1_i;
wire signed [`OutBus]		out_12_2_r;
wire signed [`OutBus]		out_12_2_i;
wire signed [`OutBus]		out_12_3_r;
wire signed [`OutBus]		out_12_3_i;
wire signed [`OutBus]		out_12_4_r;
wire signed [`OutBus]		out_12_4_i;
wire signed [`OutBus]		out_12_5_r;
wire signed [`OutBus]		out_12_5_i;
wire signed [`OutBus]		out_12_6_r;
wire signed [`OutBus]		out_12_6_i;
wire signed [`OutBus]		out_12_7_r;
wire signed [`OutBus]		out_12_7_i;
wire signed [`OutBus]		out_12_8_r;
wire signed [`OutBus]		out_12_8_i;
wire signed [`OutBus]		out_12_9_r;
wire signed [`OutBus]		out_12_9_i;
wire signed [`OutBus]		out_12_10_r;
wire signed [`OutBus]		out_12_10_i;
wire signed [`OutBus]		out_12_11_r;
wire signed [`OutBus]		out_12_11_i;
wire signed [`OutBus]		out_12_12_r;
wire signed [`OutBus]		out_12_12_i;
wire signed [`OutBus]		out_12_13_r;
wire signed [`OutBus]		out_12_13_i;
wire signed [`OutBus]		out_12_14_r;
wire signed [`OutBus]		out_12_14_i;
wire signed [`OutBus]		out_12_15_r;
wire signed [`OutBus]		out_12_15_i;
wire signed [`OutBus]		out_12_16_r;
wire signed [`OutBus]		out_12_16_i;
wire signed [`OutBus]		out_12_17_r;
wire signed [`OutBus]		out_12_17_i;
wire signed [`OutBus]		out_12_18_r;
wire signed [`OutBus]		out_12_18_i;
wire signed [`OutBus]		out_12_19_r;
wire signed [`OutBus]		out_12_19_i;
wire signed [`OutBus]		out_12_20_r;
wire signed [`OutBus]		out_12_20_i;
wire signed [`OutBus]		out_12_21_r;
wire signed [`OutBus]		out_12_21_i;
wire signed [`OutBus]		out_12_22_r;
wire signed [`OutBus]		out_12_22_i;
wire signed [`OutBus]		out_12_23_r;
wire signed [`OutBus]		out_12_23_i;
wire signed [`OutBus]		out_12_24_r;
wire signed [`OutBus]		out_12_24_i;
wire signed [`OutBus]		out_12_25_r;
wire signed [`OutBus]		out_12_25_i;
wire signed [`OutBus]		out_12_26_r;
wire signed [`OutBus]		out_12_26_i;
wire signed [`OutBus]		out_12_27_r;
wire signed [`OutBus]		out_12_27_i;
wire signed [`OutBus]		out_12_28_r;
wire signed [`OutBus]		out_12_28_i;
wire signed [`OutBus]		out_12_29_r;
wire signed [`OutBus]		out_12_29_i;
wire signed [`OutBus]		out_12_30_r;
wire signed [`OutBus]		out_12_30_i;
wire signed [`OutBus]		out_12_31_r;
wire signed [`OutBus]		out_12_31_i;
wire signed [`OutBus]		out_12_32_r;
wire signed [`OutBus]		out_12_32_i;
wire signed [`OutBus]		out_13_1_r;
wire signed [`OutBus]		out_13_1_i;
wire signed [`OutBus]		out_13_2_r;
wire signed [`OutBus]		out_13_2_i;
wire signed [`OutBus]		out_13_3_r;
wire signed [`OutBus]		out_13_3_i;
wire signed [`OutBus]		out_13_4_r;
wire signed [`OutBus]		out_13_4_i;
wire signed [`OutBus]		out_13_5_r;
wire signed [`OutBus]		out_13_5_i;
wire signed [`OutBus]		out_13_6_r;
wire signed [`OutBus]		out_13_6_i;
wire signed [`OutBus]		out_13_7_r;
wire signed [`OutBus]		out_13_7_i;
wire signed [`OutBus]		out_13_8_r;
wire signed [`OutBus]		out_13_8_i;
wire signed [`OutBus]		out_13_9_r;
wire signed [`OutBus]		out_13_9_i;
wire signed [`OutBus]		out_13_10_r;
wire signed [`OutBus]		out_13_10_i;
wire signed [`OutBus]		out_13_11_r;
wire signed [`OutBus]		out_13_11_i;
wire signed [`OutBus]		out_13_12_r;
wire signed [`OutBus]		out_13_12_i;
wire signed [`OutBus]		out_13_13_r;
wire signed [`OutBus]		out_13_13_i;
wire signed [`OutBus]		out_13_14_r;
wire signed [`OutBus]		out_13_14_i;
wire signed [`OutBus]		out_13_15_r;
wire signed [`OutBus]		out_13_15_i;
wire signed [`OutBus]		out_13_16_r;
wire signed [`OutBus]		out_13_16_i;
wire signed [`OutBus]		out_13_17_r;
wire signed [`OutBus]		out_13_17_i;
wire signed [`OutBus]		out_13_18_r;
wire signed [`OutBus]		out_13_18_i;
wire signed [`OutBus]		out_13_19_r;
wire signed [`OutBus]		out_13_19_i;
wire signed [`OutBus]		out_13_20_r;
wire signed [`OutBus]		out_13_20_i;
wire signed [`OutBus]		out_13_21_r;
wire signed [`OutBus]		out_13_21_i;
wire signed [`OutBus]		out_13_22_r;
wire signed [`OutBus]		out_13_22_i;
wire signed [`OutBus]		out_13_23_r;
wire signed [`OutBus]		out_13_23_i;
wire signed [`OutBus]		out_13_24_r;
wire signed [`OutBus]		out_13_24_i;
wire signed [`OutBus]		out_13_25_r;
wire signed [`OutBus]		out_13_25_i;
wire signed [`OutBus]		out_13_26_r;
wire signed [`OutBus]		out_13_26_i;
wire signed [`OutBus]		out_13_27_r;
wire signed [`OutBus]		out_13_27_i;
wire signed [`OutBus]		out_13_28_r;
wire signed [`OutBus]		out_13_28_i;
wire signed [`OutBus]		out_13_29_r;
wire signed [`OutBus]		out_13_29_i;
wire signed [`OutBus]		out_13_30_r;
wire signed [`OutBus]		out_13_30_i;
wire signed [`OutBus]		out_13_31_r;
wire signed [`OutBus]		out_13_31_i;
wire signed [`OutBus]		out_13_32_r;
wire signed [`OutBus]		out_13_32_i;
wire signed [`OutBus]		out_14_1_r;
wire signed [`OutBus]		out_14_1_i;
wire signed [`OutBus]		out_14_2_r;
wire signed [`OutBus]		out_14_2_i;
wire signed [`OutBus]		out_14_3_r;
wire signed [`OutBus]		out_14_3_i;
wire signed [`OutBus]		out_14_4_r;
wire signed [`OutBus]		out_14_4_i;
wire signed [`OutBus]		out_14_5_r;
wire signed [`OutBus]		out_14_5_i;
wire signed [`OutBus]		out_14_6_r;
wire signed [`OutBus]		out_14_6_i;
wire signed [`OutBus]		out_14_7_r;
wire signed [`OutBus]		out_14_7_i;
wire signed [`OutBus]		out_14_8_r;
wire signed [`OutBus]		out_14_8_i;
wire signed [`OutBus]		out_14_9_r;
wire signed [`OutBus]		out_14_9_i;
wire signed [`OutBus]		out_14_10_r;
wire signed [`OutBus]		out_14_10_i;
wire signed [`OutBus]		out_14_11_r;
wire signed [`OutBus]		out_14_11_i;
wire signed [`OutBus]		out_14_12_r;
wire signed [`OutBus]		out_14_12_i;
wire signed [`OutBus]		out_14_13_r;
wire signed [`OutBus]		out_14_13_i;
wire signed [`OutBus]		out_14_14_r;
wire signed [`OutBus]		out_14_14_i;
wire signed [`OutBus]		out_14_15_r;
wire signed [`OutBus]		out_14_15_i;
wire signed [`OutBus]		out_14_16_r;
wire signed [`OutBus]		out_14_16_i;
wire signed [`OutBus]		out_14_17_r;
wire signed [`OutBus]		out_14_17_i;
wire signed [`OutBus]		out_14_18_r;
wire signed [`OutBus]		out_14_18_i;
wire signed [`OutBus]		out_14_19_r;
wire signed [`OutBus]		out_14_19_i;
wire signed [`OutBus]		out_14_20_r;
wire signed [`OutBus]		out_14_20_i;
wire signed [`OutBus]		out_14_21_r;
wire signed [`OutBus]		out_14_21_i;
wire signed [`OutBus]		out_14_22_r;
wire signed [`OutBus]		out_14_22_i;
wire signed [`OutBus]		out_14_23_r;
wire signed [`OutBus]		out_14_23_i;
wire signed [`OutBus]		out_14_24_r;
wire signed [`OutBus]		out_14_24_i;
wire signed [`OutBus]		out_14_25_r;
wire signed [`OutBus]		out_14_25_i;
wire signed [`OutBus]		out_14_26_r;
wire signed [`OutBus]		out_14_26_i;
wire signed [`OutBus]		out_14_27_r;
wire signed [`OutBus]		out_14_27_i;
wire signed [`OutBus]		out_14_28_r;
wire signed [`OutBus]		out_14_28_i;
wire signed [`OutBus]		out_14_29_r;
wire signed [`OutBus]		out_14_29_i;
wire signed [`OutBus]		out_14_30_r;
wire signed [`OutBus]		out_14_30_i;
wire signed [`OutBus]		out_14_31_r;
wire signed [`OutBus]		out_14_31_i;
wire signed [`OutBus]		out_14_32_r;
wire signed [`OutBus]		out_14_32_i;
wire signed [`OutBus]		out_15_1_r;
wire signed [`OutBus]		out_15_1_i;
wire signed [`OutBus]		out_15_2_r;
wire signed [`OutBus]		out_15_2_i;
wire signed [`OutBus]		out_15_3_r;
wire signed [`OutBus]		out_15_3_i;
wire signed [`OutBus]		out_15_4_r;
wire signed [`OutBus]		out_15_4_i;
wire signed [`OutBus]		out_15_5_r;
wire signed [`OutBus]		out_15_5_i;
wire signed [`OutBus]		out_15_6_r;
wire signed [`OutBus]		out_15_6_i;
wire signed [`OutBus]		out_15_7_r;
wire signed [`OutBus]		out_15_7_i;
wire signed [`OutBus]		out_15_8_r;
wire signed [`OutBus]		out_15_8_i;
wire signed [`OutBus]		out_15_9_r;
wire signed [`OutBus]		out_15_9_i;
wire signed [`OutBus]		out_15_10_r;
wire signed [`OutBus]		out_15_10_i;
wire signed [`OutBus]		out_15_11_r;
wire signed [`OutBus]		out_15_11_i;
wire signed [`OutBus]		out_15_12_r;
wire signed [`OutBus]		out_15_12_i;
wire signed [`OutBus]		out_15_13_r;
wire signed [`OutBus]		out_15_13_i;
wire signed [`OutBus]		out_15_14_r;
wire signed [`OutBus]		out_15_14_i;
wire signed [`OutBus]		out_15_15_r;
wire signed [`OutBus]		out_15_15_i;
wire signed [`OutBus]		out_15_16_r;
wire signed [`OutBus]		out_15_16_i;
wire signed [`OutBus]		out_15_17_r;
wire signed [`OutBus]		out_15_17_i;
wire signed [`OutBus]		out_15_18_r;
wire signed [`OutBus]		out_15_18_i;
wire signed [`OutBus]		out_15_19_r;
wire signed [`OutBus]		out_15_19_i;
wire signed [`OutBus]		out_15_20_r;
wire signed [`OutBus]		out_15_20_i;
wire signed [`OutBus]		out_15_21_r;
wire signed [`OutBus]		out_15_21_i;
wire signed [`OutBus]		out_15_22_r;
wire signed [`OutBus]		out_15_22_i;
wire signed [`OutBus]		out_15_23_r;
wire signed [`OutBus]		out_15_23_i;
wire signed [`OutBus]		out_15_24_r;
wire signed [`OutBus]		out_15_24_i;
wire signed [`OutBus]		out_15_25_r;
wire signed [`OutBus]		out_15_25_i;
wire signed [`OutBus]		out_15_26_r;
wire signed [`OutBus]		out_15_26_i;
wire signed [`OutBus]		out_15_27_r;
wire signed [`OutBus]		out_15_27_i;
wire signed [`OutBus]		out_15_28_r;
wire signed [`OutBus]		out_15_28_i;
wire signed [`OutBus]		out_15_29_r;
wire signed [`OutBus]		out_15_29_i;
wire signed [`OutBus]		out_15_30_r;
wire signed [`OutBus]		out_15_30_i;
wire signed [`OutBus]		out_15_31_r;
wire signed [`OutBus]		out_15_31_i;
wire signed [`OutBus]		out_15_32_r;
wire signed [`OutBus]		out_15_32_i;
wire signed [`OutBus]		out_16_1_r;
wire signed [`OutBus]		out_16_1_i;
wire signed [`OutBus]		out_16_2_r;
wire signed [`OutBus]		out_16_2_i;
wire signed [`OutBus]		out_16_3_r;
wire signed [`OutBus]		out_16_3_i;
wire signed [`OutBus]		out_16_4_r;
wire signed [`OutBus]		out_16_4_i;
wire signed [`OutBus]		out_16_5_r;
wire signed [`OutBus]		out_16_5_i;
wire signed [`OutBus]		out_16_6_r;
wire signed [`OutBus]		out_16_6_i;
wire signed [`OutBus]		out_16_7_r;
wire signed [`OutBus]		out_16_7_i;
wire signed [`OutBus]		out_16_8_r;
wire signed [`OutBus]		out_16_8_i;
wire signed [`OutBus]		out_16_9_r;
wire signed [`OutBus]		out_16_9_i;
wire signed [`OutBus]		out_16_10_r;
wire signed [`OutBus]		out_16_10_i;
wire signed [`OutBus]		out_16_11_r;
wire signed [`OutBus]		out_16_11_i;
wire signed [`OutBus]		out_16_12_r;
wire signed [`OutBus]		out_16_12_i;
wire signed [`OutBus]		out_16_13_r;
wire signed [`OutBus]		out_16_13_i;
wire signed [`OutBus]		out_16_14_r;
wire signed [`OutBus]		out_16_14_i;
wire signed [`OutBus]		out_16_15_r;
wire signed [`OutBus]		out_16_15_i;
wire signed [`OutBus]		out_16_16_r;
wire signed [`OutBus]		out_16_16_i;
wire signed [`OutBus]		out_16_17_r;
wire signed [`OutBus]		out_16_17_i;
wire signed [`OutBus]		out_16_18_r;
wire signed [`OutBus]		out_16_18_i;
wire signed [`OutBus]		out_16_19_r;
wire signed [`OutBus]		out_16_19_i;
wire signed [`OutBus]		out_16_20_r;
wire signed [`OutBus]		out_16_20_i;
wire signed [`OutBus]		out_16_21_r;
wire signed [`OutBus]		out_16_21_i;
wire signed [`OutBus]		out_16_22_r;
wire signed [`OutBus]		out_16_22_i;
wire signed [`OutBus]		out_16_23_r;
wire signed [`OutBus]		out_16_23_i;
wire signed [`OutBus]		out_16_24_r;
wire signed [`OutBus]		out_16_24_i;
wire signed [`OutBus]		out_16_25_r;
wire signed [`OutBus]		out_16_25_i;
wire signed [`OutBus]		out_16_26_r;
wire signed [`OutBus]		out_16_26_i;
wire signed [`OutBus]		out_16_27_r;
wire signed [`OutBus]		out_16_27_i;
wire signed [`OutBus]		out_16_28_r;
wire signed [`OutBus]		out_16_28_i;
wire signed [`OutBus]		out_16_29_r;
wire signed [`OutBus]		out_16_29_i;
wire signed [`OutBus]		out_16_30_r;
wire signed [`OutBus]		out_16_30_i;
wire signed [`OutBus]		out_16_31_r;
wire signed [`OutBus]		out_16_31_i;
wire signed [`OutBus]		out_16_32_r;
wire signed [`OutBus]		out_16_32_i;
wire signed [`OutBus]		out_17_1_r;
wire signed [`OutBus]		out_17_1_i;
wire signed [`OutBus]		out_17_2_r;
wire signed [`OutBus]		out_17_2_i;
wire signed [`OutBus]		out_17_3_r;
wire signed [`OutBus]		out_17_3_i;
wire signed [`OutBus]		out_17_4_r;
wire signed [`OutBus]		out_17_4_i;
wire signed [`OutBus]		out_17_5_r;
wire signed [`OutBus]		out_17_5_i;
wire signed [`OutBus]		out_17_6_r;
wire signed [`OutBus]		out_17_6_i;
wire signed [`OutBus]		out_17_7_r;
wire signed [`OutBus]		out_17_7_i;
wire signed [`OutBus]		out_17_8_r;
wire signed [`OutBus]		out_17_8_i;
wire signed [`OutBus]		out_17_9_r;
wire signed [`OutBus]		out_17_9_i;
wire signed [`OutBus]		out_17_10_r;
wire signed [`OutBus]		out_17_10_i;
wire signed [`OutBus]		out_17_11_r;
wire signed [`OutBus]		out_17_11_i;
wire signed [`OutBus]		out_17_12_r;
wire signed [`OutBus]		out_17_12_i;
wire signed [`OutBus]		out_17_13_r;
wire signed [`OutBus]		out_17_13_i;
wire signed [`OutBus]		out_17_14_r;
wire signed [`OutBus]		out_17_14_i;
wire signed [`OutBus]		out_17_15_r;
wire signed [`OutBus]		out_17_15_i;
wire signed [`OutBus]		out_17_16_r;
wire signed [`OutBus]		out_17_16_i;
wire signed [`OutBus]		out_17_17_r;
wire signed [`OutBus]		out_17_17_i;
wire signed [`OutBus]		out_17_18_r;
wire signed [`OutBus]		out_17_18_i;
wire signed [`OutBus]		out_17_19_r;
wire signed [`OutBus]		out_17_19_i;
wire signed [`OutBus]		out_17_20_r;
wire signed [`OutBus]		out_17_20_i;
wire signed [`OutBus]		out_17_21_r;
wire signed [`OutBus]		out_17_21_i;
wire signed [`OutBus]		out_17_22_r;
wire signed [`OutBus]		out_17_22_i;
wire signed [`OutBus]		out_17_23_r;
wire signed [`OutBus]		out_17_23_i;
wire signed [`OutBus]		out_17_24_r;
wire signed [`OutBus]		out_17_24_i;
wire signed [`OutBus]		out_17_25_r;
wire signed [`OutBus]		out_17_25_i;
wire signed [`OutBus]		out_17_26_r;
wire signed [`OutBus]		out_17_26_i;
wire signed [`OutBus]		out_17_27_r;
wire signed [`OutBus]		out_17_27_i;
wire signed [`OutBus]		out_17_28_r;
wire signed [`OutBus]		out_17_28_i;
wire signed [`OutBus]		out_17_29_r;
wire signed [`OutBus]		out_17_29_i;
wire signed [`OutBus]		out_17_30_r;
wire signed [`OutBus]		out_17_30_i;
wire signed [`OutBus]		out_17_31_r;
wire signed [`OutBus]		out_17_31_i;
wire signed [`OutBus]		out_17_32_r;
wire signed [`OutBus]		out_17_32_i;
wire signed [`OutBus]		out_18_1_r;
wire signed [`OutBus]		out_18_1_i;
wire signed [`OutBus]		out_18_2_r;
wire signed [`OutBus]		out_18_2_i;
wire signed [`OutBus]		out_18_3_r;
wire signed [`OutBus]		out_18_3_i;
wire signed [`OutBus]		out_18_4_r;
wire signed [`OutBus]		out_18_4_i;
wire signed [`OutBus]		out_18_5_r;
wire signed [`OutBus]		out_18_5_i;
wire signed [`OutBus]		out_18_6_r;
wire signed [`OutBus]		out_18_6_i;
wire signed [`OutBus]		out_18_7_r;
wire signed [`OutBus]		out_18_7_i;
wire signed [`OutBus]		out_18_8_r;
wire signed [`OutBus]		out_18_8_i;
wire signed [`OutBus]		out_18_9_r;
wire signed [`OutBus]		out_18_9_i;
wire signed [`OutBus]		out_18_10_r;
wire signed [`OutBus]		out_18_10_i;
wire signed [`OutBus]		out_18_11_r;
wire signed [`OutBus]		out_18_11_i;
wire signed [`OutBus]		out_18_12_r;
wire signed [`OutBus]		out_18_12_i;
wire signed [`OutBus]		out_18_13_r;
wire signed [`OutBus]		out_18_13_i;
wire signed [`OutBus]		out_18_14_r;
wire signed [`OutBus]		out_18_14_i;
wire signed [`OutBus]		out_18_15_r;
wire signed [`OutBus]		out_18_15_i;
wire signed [`OutBus]		out_18_16_r;
wire signed [`OutBus]		out_18_16_i;
wire signed [`OutBus]		out_18_17_r;
wire signed [`OutBus]		out_18_17_i;
wire signed [`OutBus]		out_18_18_r;
wire signed [`OutBus]		out_18_18_i;
wire signed [`OutBus]		out_18_19_r;
wire signed [`OutBus]		out_18_19_i;
wire signed [`OutBus]		out_18_20_r;
wire signed [`OutBus]		out_18_20_i;
wire signed [`OutBus]		out_18_21_r;
wire signed [`OutBus]		out_18_21_i;
wire signed [`OutBus]		out_18_22_r;
wire signed [`OutBus]		out_18_22_i;
wire signed [`OutBus]		out_18_23_r;
wire signed [`OutBus]		out_18_23_i;
wire signed [`OutBus]		out_18_24_r;
wire signed [`OutBus]		out_18_24_i;
wire signed [`OutBus]		out_18_25_r;
wire signed [`OutBus]		out_18_25_i;
wire signed [`OutBus]		out_18_26_r;
wire signed [`OutBus]		out_18_26_i;
wire signed [`OutBus]		out_18_27_r;
wire signed [`OutBus]		out_18_27_i;
wire signed [`OutBus]		out_18_28_r;
wire signed [`OutBus]		out_18_28_i;
wire signed [`OutBus]		out_18_29_r;
wire signed [`OutBus]		out_18_29_i;
wire signed [`OutBus]		out_18_30_r;
wire signed [`OutBus]		out_18_30_i;
wire signed [`OutBus]		out_18_31_r;
wire signed [`OutBus]		out_18_31_i;
wire signed [`OutBus]		out_18_32_r;
wire signed [`OutBus]		out_18_32_i;
wire signed [`OutBus]		out_19_1_r;
wire signed [`OutBus]		out_19_1_i;
wire signed [`OutBus]		out_19_2_r;
wire signed [`OutBus]		out_19_2_i;
wire signed [`OutBus]		out_19_3_r;
wire signed [`OutBus]		out_19_3_i;
wire signed [`OutBus]		out_19_4_r;
wire signed [`OutBus]		out_19_4_i;
wire signed [`OutBus]		out_19_5_r;
wire signed [`OutBus]		out_19_5_i;
wire signed [`OutBus]		out_19_6_r;
wire signed [`OutBus]		out_19_6_i;
wire signed [`OutBus]		out_19_7_r;
wire signed [`OutBus]		out_19_7_i;
wire signed [`OutBus]		out_19_8_r;
wire signed [`OutBus]		out_19_8_i;
wire signed [`OutBus]		out_19_9_r;
wire signed [`OutBus]		out_19_9_i;
wire signed [`OutBus]		out_19_10_r;
wire signed [`OutBus]		out_19_10_i;
wire signed [`OutBus]		out_19_11_r;
wire signed [`OutBus]		out_19_11_i;
wire signed [`OutBus]		out_19_12_r;
wire signed [`OutBus]		out_19_12_i;
wire signed [`OutBus]		out_19_13_r;
wire signed [`OutBus]		out_19_13_i;
wire signed [`OutBus]		out_19_14_r;
wire signed [`OutBus]		out_19_14_i;
wire signed [`OutBus]		out_19_15_r;
wire signed [`OutBus]		out_19_15_i;
wire signed [`OutBus]		out_19_16_r;
wire signed [`OutBus]		out_19_16_i;
wire signed [`OutBus]		out_19_17_r;
wire signed [`OutBus]		out_19_17_i;
wire signed [`OutBus]		out_19_18_r;
wire signed [`OutBus]		out_19_18_i;
wire signed [`OutBus]		out_19_19_r;
wire signed [`OutBus]		out_19_19_i;
wire signed [`OutBus]		out_19_20_r;
wire signed [`OutBus]		out_19_20_i;
wire signed [`OutBus]		out_19_21_r;
wire signed [`OutBus]		out_19_21_i;
wire signed [`OutBus]		out_19_22_r;
wire signed [`OutBus]		out_19_22_i;
wire signed [`OutBus]		out_19_23_r;
wire signed [`OutBus]		out_19_23_i;
wire signed [`OutBus]		out_19_24_r;
wire signed [`OutBus]		out_19_24_i;
wire signed [`OutBus]		out_19_25_r;
wire signed [`OutBus]		out_19_25_i;
wire signed [`OutBus]		out_19_26_r;
wire signed [`OutBus]		out_19_26_i;
wire signed [`OutBus]		out_19_27_r;
wire signed [`OutBus]		out_19_27_i;
wire signed [`OutBus]		out_19_28_r;
wire signed [`OutBus]		out_19_28_i;
wire signed [`OutBus]		out_19_29_r;
wire signed [`OutBus]		out_19_29_i;
wire signed [`OutBus]		out_19_30_r;
wire signed [`OutBus]		out_19_30_i;
wire signed [`OutBus]		out_19_31_r;
wire signed [`OutBus]		out_19_31_i;
wire signed [`OutBus]		out_19_32_r;
wire signed [`OutBus]		out_19_32_i;
wire signed [`OutBus]		out_20_1_r;
wire signed [`OutBus]		out_20_1_i;
wire signed [`OutBus]		out_20_2_r;
wire signed [`OutBus]		out_20_2_i;
wire signed [`OutBus]		out_20_3_r;
wire signed [`OutBus]		out_20_3_i;
wire signed [`OutBus]		out_20_4_r;
wire signed [`OutBus]		out_20_4_i;
wire signed [`OutBus]		out_20_5_r;
wire signed [`OutBus]		out_20_5_i;
wire signed [`OutBus]		out_20_6_r;
wire signed [`OutBus]		out_20_6_i;
wire signed [`OutBus]		out_20_7_r;
wire signed [`OutBus]		out_20_7_i;
wire signed [`OutBus]		out_20_8_r;
wire signed [`OutBus]		out_20_8_i;
wire signed [`OutBus]		out_20_9_r;
wire signed [`OutBus]		out_20_9_i;
wire signed [`OutBus]		out_20_10_r;
wire signed [`OutBus]		out_20_10_i;
wire signed [`OutBus]		out_20_11_r;
wire signed [`OutBus]		out_20_11_i;
wire signed [`OutBus]		out_20_12_r;
wire signed [`OutBus]		out_20_12_i;
wire signed [`OutBus]		out_20_13_r;
wire signed [`OutBus]		out_20_13_i;
wire signed [`OutBus]		out_20_14_r;
wire signed [`OutBus]		out_20_14_i;
wire signed [`OutBus]		out_20_15_r;
wire signed [`OutBus]		out_20_15_i;
wire signed [`OutBus]		out_20_16_r;
wire signed [`OutBus]		out_20_16_i;
wire signed [`OutBus]		out_20_17_r;
wire signed [`OutBus]		out_20_17_i;
wire signed [`OutBus]		out_20_18_r;
wire signed [`OutBus]		out_20_18_i;
wire signed [`OutBus]		out_20_19_r;
wire signed [`OutBus]		out_20_19_i;
wire signed [`OutBus]		out_20_20_r;
wire signed [`OutBus]		out_20_20_i;
wire signed [`OutBus]		out_20_21_r;
wire signed [`OutBus]		out_20_21_i;
wire signed [`OutBus]		out_20_22_r;
wire signed [`OutBus]		out_20_22_i;
wire signed [`OutBus]		out_20_23_r;
wire signed [`OutBus]		out_20_23_i;
wire signed [`OutBus]		out_20_24_r;
wire signed [`OutBus]		out_20_24_i;
wire signed [`OutBus]		out_20_25_r;
wire signed [`OutBus]		out_20_25_i;
wire signed [`OutBus]		out_20_26_r;
wire signed [`OutBus]		out_20_26_i;
wire signed [`OutBus]		out_20_27_r;
wire signed [`OutBus]		out_20_27_i;
wire signed [`OutBus]		out_20_28_r;
wire signed [`OutBus]		out_20_28_i;
wire signed [`OutBus]		out_20_29_r;
wire signed [`OutBus]		out_20_29_i;
wire signed [`OutBus]		out_20_30_r;
wire signed [`OutBus]		out_20_30_i;
wire signed [`OutBus]		out_20_31_r;
wire signed [`OutBus]		out_20_31_i;
wire signed [`OutBus]		out_20_32_r;
wire signed [`OutBus]		out_20_32_i;
wire signed [`OutBus]		out_21_1_r;
wire signed [`OutBus]		out_21_1_i;
wire signed [`OutBus]		out_21_2_r;
wire signed [`OutBus]		out_21_2_i;
wire signed [`OutBus]		out_21_3_r;
wire signed [`OutBus]		out_21_3_i;
wire signed [`OutBus]		out_21_4_r;
wire signed [`OutBus]		out_21_4_i;
wire signed [`OutBus]		out_21_5_r;
wire signed [`OutBus]		out_21_5_i;
wire signed [`OutBus]		out_21_6_r;
wire signed [`OutBus]		out_21_6_i;
wire signed [`OutBus]		out_21_7_r;
wire signed [`OutBus]		out_21_7_i;
wire signed [`OutBus]		out_21_8_r;
wire signed [`OutBus]		out_21_8_i;
wire signed [`OutBus]		out_21_9_r;
wire signed [`OutBus]		out_21_9_i;
wire signed [`OutBus]		out_21_10_r;
wire signed [`OutBus]		out_21_10_i;
wire signed [`OutBus]		out_21_11_r;
wire signed [`OutBus]		out_21_11_i;
wire signed [`OutBus]		out_21_12_r;
wire signed [`OutBus]		out_21_12_i;
wire signed [`OutBus]		out_21_13_r;
wire signed [`OutBus]		out_21_13_i;
wire signed [`OutBus]		out_21_14_r;
wire signed [`OutBus]		out_21_14_i;
wire signed [`OutBus]		out_21_15_r;
wire signed [`OutBus]		out_21_15_i;
wire signed [`OutBus]		out_21_16_r;
wire signed [`OutBus]		out_21_16_i;
wire signed [`OutBus]		out_21_17_r;
wire signed [`OutBus]		out_21_17_i;
wire signed [`OutBus]		out_21_18_r;
wire signed [`OutBus]		out_21_18_i;
wire signed [`OutBus]		out_21_19_r;
wire signed [`OutBus]		out_21_19_i;
wire signed [`OutBus]		out_21_20_r;
wire signed [`OutBus]		out_21_20_i;
wire signed [`OutBus]		out_21_21_r;
wire signed [`OutBus]		out_21_21_i;
wire signed [`OutBus]		out_21_22_r;
wire signed [`OutBus]		out_21_22_i;
wire signed [`OutBus]		out_21_23_r;
wire signed [`OutBus]		out_21_23_i;
wire signed [`OutBus]		out_21_24_r;
wire signed [`OutBus]		out_21_24_i;
wire signed [`OutBus]		out_21_25_r;
wire signed [`OutBus]		out_21_25_i;
wire signed [`OutBus]		out_21_26_r;
wire signed [`OutBus]		out_21_26_i;
wire signed [`OutBus]		out_21_27_r;
wire signed [`OutBus]		out_21_27_i;
wire signed [`OutBus]		out_21_28_r;
wire signed [`OutBus]		out_21_28_i;
wire signed [`OutBus]		out_21_29_r;
wire signed [`OutBus]		out_21_29_i;
wire signed [`OutBus]		out_21_30_r;
wire signed [`OutBus]		out_21_30_i;
wire signed [`OutBus]		out_21_31_r;
wire signed [`OutBus]		out_21_31_i;
wire signed [`OutBus]		out_21_32_r;
wire signed [`OutBus]		out_21_32_i;
wire signed [`OutBus]		out_22_1_r;
wire signed [`OutBus]		out_22_1_i;
wire signed [`OutBus]		out_22_2_r;
wire signed [`OutBus]		out_22_2_i;
wire signed [`OutBus]		out_22_3_r;
wire signed [`OutBus]		out_22_3_i;
wire signed [`OutBus]		out_22_4_r;
wire signed [`OutBus]		out_22_4_i;
wire signed [`OutBus]		out_22_5_r;
wire signed [`OutBus]		out_22_5_i;
wire signed [`OutBus]		out_22_6_r;
wire signed [`OutBus]		out_22_6_i;
wire signed [`OutBus]		out_22_7_r;
wire signed [`OutBus]		out_22_7_i;
wire signed [`OutBus]		out_22_8_r;
wire signed [`OutBus]		out_22_8_i;
wire signed [`OutBus]		out_22_9_r;
wire signed [`OutBus]		out_22_9_i;
wire signed [`OutBus]		out_22_10_r;
wire signed [`OutBus]		out_22_10_i;
wire signed [`OutBus]		out_22_11_r;
wire signed [`OutBus]		out_22_11_i;
wire signed [`OutBus]		out_22_12_r;
wire signed [`OutBus]		out_22_12_i;
wire signed [`OutBus]		out_22_13_r;
wire signed [`OutBus]		out_22_13_i;
wire signed [`OutBus]		out_22_14_r;
wire signed [`OutBus]		out_22_14_i;
wire signed [`OutBus]		out_22_15_r;
wire signed [`OutBus]		out_22_15_i;
wire signed [`OutBus]		out_22_16_r;
wire signed [`OutBus]		out_22_16_i;
wire signed [`OutBus]		out_22_17_r;
wire signed [`OutBus]		out_22_17_i;
wire signed [`OutBus]		out_22_18_r;
wire signed [`OutBus]		out_22_18_i;
wire signed [`OutBus]		out_22_19_r;
wire signed [`OutBus]		out_22_19_i;
wire signed [`OutBus]		out_22_20_r;
wire signed [`OutBus]		out_22_20_i;
wire signed [`OutBus]		out_22_21_r;
wire signed [`OutBus]		out_22_21_i;
wire signed [`OutBus]		out_22_22_r;
wire signed [`OutBus]		out_22_22_i;
wire signed [`OutBus]		out_22_23_r;
wire signed [`OutBus]		out_22_23_i;
wire signed [`OutBus]		out_22_24_r;
wire signed [`OutBus]		out_22_24_i;
wire signed [`OutBus]		out_22_25_r;
wire signed [`OutBus]		out_22_25_i;
wire signed [`OutBus]		out_22_26_r;
wire signed [`OutBus]		out_22_26_i;
wire signed [`OutBus]		out_22_27_r;
wire signed [`OutBus]		out_22_27_i;
wire signed [`OutBus]		out_22_28_r;
wire signed [`OutBus]		out_22_28_i;
wire signed [`OutBus]		out_22_29_r;
wire signed [`OutBus]		out_22_29_i;
wire signed [`OutBus]		out_22_30_r;
wire signed [`OutBus]		out_22_30_i;
wire signed [`OutBus]		out_22_31_r;
wire signed [`OutBus]		out_22_31_i;
wire signed [`OutBus]		out_22_32_r;
wire signed [`OutBus]		out_22_32_i;
wire signed [`OutBus]		out_23_1_r;
wire signed [`OutBus]		out_23_1_i;
wire signed [`OutBus]		out_23_2_r;
wire signed [`OutBus]		out_23_2_i;
wire signed [`OutBus]		out_23_3_r;
wire signed [`OutBus]		out_23_3_i;
wire signed [`OutBus]		out_23_4_r;
wire signed [`OutBus]		out_23_4_i;
wire signed [`OutBus]		out_23_5_r;
wire signed [`OutBus]		out_23_5_i;
wire signed [`OutBus]		out_23_6_r;
wire signed [`OutBus]		out_23_6_i;
wire signed [`OutBus]		out_23_7_r;
wire signed [`OutBus]		out_23_7_i;
wire signed [`OutBus]		out_23_8_r;
wire signed [`OutBus]		out_23_8_i;
wire signed [`OutBus]		out_23_9_r;
wire signed [`OutBus]		out_23_9_i;
wire signed [`OutBus]		out_23_10_r;
wire signed [`OutBus]		out_23_10_i;
wire signed [`OutBus]		out_23_11_r;
wire signed [`OutBus]		out_23_11_i;
wire signed [`OutBus]		out_23_12_r;
wire signed [`OutBus]		out_23_12_i;
wire signed [`OutBus]		out_23_13_r;
wire signed [`OutBus]		out_23_13_i;
wire signed [`OutBus]		out_23_14_r;
wire signed [`OutBus]		out_23_14_i;
wire signed [`OutBus]		out_23_15_r;
wire signed [`OutBus]		out_23_15_i;
wire signed [`OutBus]		out_23_16_r;
wire signed [`OutBus]		out_23_16_i;
wire signed [`OutBus]		out_23_17_r;
wire signed [`OutBus]		out_23_17_i;
wire signed [`OutBus]		out_23_18_r;
wire signed [`OutBus]		out_23_18_i;
wire signed [`OutBus]		out_23_19_r;
wire signed [`OutBus]		out_23_19_i;
wire signed [`OutBus]		out_23_20_r;
wire signed [`OutBus]		out_23_20_i;
wire signed [`OutBus]		out_23_21_r;
wire signed [`OutBus]		out_23_21_i;
wire signed [`OutBus]		out_23_22_r;
wire signed [`OutBus]		out_23_22_i;
wire signed [`OutBus]		out_23_23_r;
wire signed [`OutBus]		out_23_23_i;
wire signed [`OutBus]		out_23_24_r;
wire signed [`OutBus]		out_23_24_i;
wire signed [`OutBus]		out_23_25_r;
wire signed [`OutBus]		out_23_25_i;
wire signed [`OutBus]		out_23_26_r;
wire signed [`OutBus]		out_23_26_i;
wire signed [`OutBus]		out_23_27_r;
wire signed [`OutBus]		out_23_27_i;
wire signed [`OutBus]		out_23_28_r;
wire signed [`OutBus]		out_23_28_i;
wire signed [`OutBus]		out_23_29_r;
wire signed [`OutBus]		out_23_29_i;
wire signed [`OutBus]		out_23_30_r;
wire signed [`OutBus]		out_23_30_i;
wire signed [`OutBus]		out_23_31_r;
wire signed [`OutBus]		out_23_31_i;
wire signed [`OutBus]		out_23_32_r;
wire signed [`OutBus]		out_23_32_i;
wire signed [`OutBus]		out_24_1_r;
wire signed [`OutBus]		out_24_1_i;
wire signed [`OutBus]		out_24_2_r;
wire signed [`OutBus]		out_24_2_i;
wire signed [`OutBus]		out_24_3_r;
wire signed [`OutBus]		out_24_3_i;
wire signed [`OutBus]		out_24_4_r;
wire signed [`OutBus]		out_24_4_i;
wire signed [`OutBus]		out_24_5_r;
wire signed [`OutBus]		out_24_5_i;
wire signed [`OutBus]		out_24_6_r;
wire signed [`OutBus]		out_24_6_i;
wire signed [`OutBus]		out_24_7_r;
wire signed [`OutBus]		out_24_7_i;
wire signed [`OutBus]		out_24_8_r;
wire signed [`OutBus]		out_24_8_i;
wire signed [`OutBus]		out_24_9_r;
wire signed [`OutBus]		out_24_9_i;
wire signed [`OutBus]		out_24_10_r;
wire signed [`OutBus]		out_24_10_i;
wire signed [`OutBus]		out_24_11_r;
wire signed [`OutBus]		out_24_11_i;
wire signed [`OutBus]		out_24_12_r;
wire signed [`OutBus]		out_24_12_i;
wire signed [`OutBus]		out_24_13_r;
wire signed [`OutBus]		out_24_13_i;
wire signed [`OutBus]		out_24_14_r;
wire signed [`OutBus]		out_24_14_i;
wire signed [`OutBus]		out_24_15_r;
wire signed [`OutBus]		out_24_15_i;
wire signed [`OutBus]		out_24_16_r;
wire signed [`OutBus]		out_24_16_i;
wire signed [`OutBus]		out_24_17_r;
wire signed [`OutBus]		out_24_17_i;
wire signed [`OutBus]		out_24_18_r;
wire signed [`OutBus]		out_24_18_i;
wire signed [`OutBus]		out_24_19_r;
wire signed [`OutBus]		out_24_19_i;
wire signed [`OutBus]		out_24_20_r;
wire signed [`OutBus]		out_24_20_i;
wire signed [`OutBus]		out_24_21_r;
wire signed [`OutBus]		out_24_21_i;
wire signed [`OutBus]		out_24_22_r;
wire signed [`OutBus]		out_24_22_i;
wire signed [`OutBus]		out_24_23_r;
wire signed [`OutBus]		out_24_23_i;
wire signed [`OutBus]		out_24_24_r;
wire signed [`OutBus]		out_24_24_i;
wire signed [`OutBus]		out_24_25_r;
wire signed [`OutBus]		out_24_25_i;
wire signed [`OutBus]		out_24_26_r;
wire signed [`OutBus]		out_24_26_i;
wire signed [`OutBus]		out_24_27_r;
wire signed [`OutBus]		out_24_27_i;
wire signed [`OutBus]		out_24_28_r;
wire signed [`OutBus]		out_24_28_i;
wire signed [`OutBus]		out_24_29_r;
wire signed [`OutBus]		out_24_29_i;
wire signed [`OutBus]		out_24_30_r;
wire signed [`OutBus]		out_24_30_i;
wire signed [`OutBus]		out_24_31_r;
wire signed [`OutBus]		out_24_31_i;
wire signed [`OutBus]		out_24_32_r;
wire signed [`OutBus]		out_24_32_i;
wire signed [`OutBus]		out_25_1_r;
wire signed [`OutBus]		out_25_1_i;
wire signed [`OutBus]		out_25_2_r;
wire signed [`OutBus]		out_25_2_i;
wire signed [`OutBus]		out_25_3_r;
wire signed [`OutBus]		out_25_3_i;
wire signed [`OutBus]		out_25_4_r;
wire signed [`OutBus]		out_25_4_i;
wire signed [`OutBus]		out_25_5_r;
wire signed [`OutBus]		out_25_5_i;
wire signed [`OutBus]		out_25_6_r;
wire signed [`OutBus]		out_25_6_i;
wire signed [`OutBus]		out_25_7_r;
wire signed [`OutBus]		out_25_7_i;
wire signed [`OutBus]		out_25_8_r;
wire signed [`OutBus]		out_25_8_i;
wire signed [`OutBus]		out_25_9_r;
wire signed [`OutBus]		out_25_9_i;
wire signed [`OutBus]		out_25_10_r;
wire signed [`OutBus]		out_25_10_i;
wire signed [`OutBus]		out_25_11_r;
wire signed [`OutBus]		out_25_11_i;
wire signed [`OutBus]		out_25_12_r;
wire signed [`OutBus]		out_25_12_i;
wire signed [`OutBus]		out_25_13_r;
wire signed [`OutBus]		out_25_13_i;
wire signed [`OutBus]		out_25_14_r;
wire signed [`OutBus]		out_25_14_i;
wire signed [`OutBus]		out_25_15_r;
wire signed [`OutBus]		out_25_15_i;
wire signed [`OutBus]		out_25_16_r;
wire signed [`OutBus]		out_25_16_i;
wire signed [`OutBus]		out_25_17_r;
wire signed [`OutBus]		out_25_17_i;
wire signed [`OutBus]		out_25_18_r;
wire signed [`OutBus]		out_25_18_i;
wire signed [`OutBus]		out_25_19_r;
wire signed [`OutBus]		out_25_19_i;
wire signed [`OutBus]		out_25_20_r;
wire signed [`OutBus]		out_25_20_i;
wire signed [`OutBus]		out_25_21_r;
wire signed [`OutBus]		out_25_21_i;
wire signed [`OutBus]		out_25_22_r;
wire signed [`OutBus]		out_25_22_i;
wire signed [`OutBus]		out_25_23_r;
wire signed [`OutBus]		out_25_23_i;
wire signed [`OutBus]		out_25_24_r;
wire signed [`OutBus]		out_25_24_i;
wire signed [`OutBus]		out_25_25_r;
wire signed [`OutBus]		out_25_25_i;
wire signed [`OutBus]		out_25_26_r;
wire signed [`OutBus]		out_25_26_i;
wire signed [`OutBus]		out_25_27_r;
wire signed [`OutBus]		out_25_27_i;
wire signed [`OutBus]		out_25_28_r;
wire signed [`OutBus]		out_25_28_i;
wire signed [`OutBus]		out_25_29_r;
wire signed [`OutBus]		out_25_29_i;
wire signed [`OutBus]		out_25_30_r;
wire signed [`OutBus]		out_25_30_i;
wire signed [`OutBus]		out_25_31_r;
wire signed [`OutBus]		out_25_31_i;
wire signed [`OutBus]		out_25_32_r;
wire signed [`OutBus]		out_25_32_i;
wire signed [`OutBus]		out_26_1_r;
wire signed [`OutBus]		out_26_1_i;
wire signed [`OutBus]		out_26_2_r;
wire signed [`OutBus]		out_26_2_i;
wire signed [`OutBus]		out_26_3_r;
wire signed [`OutBus]		out_26_3_i;
wire signed [`OutBus]		out_26_4_r;
wire signed [`OutBus]		out_26_4_i;
wire signed [`OutBus]		out_26_5_r;
wire signed [`OutBus]		out_26_5_i;
wire signed [`OutBus]		out_26_6_r;
wire signed [`OutBus]		out_26_6_i;
wire signed [`OutBus]		out_26_7_r;
wire signed [`OutBus]		out_26_7_i;
wire signed [`OutBus]		out_26_8_r;
wire signed [`OutBus]		out_26_8_i;
wire signed [`OutBus]		out_26_9_r;
wire signed [`OutBus]		out_26_9_i;
wire signed [`OutBus]		out_26_10_r;
wire signed [`OutBus]		out_26_10_i;
wire signed [`OutBus]		out_26_11_r;
wire signed [`OutBus]		out_26_11_i;
wire signed [`OutBus]		out_26_12_r;
wire signed [`OutBus]		out_26_12_i;
wire signed [`OutBus]		out_26_13_r;
wire signed [`OutBus]		out_26_13_i;
wire signed [`OutBus]		out_26_14_r;
wire signed [`OutBus]		out_26_14_i;
wire signed [`OutBus]		out_26_15_r;
wire signed [`OutBus]		out_26_15_i;
wire signed [`OutBus]		out_26_16_r;
wire signed [`OutBus]		out_26_16_i;
wire signed [`OutBus]		out_26_17_r;
wire signed [`OutBus]		out_26_17_i;
wire signed [`OutBus]		out_26_18_r;
wire signed [`OutBus]		out_26_18_i;
wire signed [`OutBus]		out_26_19_r;
wire signed [`OutBus]		out_26_19_i;
wire signed [`OutBus]		out_26_20_r;
wire signed [`OutBus]		out_26_20_i;
wire signed [`OutBus]		out_26_21_r;
wire signed [`OutBus]		out_26_21_i;
wire signed [`OutBus]		out_26_22_r;
wire signed [`OutBus]		out_26_22_i;
wire signed [`OutBus]		out_26_23_r;
wire signed [`OutBus]		out_26_23_i;
wire signed [`OutBus]		out_26_24_r;
wire signed [`OutBus]		out_26_24_i;
wire signed [`OutBus]		out_26_25_r;
wire signed [`OutBus]		out_26_25_i;
wire signed [`OutBus]		out_26_26_r;
wire signed [`OutBus]		out_26_26_i;
wire signed [`OutBus]		out_26_27_r;
wire signed [`OutBus]		out_26_27_i;
wire signed [`OutBus]		out_26_28_r;
wire signed [`OutBus]		out_26_28_i;
wire signed [`OutBus]		out_26_29_r;
wire signed [`OutBus]		out_26_29_i;
wire signed [`OutBus]		out_26_30_r;
wire signed [`OutBus]		out_26_30_i;
wire signed [`OutBus]		out_26_31_r;
wire signed [`OutBus]		out_26_31_i;
wire signed [`OutBus]		out_26_32_r;
wire signed [`OutBus]		out_26_32_i;
wire signed [`OutBus]		out_27_1_r;
wire signed [`OutBus]		out_27_1_i;
wire signed [`OutBus]		out_27_2_r;
wire signed [`OutBus]		out_27_2_i;
wire signed [`OutBus]		out_27_3_r;
wire signed [`OutBus]		out_27_3_i;
wire signed [`OutBus]		out_27_4_r;
wire signed [`OutBus]		out_27_4_i;
wire signed [`OutBus]		out_27_5_r;
wire signed [`OutBus]		out_27_5_i;
wire signed [`OutBus]		out_27_6_r;
wire signed [`OutBus]		out_27_6_i;
wire signed [`OutBus]		out_27_7_r;
wire signed [`OutBus]		out_27_7_i;
wire signed [`OutBus]		out_27_8_r;
wire signed [`OutBus]		out_27_8_i;
wire signed [`OutBus]		out_27_9_r;
wire signed [`OutBus]		out_27_9_i;
wire signed [`OutBus]		out_27_10_r;
wire signed [`OutBus]		out_27_10_i;
wire signed [`OutBus]		out_27_11_r;
wire signed [`OutBus]		out_27_11_i;
wire signed [`OutBus]		out_27_12_r;
wire signed [`OutBus]		out_27_12_i;
wire signed [`OutBus]		out_27_13_r;
wire signed [`OutBus]		out_27_13_i;
wire signed [`OutBus]		out_27_14_r;
wire signed [`OutBus]		out_27_14_i;
wire signed [`OutBus]		out_27_15_r;
wire signed [`OutBus]		out_27_15_i;
wire signed [`OutBus]		out_27_16_r;
wire signed [`OutBus]		out_27_16_i;
wire signed [`OutBus]		out_27_17_r;
wire signed [`OutBus]		out_27_17_i;
wire signed [`OutBus]		out_27_18_r;
wire signed [`OutBus]		out_27_18_i;
wire signed [`OutBus]		out_27_19_r;
wire signed [`OutBus]		out_27_19_i;
wire signed [`OutBus]		out_27_20_r;
wire signed [`OutBus]		out_27_20_i;
wire signed [`OutBus]		out_27_21_r;
wire signed [`OutBus]		out_27_21_i;
wire signed [`OutBus]		out_27_22_r;
wire signed [`OutBus]		out_27_22_i;
wire signed [`OutBus]		out_27_23_r;
wire signed [`OutBus]		out_27_23_i;
wire signed [`OutBus]		out_27_24_r;
wire signed [`OutBus]		out_27_24_i;
wire signed [`OutBus]		out_27_25_r;
wire signed [`OutBus]		out_27_25_i;
wire signed [`OutBus]		out_27_26_r;
wire signed [`OutBus]		out_27_26_i;
wire signed [`OutBus]		out_27_27_r;
wire signed [`OutBus]		out_27_27_i;
wire signed [`OutBus]		out_27_28_r;
wire signed [`OutBus]		out_27_28_i;
wire signed [`OutBus]		out_27_29_r;
wire signed [`OutBus]		out_27_29_i;
wire signed [`OutBus]		out_27_30_r;
wire signed [`OutBus]		out_27_30_i;
wire signed [`OutBus]		out_27_31_r;
wire signed [`OutBus]		out_27_31_i;
wire signed [`OutBus]		out_27_32_r;
wire signed [`OutBus]		out_27_32_i;
wire signed [`OutBus]		out_28_1_r;
wire signed [`OutBus]		out_28_1_i;
wire signed [`OutBus]		out_28_2_r;
wire signed [`OutBus]		out_28_2_i;
wire signed [`OutBus]		out_28_3_r;
wire signed [`OutBus]		out_28_3_i;
wire signed [`OutBus]		out_28_4_r;
wire signed [`OutBus]		out_28_4_i;
wire signed [`OutBus]		out_28_5_r;
wire signed [`OutBus]		out_28_5_i;
wire signed [`OutBus]		out_28_6_r;
wire signed [`OutBus]		out_28_6_i;
wire signed [`OutBus]		out_28_7_r;
wire signed [`OutBus]		out_28_7_i;
wire signed [`OutBus]		out_28_8_r;
wire signed [`OutBus]		out_28_8_i;
wire signed [`OutBus]		out_28_9_r;
wire signed [`OutBus]		out_28_9_i;
wire signed [`OutBus]		out_28_10_r;
wire signed [`OutBus]		out_28_10_i;
wire signed [`OutBus]		out_28_11_r;
wire signed [`OutBus]		out_28_11_i;
wire signed [`OutBus]		out_28_12_r;
wire signed [`OutBus]		out_28_12_i;
wire signed [`OutBus]		out_28_13_r;
wire signed [`OutBus]		out_28_13_i;
wire signed [`OutBus]		out_28_14_r;
wire signed [`OutBus]		out_28_14_i;
wire signed [`OutBus]		out_28_15_r;
wire signed [`OutBus]		out_28_15_i;
wire signed [`OutBus]		out_28_16_r;
wire signed [`OutBus]		out_28_16_i;
wire signed [`OutBus]		out_28_17_r;
wire signed [`OutBus]		out_28_17_i;
wire signed [`OutBus]		out_28_18_r;
wire signed [`OutBus]		out_28_18_i;
wire signed [`OutBus]		out_28_19_r;
wire signed [`OutBus]		out_28_19_i;
wire signed [`OutBus]		out_28_20_r;
wire signed [`OutBus]		out_28_20_i;
wire signed [`OutBus]		out_28_21_r;
wire signed [`OutBus]		out_28_21_i;
wire signed [`OutBus]		out_28_22_r;
wire signed [`OutBus]		out_28_22_i;
wire signed [`OutBus]		out_28_23_r;
wire signed [`OutBus]		out_28_23_i;
wire signed [`OutBus]		out_28_24_r;
wire signed [`OutBus]		out_28_24_i;
wire signed [`OutBus]		out_28_25_r;
wire signed [`OutBus]		out_28_25_i;
wire signed [`OutBus]		out_28_26_r;
wire signed [`OutBus]		out_28_26_i;
wire signed [`OutBus]		out_28_27_r;
wire signed [`OutBus]		out_28_27_i;
wire signed [`OutBus]		out_28_28_r;
wire signed [`OutBus]		out_28_28_i;
wire signed [`OutBus]		out_28_29_r;
wire signed [`OutBus]		out_28_29_i;
wire signed [`OutBus]		out_28_30_r;
wire signed [`OutBus]		out_28_30_i;
wire signed [`OutBus]		out_28_31_r;
wire signed [`OutBus]		out_28_31_i;
wire signed [`OutBus]		out_28_32_r;
wire signed [`OutBus]		out_28_32_i;
wire signed [`OutBus]		out_29_1_r;
wire signed [`OutBus]		out_29_1_i;
wire signed [`OutBus]		out_29_2_r;
wire signed [`OutBus]		out_29_2_i;
wire signed [`OutBus]		out_29_3_r;
wire signed [`OutBus]		out_29_3_i;
wire signed [`OutBus]		out_29_4_r;
wire signed [`OutBus]		out_29_4_i;
wire signed [`OutBus]		out_29_5_r;
wire signed [`OutBus]		out_29_5_i;
wire signed [`OutBus]		out_29_6_r;
wire signed [`OutBus]		out_29_6_i;
wire signed [`OutBus]		out_29_7_r;
wire signed [`OutBus]		out_29_7_i;
wire signed [`OutBus]		out_29_8_r;
wire signed [`OutBus]		out_29_8_i;
wire signed [`OutBus]		out_29_9_r;
wire signed [`OutBus]		out_29_9_i;
wire signed [`OutBus]		out_29_10_r;
wire signed [`OutBus]		out_29_10_i;
wire signed [`OutBus]		out_29_11_r;
wire signed [`OutBus]		out_29_11_i;
wire signed [`OutBus]		out_29_12_r;
wire signed [`OutBus]		out_29_12_i;
wire signed [`OutBus]		out_29_13_r;
wire signed [`OutBus]		out_29_13_i;
wire signed [`OutBus]		out_29_14_r;
wire signed [`OutBus]		out_29_14_i;
wire signed [`OutBus]		out_29_15_r;
wire signed [`OutBus]		out_29_15_i;
wire signed [`OutBus]		out_29_16_r;
wire signed [`OutBus]		out_29_16_i;
wire signed [`OutBus]		out_29_17_r;
wire signed [`OutBus]		out_29_17_i;
wire signed [`OutBus]		out_29_18_r;
wire signed [`OutBus]		out_29_18_i;
wire signed [`OutBus]		out_29_19_r;
wire signed [`OutBus]		out_29_19_i;
wire signed [`OutBus]		out_29_20_r;
wire signed [`OutBus]		out_29_20_i;
wire signed [`OutBus]		out_29_21_r;
wire signed [`OutBus]		out_29_21_i;
wire signed [`OutBus]		out_29_22_r;
wire signed [`OutBus]		out_29_22_i;
wire signed [`OutBus]		out_29_23_r;
wire signed [`OutBus]		out_29_23_i;
wire signed [`OutBus]		out_29_24_r;
wire signed [`OutBus]		out_29_24_i;
wire signed [`OutBus]		out_29_25_r;
wire signed [`OutBus]		out_29_25_i;
wire signed [`OutBus]		out_29_26_r;
wire signed [`OutBus]		out_29_26_i;
wire signed [`OutBus]		out_29_27_r;
wire signed [`OutBus]		out_29_27_i;
wire signed [`OutBus]		out_29_28_r;
wire signed [`OutBus]		out_29_28_i;
wire signed [`OutBus]		out_29_29_r;
wire signed [`OutBus]		out_29_29_i;
wire signed [`OutBus]		out_29_30_r;
wire signed [`OutBus]		out_29_30_i;
wire signed [`OutBus]		out_29_31_r;
wire signed [`OutBus]		out_29_31_i;
wire signed [`OutBus]		out_29_32_r;
wire signed [`OutBus]		out_29_32_i;
wire signed [`OutBus]		out_30_1_r;
wire signed [`OutBus]		out_30_1_i;
wire signed [`OutBus]		out_30_2_r;
wire signed [`OutBus]		out_30_2_i;
wire signed [`OutBus]		out_30_3_r;
wire signed [`OutBus]		out_30_3_i;
wire signed [`OutBus]		out_30_4_r;
wire signed [`OutBus]		out_30_4_i;
wire signed [`OutBus]		out_30_5_r;
wire signed [`OutBus]		out_30_5_i;
wire signed [`OutBus]		out_30_6_r;
wire signed [`OutBus]		out_30_6_i;
wire signed [`OutBus]		out_30_7_r;
wire signed [`OutBus]		out_30_7_i;
wire signed [`OutBus]		out_30_8_r;
wire signed [`OutBus]		out_30_8_i;
wire signed [`OutBus]		out_30_9_r;
wire signed [`OutBus]		out_30_9_i;
wire signed [`OutBus]		out_30_10_r;
wire signed [`OutBus]		out_30_10_i;
wire signed [`OutBus]		out_30_11_r;
wire signed [`OutBus]		out_30_11_i;
wire signed [`OutBus]		out_30_12_r;
wire signed [`OutBus]		out_30_12_i;
wire signed [`OutBus]		out_30_13_r;
wire signed [`OutBus]		out_30_13_i;
wire signed [`OutBus]		out_30_14_r;
wire signed [`OutBus]		out_30_14_i;
wire signed [`OutBus]		out_30_15_r;
wire signed [`OutBus]		out_30_15_i;
wire signed [`OutBus]		out_30_16_r;
wire signed [`OutBus]		out_30_16_i;
wire signed [`OutBus]		out_30_17_r;
wire signed [`OutBus]		out_30_17_i;
wire signed [`OutBus]		out_30_18_r;
wire signed [`OutBus]		out_30_18_i;
wire signed [`OutBus]		out_30_19_r;
wire signed [`OutBus]		out_30_19_i;
wire signed [`OutBus]		out_30_20_r;
wire signed [`OutBus]		out_30_20_i;
wire signed [`OutBus]		out_30_21_r;
wire signed [`OutBus]		out_30_21_i;
wire signed [`OutBus]		out_30_22_r;
wire signed [`OutBus]		out_30_22_i;
wire signed [`OutBus]		out_30_23_r;
wire signed [`OutBus]		out_30_23_i;
wire signed [`OutBus]		out_30_24_r;
wire signed [`OutBus]		out_30_24_i;
wire signed [`OutBus]		out_30_25_r;
wire signed [`OutBus]		out_30_25_i;
wire signed [`OutBus]		out_30_26_r;
wire signed [`OutBus]		out_30_26_i;
wire signed [`OutBus]		out_30_27_r;
wire signed [`OutBus]		out_30_27_i;
wire signed [`OutBus]		out_30_28_r;
wire signed [`OutBus]		out_30_28_i;
wire signed [`OutBus]		out_30_29_r;
wire signed [`OutBus]		out_30_29_i;
wire signed [`OutBus]		out_30_30_r;
wire signed [`OutBus]		out_30_30_i;
wire signed [`OutBus]		out_30_31_r;
wire signed [`OutBus]		out_30_31_i;
wire signed [`OutBus]		out_30_32_r;
wire signed [`OutBus]		out_30_32_i;
wire signed [`OutBus]		out_31_1_r;
wire signed [`OutBus]		out_31_1_i;
wire signed [`OutBus]		out_31_2_r;
wire signed [`OutBus]		out_31_2_i;
wire signed [`OutBus]		out_31_3_r;
wire signed [`OutBus]		out_31_3_i;
wire signed [`OutBus]		out_31_4_r;
wire signed [`OutBus]		out_31_4_i;
wire signed [`OutBus]		out_31_5_r;
wire signed [`OutBus]		out_31_5_i;
wire signed [`OutBus]		out_31_6_r;
wire signed [`OutBus]		out_31_6_i;
wire signed [`OutBus]		out_31_7_r;
wire signed [`OutBus]		out_31_7_i;
wire signed [`OutBus]		out_31_8_r;
wire signed [`OutBus]		out_31_8_i;
wire signed [`OutBus]		out_31_9_r;
wire signed [`OutBus]		out_31_9_i;
wire signed [`OutBus]		out_31_10_r;
wire signed [`OutBus]		out_31_10_i;
wire signed [`OutBus]		out_31_11_r;
wire signed [`OutBus]		out_31_11_i;
wire signed [`OutBus]		out_31_12_r;
wire signed [`OutBus]		out_31_12_i;
wire signed [`OutBus]		out_31_13_r;
wire signed [`OutBus]		out_31_13_i;
wire signed [`OutBus]		out_31_14_r;
wire signed [`OutBus]		out_31_14_i;
wire signed [`OutBus]		out_31_15_r;
wire signed [`OutBus]		out_31_15_i;
wire signed [`OutBus]		out_31_16_r;
wire signed [`OutBus]		out_31_16_i;
wire signed [`OutBus]		out_31_17_r;
wire signed [`OutBus]		out_31_17_i;
wire signed [`OutBus]		out_31_18_r;
wire signed [`OutBus]		out_31_18_i;
wire signed [`OutBus]		out_31_19_r;
wire signed [`OutBus]		out_31_19_i;
wire signed [`OutBus]		out_31_20_r;
wire signed [`OutBus]		out_31_20_i;
wire signed [`OutBus]		out_31_21_r;
wire signed [`OutBus]		out_31_21_i;
wire signed [`OutBus]		out_31_22_r;
wire signed [`OutBus]		out_31_22_i;
wire signed [`OutBus]		out_31_23_r;
wire signed [`OutBus]		out_31_23_i;
wire signed [`OutBus]		out_31_24_r;
wire signed [`OutBus]		out_31_24_i;
wire signed [`OutBus]		out_31_25_r;
wire signed [`OutBus]		out_31_25_i;
wire signed [`OutBus]		out_31_26_r;
wire signed [`OutBus]		out_31_26_i;
wire signed [`OutBus]		out_31_27_r;
wire signed [`OutBus]		out_31_27_i;
wire signed [`OutBus]		out_31_28_r;
wire signed [`OutBus]		out_31_28_i;
wire signed [`OutBus]		out_31_29_r;
wire signed [`OutBus]		out_31_29_i;
wire signed [`OutBus]		out_31_30_r;
wire signed [`OutBus]		out_31_30_i;
wire signed [`OutBus]		out_31_31_r;
wire signed [`OutBus]		out_31_31_i;
wire signed [`OutBus]		out_31_32_r;
wire signed [`OutBus]		out_31_32_i;
wire signed [`OutBus]		out_32_1_r;
wire signed [`OutBus]		out_32_1_i;
wire signed [`OutBus]		out_32_2_r;
wire signed [`OutBus]		out_32_2_i;
wire signed [`OutBus]		out_32_3_r;
wire signed [`OutBus]		out_32_3_i;
wire signed [`OutBus]		out_32_4_r;
wire signed [`OutBus]		out_32_4_i;
wire signed [`OutBus]		out_32_5_r;
wire signed [`OutBus]		out_32_5_i;
wire signed [`OutBus]		out_32_6_r;
wire signed [`OutBus]		out_32_6_i;
wire signed [`OutBus]		out_32_7_r;
wire signed [`OutBus]		out_32_7_i;
wire signed [`OutBus]		out_32_8_r;
wire signed [`OutBus]		out_32_8_i;
wire signed [`OutBus]		out_32_9_r;
wire signed [`OutBus]		out_32_9_i;
wire signed [`OutBus]		out_32_10_r;
wire signed [`OutBus]		out_32_10_i;
wire signed [`OutBus]		out_32_11_r;
wire signed [`OutBus]		out_32_11_i;
wire signed [`OutBus]		out_32_12_r;
wire signed [`OutBus]		out_32_12_i;
wire signed [`OutBus]		out_32_13_r;
wire signed [`OutBus]		out_32_13_i;
wire signed [`OutBus]		out_32_14_r;
wire signed [`OutBus]		out_32_14_i;
wire signed [`OutBus]		out_32_15_r;
wire signed [`OutBus]		out_32_15_i;
wire signed [`OutBus]		out_32_16_r;
wire signed [`OutBus]		out_32_16_i;
wire signed [`OutBus]		out_32_17_r;
wire signed [`OutBus]		out_32_17_i;
wire signed [`OutBus]		out_32_18_r;
wire signed [`OutBus]		out_32_18_i;
wire signed [`OutBus]		out_32_19_r;
wire signed [`OutBus]		out_32_19_i;
wire signed [`OutBus]		out_32_20_r;
wire signed [`OutBus]		out_32_20_i;
wire signed [`OutBus]		out_32_21_r;
wire signed [`OutBus]		out_32_21_i;
wire signed [`OutBus]		out_32_22_r;
wire signed [`OutBus]		out_32_22_i;
wire signed [`OutBus]		out_32_23_r;
wire signed [`OutBus]		out_32_23_i;
wire signed [`OutBus]		out_32_24_r;
wire signed [`OutBus]		out_32_24_i;
wire signed [`OutBus]		out_32_25_r;
wire signed [`OutBus]		out_32_25_i;
wire signed [`OutBus]		out_32_26_r;
wire signed [`OutBus]		out_32_26_i;
wire signed [`OutBus]		out_32_27_r;
wire signed [`OutBus]		out_32_27_i;
wire signed [`OutBus]		out_32_28_r;
wire signed [`OutBus]		out_32_28_i;
wire signed [`OutBus]		out_32_29_r;
wire signed [`OutBus]		out_32_29_i;
wire signed [`OutBus]		out_32_30_r;
wire signed [`OutBus]		out_32_30_i;
wire signed [`OutBus]		out_32_31_r;
wire signed [`OutBus]		out_32_31_i;
wire signed [`OutBus]		out_32_32_r;
wire signed [`OutBus]		out_32_32_i;

/************************temp MUX butterfly***********************/
wire signed [`CalcTempBus]          temp_m1_1_1_r;
wire signed [`CalcTempBus]          temp_m1_1_1_i;
wire signed [`CalcTempBus]          temp_m1_1_2_r;
wire signed [`CalcTempBus]          temp_m1_1_2_i;
wire signed [`CalcTempBus]          temp_m1_1_3_r;
wire signed [`CalcTempBus]          temp_m1_1_3_i;
wire signed [`CalcTempBus]          temp_m1_1_4_r;
wire signed [`CalcTempBus]          temp_m1_1_4_i;
wire signed [`CalcTempBus]          temp_m1_1_5_r;
wire signed [`CalcTempBus]          temp_m1_1_5_i;
wire signed [`CalcTempBus]          temp_m1_1_6_r;
wire signed [`CalcTempBus]          temp_m1_1_6_i;
wire signed [`CalcTempBus]          temp_m1_1_7_r;
wire signed [`CalcTempBus]          temp_m1_1_7_i;
wire signed [`CalcTempBus]          temp_m1_1_8_r;
wire signed [`CalcTempBus]          temp_m1_1_8_i;
wire signed [`CalcTempBus]          temp_m1_1_9_r;
wire signed [`CalcTempBus]          temp_m1_1_9_i;
wire signed [`CalcTempBus]          temp_m1_1_10_r;
wire signed [`CalcTempBus]          temp_m1_1_10_i;
wire signed [`CalcTempBus]          temp_m1_1_11_r;
wire signed [`CalcTempBus]          temp_m1_1_11_i;
wire signed [`CalcTempBus]          temp_m1_1_12_r;
wire signed [`CalcTempBus]          temp_m1_1_12_i;
wire signed [`CalcTempBus]          temp_m1_1_13_r;
wire signed [`CalcTempBus]          temp_m1_1_13_i;
wire signed [`CalcTempBus]          temp_m1_1_14_r;
wire signed [`CalcTempBus]          temp_m1_1_14_i;
wire signed [`CalcTempBus]          temp_m1_1_15_r;
wire signed [`CalcTempBus]          temp_m1_1_15_i;
wire signed [`CalcTempBus]          temp_m1_1_16_r;
wire signed [`CalcTempBus]          temp_m1_1_16_i;
wire signed [`CalcTempBus]          temp_m1_1_17_r;
wire signed [`CalcTempBus]          temp_m1_1_17_i;
wire signed [`CalcTempBus]          temp_m1_1_18_r;
wire signed [`CalcTempBus]          temp_m1_1_18_i;
wire signed [`CalcTempBus]          temp_m1_1_19_r;
wire signed [`CalcTempBus]          temp_m1_1_19_i;
wire signed [`CalcTempBus]          temp_m1_1_20_r;
wire signed [`CalcTempBus]          temp_m1_1_20_i;
wire signed [`CalcTempBus]          temp_m1_1_21_r;
wire signed [`CalcTempBus]          temp_m1_1_21_i;
wire signed [`CalcTempBus]          temp_m1_1_22_r;
wire signed [`CalcTempBus]          temp_m1_1_22_i;
wire signed [`CalcTempBus]          temp_m1_1_23_r;
wire signed [`CalcTempBus]          temp_m1_1_23_i;
wire signed [`CalcTempBus]          temp_m1_1_24_r;
wire signed [`CalcTempBus]          temp_m1_1_24_i;
wire signed [`CalcTempBus]          temp_m1_1_25_r;
wire signed [`CalcTempBus]          temp_m1_1_25_i;
wire signed [`CalcTempBus]          temp_m1_1_26_r;
wire signed [`CalcTempBus]          temp_m1_1_26_i;
wire signed [`CalcTempBus]          temp_m1_1_27_r;
wire signed [`CalcTempBus]          temp_m1_1_27_i;
wire signed [`CalcTempBus]          temp_m1_1_28_r;
wire signed [`CalcTempBus]          temp_m1_1_28_i;
wire signed [`CalcTempBus]          temp_m1_1_29_r;
wire signed [`CalcTempBus]          temp_m1_1_29_i;
wire signed [`CalcTempBus]          temp_m1_1_30_r;
wire signed [`CalcTempBus]          temp_m1_1_30_i;
wire signed [`CalcTempBus]          temp_m1_1_31_r;
wire signed [`CalcTempBus]          temp_m1_1_31_i;
wire signed [`CalcTempBus]          temp_m1_1_32_r;
wire signed [`CalcTempBus]          temp_m1_1_32_i;
wire signed [`CalcTempBus]          temp_m1_2_1_r;
wire signed [`CalcTempBus]          temp_m1_2_1_i;
wire signed [`CalcTempBus]          temp_m1_2_2_r;
wire signed [`CalcTempBus]          temp_m1_2_2_i;
wire signed [`CalcTempBus]          temp_m1_2_3_r;
wire signed [`CalcTempBus]          temp_m1_2_3_i;
wire signed [`CalcTempBus]          temp_m1_2_4_r;
wire signed [`CalcTempBus]          temp_m1_2_4_i;
wire signed [`CalcTempBus]          temp_m1_2_5_r;
wire signed [`CalcTempBus]          temp_m1_2_5_i;
wire signed [`CalcTempBus]          temp_m1_2_6_r;
wire signed [`CalcTempBus]          temp_m1_2_6_i;
wire signed [`CalcTempBus]          temp_m1_2_7_r;
wire signed [`CalcTempBus]          temp_m1_2_7_i;
wire signed [`CalcTempBus]          temp_m1_2_8_r;
wire signed [`CalcTempBus]          temp_m1_2_8_i;
wire signed [`CalcTempBus]          temp_m1_2_9_r;
wire signed [`CalcTempBus]          temp_m1_2_9_i;
wire signed [`CalcTempBus]          temp_m1_2_10_r;
wire signed [`CalcTempBus]          temp_m1_2_10_i;
wire signed [`CalcTempBus]          temp_m1_2_11_r;
wire signed [`CalcTempBus]          temp_m1_2_11_i;
wire signed [`CalcTempBus]          temp_m1_2_12_r;
wire signed [`CalcTempBus]          temp_m1_2_12_i;
wire signed [`CalcTempBus]          temp_m1_2_13_r;
wire signed [`CalcTempBus]          temp_m1_2_13_i;
wire signed [`CalcTempBus]          temp_m1_2_14_r;
wire signed [`CalcTempBus]          temp_m1_2_14_i;
wire signed [`CalcTempBus]          temp_m1_2_15_r;
wire signed [`CalcTempBus]          temp_m1_2_15_i;
wire signed [`CalcTempBus]          temp_m1_2_16_r;
wire signed [`CalcTempBus]          temp_m1_2_16_i;
wire signed [`CalcTempBus]          temp_m1_2_17_r;
wire signed [`CalcTempBus]          temp_m1_2_17_i;
wire signed [`CalcTempBus]          temp_m1_2_18_r;
wire signed [`CalcTempBus]          temp_m1_2_18_i;
wire signed [`CalcTempBus]          temp_m1_2_19_r;
wire signed [`CalcTempBus]          temp_m1_2_19_i;
wire signed [`CalcTempBus]          temp_m1_2_20_r;
wire signed [`CalcTempBus]          temp_m1_2_20_i;
wire signed [`CalcTempBus]          temp_m1_2_21_r;
wire signed [`CalcTempBus]          temp_m1_2_21_i;
wire signed [`CalcTempBus]          temp_m1_2_22_r;
wire signed [`CalcTempBus]          temp_m1_2_22_i;
wire signed [`CalcTempBus]          temp_m1_2_23_r;
wire signed [`CalcTempBus]          temp_m1_2_23_i;
wire signed [`CalcTempBus]          temp_m1_2_24_r;
wire signed [`CalcTempBus]          temp_m1_2_24_i;
wire signed [`CalcTempBus]          temp_m1_2_25_r;
wire signed [`CalcTempBus]          temp_m1_2_25_i;
wire signed [`CalcTempBus]          temp_m1_2_26_r;
wire signed [`CalcTempBus]          temp_m1_2_26_i;
wire signed [`CalcTempBus]          temp_m1_2_27_r;
wire signed [`CalcTempBus]          temp_m1_2_27_i;
wire signed [`CalcTempBus]          temp_m1_2_28_r;
wire signed [`CalcTempBus]          temp_m1_2_28_i;
wire signed [`CalcTempBus]          temp_m1_2_29_r;
wire signed [`CalcTempBus]          temp_m1_2_29_i;
wire signed [`CalcTempBus]          temp_m1_2_30_r;
wire signed [`CalcTempBus]          temp_m1_2_30_i;
wire signed [`CalcTempBus]          temp_m1_2_31_r;
wire signed [`CalcTempBus]          temp_m1_2_31_i;
wire signed [`CalcTempBus]          temp_m1_2_32_r;
wire signed [`CalcTempBus]          temp_m1_2_32_i;
wire signed [`CalcTempBus]          temp_m1_3_1_r;
wire signed [`CalcTempBus]          temp_m1_3_1_i;
wire signed [`CalcTempBus]          temp_m1_3_2_r;
wire signed [`CalcTempBus]          temp_m1_3_2_i;
wire signed [`CalcTempBus]          temp_m1_3_3_r;
wire signed [`CalcTempBus]          temp_m1_3_3_i;
wire signed [`CalcTempBus]          temp_m1_3_4_r;
wire signed [`CalcTempBus]          temp_m1_3_4_i;
wire signed [`CalcTempBus]          temp_m1_3_5_r;
wire signed [`CalcTempBus]          temp_m1_3_5_i;
wire signed [`CalcTempBus]          temp_m1_3_6_r;
wire signed [`CalcTempBus]          temp_m1_3_6_i;
wire signed [`CalcTempBus]          temp_m1_3_7_r;
wire signed [`CalcTempBus]          temp_m1_3_7_i;
wire signed [`CalcTempBus]          temp_m1_3_8_r;
wire signed [`CalcTempBus]          temp_m1_3_8_i;
wire signed [`CalcTempBus]          temp_m1_3_9_r;
wire signed [`CalcTempBus]          temp_m1_3_9_i;
wire signed [`CalcTempBus]          temp_m1_3_10_r;
wire signed [`CalcTempBus]          temp_m1_3_10_i;
wire signed [`CalcTempBus]          temp_m1_3_11_r;
wire signed [`CalcTempBus]          temp_m1_3_11_i;
wire signed [`CalcTempBus]          temp_m1_3_12_r;
wire signed [`CalcTempBus]          temp_m1_3_12_i;
wire signed [`CalcTempBus]          temp_m1_3_13_r;
wire signed [`CalcTempBus]          temp_m1_3_13_i;
wire signed [`CalcTempBus]          temp_m1_3_14_r;
wire signed [`CalcTempBus]          temp_m1_3_14_i;
wire signed [`CalcTempBus]          temp_m1_3_15_r;
wire signed [`CalcTempBus]          temp_m1_3_15_i;
wire signed [`CalcTempBus]          temp_m1_3_16_r;
wire signed [`CalcTempBus]          temp_m1_3_16_i;
wire signed [`CalcTempBus]          temp_m1_3_17_r;
wire signed [`CalcTempBus]          temp_m1_3_17_i;
wire signed [`CalcTempBus]          temp_m1_3_18_r;
wire signed [`CalcTempBus]          temp_m1_3_18_i;
wire signed [`CalcTempBus]          temp_m1_3_19_r;
wire signed [`CalcTempBus]          temp_m1_3_19_i;
wire signed [`CalcTempBus]          temp_m1_3_20_r;
wire signed [`CalcTempBus]          temp_m1_3_20_i;
wire signed [`CalcTempBus]          temp_m1_3_21_r;
wire signed [`CalcTempBus]          temp_m1_3_21_i;
wire signed [`CalcTempBus]          temp_m1_3_22_r;
wire signed [`CalcTempBus]          temp_m1_3_22_i;
wire signed [`CalcTempBus]          temp_m1_3_23_r;
wire signed [`CalcTempBus]          temp_m1_3_23_i;
wire signed [`CalcTempBus]          temp_m1_3_24_r;
wire signed [`CalcTempBus]          temp_m1_3_24_i;
wire signed [`CalcTempBus]          temp_m1_3_25_r;
wire signed [`CalcTempBus]          temp_m1_3_25_i;
wire signed [`CalcTempBus]          temp_m1_3_26_r;
wire signed [`CalcTempBus]          temp_m1_3_26_i;
wire signed [`CalcTempBus]          temp_m1_3_27_r;
wire signed [`CalcTempBus]          temp_m1_3_27_i;
wire signed [`CalcTempBus]          temp_m1_3_28_r;
wire signed [`CalcTempBus]          temp_m1_3_28_i;
wire signed [`CalcTempBus]          temp_m1_3_29_r;
wire signed [`CalcTempBus]          temp_m1_3_29_i;
wire signed [`CalcTempBus]          temp_m1_3_30_r;
wire signed [`CalcTempBus]          temp_m1_3_30_i;
wire signed [`CalcTempBus]          temp_m1_3_31_r;
wire signed [`CalcTempBus]          temp_m1_3_31_i;
wire signed [`CalcTempBus]          temp_m1_3_32_r;
wire signed [`CalcTempBus]          temp_m1_3_32_i;
wire signed [`CalcTempBus]          temp_m1_4_1_r;
wire signed [`CalcTempBus]          temp_m1_4_1_i;
wire signed [`CalcTempBus]          temp_m1_4_2_r;
wire signed [`CalcTempBus]          temp_m1_4_2_i;
wire signed [`CalcTempBus]          temp_m1_4_3_r;
wire signed [`CalcTempBus]          temp_m1_4_3_i;
wire signed [`CalcTempBus]          temp_m1_4_4_r;
wire signed [`CalcTempBus]          temp_m1_4_4_i;
wire signed [`CalcTempBus]          temp_m1_4_5_r;
wire signed [`CalcTempBus]          temp_m1_4_5_i;
wire signed [`CalcTempBus]          temp_m1_4_6_r;
wire signed [`CalcTempBus]          temp_m1_4_6_i;
wire signed [`CalcTempBus]          temp_m1_4_7_r;
wire signed [`CalcTempBus]          temp_m1_4_7_i;
wire signed [`CalcTempBus]          temp_m1_4_8_r;
wire signed [`CalcTempBus]          temp_m1_4_8_i;
wire signed [`CalcTempBus]          temp_m1_4_9_r;
wire signed [`CalcTempBus]          temp_m1_4_9_i;
wire signed [`CalcTempBus]          temp_m1_4_10_r;
wire signed [`CalcTempBus]          temp_m1_4_10_i;
wire signed [`CalcTempBus]          temp_m1_4_11_r;
wire signed [`CalcTempBus]          temp_m1_4_11_i;
wire signed [`CalcTempBus]          temp_m1_4_12_r;
wire signed [`CalcTempBus]          temp_m1_4_12_i;
wire signed [`CalcTempBus]          temp_m1_4_13_r;
wire signed [`CalcTempBus]          temp_m1_4_13_i;
wire signed [`CalcTempBus]          temp_m1_4_14_r;
wire signed [`CalcTempBus]          temp_m1_4_14_i;
wire signed [`CalcTempBus]          temp_m1_4_15_r;
wire signed [`CalcTempBus]          temp_m1_4_15_i;
wire signed [`CalcTempBus]          temp_m1_4_16_r;
wire signed [`CalcTempBus]          temp_m1_4_16_i;
wire signed [`CalcTempBus]          temp_m1_4_17_r;
wire signed [`CalcTempBus]          temp_m1_4_17_i;
wire signed [`CalcTempBus]          temp_m1_4_18_r;
wire signed [`CalcTempBus]          temp_m1_4_18_i;
wire signed [`CalcTempBus]          temp_m1_4_19_r;
wire signed [`CalcTempBus]          temp_m1_4_19_i;
wire signed [`CalcTempBus]          temp_m1_4_20_r;
wire signed [`CalcTempBus]          temp_m1_4_20_i;
wire signed [`CalcTempBus]          temp_m1_4_21_r;
wire signed [`CalcTempBus]          temp_m1_4_21_i;
wire signed [`CalcTempBus]          temp_m1_4_22_r;
wire signed [`CalcTempBus]          temp_m1_4_22_i;
wire signed [`CalcTempBus]          temp_m1_4_23_r;
wire signed [`CalcTempBus]          temp_m1_4_23_i;
wire signed [`CalcTempBus]          temp_m1_4_24_r;
wire signed [`CalcTempBus]          temp_m1_4_24_i;
wire signed [`CalcTempBus]          temp_m1_4_25_r;
wire signed [`CalcTempBus]          temp_m1_4_25_i;
wire signed [`CalcTempBus]          temp_m1_4_26_r;
wire signed [`CalcTempBus]          temp_m1_4_26_i;
wire signed [`CalcTempBus]          temp_m1_4_27_r;
wire signed [`CalcTempBus]          temp_m1_4_27_i;
wire signed [`CalcTempBus]          temp_m1_4_28_r;
wire signed [`CalcTempBus]          temp_m1_4_28_i;
wire signed [`CalcTempBus]          temp_m1_4_29_r;
wire signed [`CalcTempBus]          temp_m1_4_29_i;
wire signed [`CalcTempBus]          temp_m1_4_30_r;
wire signed [`CalcTempBus]          temp_m1_4_30_i;
wire signed [`CalcTempBus]          temp_m1_4_31_r;
wire signed [`CalcTempBus]          temp_m1_4_31_i;
wire signed [`CalcTempBus]          temp_m1_4_32_r;
wire signed [`CalcTempBus]          temp_m1_4_32_i;
wire signed [`CalcTempBus]          temp_m1_5_1_r;
wire signed [`CalcTempBus]          temp_m1_5_1_i;
wire signed [`CalcTempBus]          temp_m1_5_2_r;
wire signed [`CalcTempBus]          temp_m1_5_2_i;
wire signed [`CalcTempBus]          temp_m1_5_3_r;
wire signed [`CalcTempBus]          temp_m1_5_3_i;
wire signed [`CalcTempBus]          temp_m1_5_4_r;
wire signed [`CalcTempBus]          temp_m1_5_4_i;
wire signed [`CalcTempBus]          temp_m1_5_5_r;
wire signed [`CalcTempBus]          temp_m1_5_5_i;
wire signed [`CalcTempBus]          temp_m1_5_6_r;
wire signed [`CalcTempBus]          temp_m1_5_6_i;
wire signed [`CalcTempBus]          temp_m1_5_7_r;
wire signed [`CalcTempBus]          temp_m1_5_7_i;
wire signed [`CalcTempBus]          temp_m1_5_8_r;
wire signed [`CalcTempBus]          temp_m1_5_8_i;
wire signed [`CalcTempBus]          temp_m1_5_9_r;
wire signed [`CalcTempBus]          temp_m1_5_9_i;
wire signed [`CalcTempBus]          temp_m1_5_10_r;
wire signed [`CalcTempBus]          temp_m1_5_10_i;
wire signed [`CalcTempBus]          temp_m1_5_11_r;
wire signed [`CalcTempBus]          temp_m1_5_11_i;
wire signed [`CalcTempBus]          temp_m1_5_12_r;
wire signed [`CalcTempBus]          temp_m1_5_12_i;
wire signed [`CalcTempBus]          temp_m1_5_13_r;
wire signed [`CalcTempBus]          temp_m1_5_13_i;
wire signed [`CalcTempBus]          temp_m1_5_14_r;
wire signed [`CalcTempBus]          temp_m1_5_14_i;
wire signed [`CalcTempBus]          temp_m1_5_15_r;
wire signed [`CalcTempBus]          temp_m1_5_15_i;
wire signed [`CalcTempBus]          temp_m1_5_16_r;
wire signed [`CalcTempBus]          temp_m1_5_16_i;
wire signed [`CalcTempBus]          temp_m1_5_17_r;
wire signed [`CalcTempBus]          temp_m1_5_17_i;
wire signed [`CalcTempBus]          temp_m1_5_18_r;
wire signed [`CalcTempBus]          temp_m1_5_18_i;
wire signed [`CalcTempBus]          temp_m1_5_19_r;
wire signed [`CalcTempBus]          temp_m1_5_19_i;
wire signed [`CalcTempBus]          temp_m1_5_20_r;
wire signed [`CalcTempBus]          temp_m1_5_20_i;
wire signed [`CalcTempBus]          temp_m1_5_21_r;
wire signed [`CalcTempBus]          temp_m1_5_21_i;
wire signed [`CalcTempBus]          temp_m1_5_22_r;
wire signed [`CalcTempBus]          temp_m1_5_22_i;
wire signed [`CalcTempBus]          temp_m1_5_23_r;
wire signed [`CalcTempBus]          temp_m1_5_23_i;
wire signed [`CalcTempBus]          temp_m1_5_24_r;
wire signed [`CalcTempBus]          temp_m1_5_24_i;
wire signed [`CalcTempBus]          temp_m1_5_25_r;
wire signed [`CalcTempBus]          temp_m1_5_25_i;
wire signed [`CalcTempBus]          temp_m1_5_26_r;
wire signed [`CalcTempBus]          temp_m1_5_26_i;
wire signed [`CalcTempBus]          temp_m1_5_27_r;
wire signed [`CalcTempBus]          temp_m1_5_27_i;
wire signed [`CalcTempBus]          temp_m1_5_28_r;
wire signed [`CalcTempBus]          temp_m1_5_28_i;
wire signed [`CalcTempBus]          temp_m1_5_29_r;
wire signed [`CalcTempBus]          temp_m1_5_29_i;
wire signed [`CalcTempBus]          temp_m1_5_30_r;
wire signed [`CalcTempBus]          temp_m1_5_30_i;
wire signed [`CalcTempBus]          temp_m1_5_31_r;
wire signed [`CalcTempBus]          temp_m1_5_31_i;
wire signed [`CalcTempBus]          temp_m1_5_32_r;
wire signed [`CalcTempBus]          temp_m1_5_32_i;
wire signed [`CalcTempBus]          temp_m1_6_1_r;
wire signed [`CalcTempBus]          temp_m1_6_1_i;
wire signed [`CalcTempBus]          temp_m1_6_2_r;
wire signed [`CalcTempBus]          temp_m1_6_2_i;
wire signed [`CalcTempBus]          temp_m1_6_3_r;
wire signed [`CalcTempBus]          temp_m1_6_3_i;
wire signed [`CalcTempBus]          temp_m1_6_4_r;
wire signed [`CalcTempBus]          temp_m1_6_4_i;
wire signed [`CalcTempBus]          temp_m1_6_5_r;
wire signed [`CalcTempBus]          temp_m1_6_5_i;
wire signed [`CalcTempBus]          temp_m1_6_6_r;
wire signed [`CalcTempBus]          temp_m1_6_6_i;
wire signed [`CalcTempBus]          temp_m1_6_7_r;
wire signed [`CalcTempBus]          temp_m1_6_7_i;
wire signed [`CalcTempBus]          temp_m1_6_8_r;
wire signed [`CalcTempBus]          temp_m1_6_8_i;
wire signed [`CalcTempBus]          temp_m1_6_9_r;
wire signed [`CalcTempBus]          temp_m1_6_9_i;
wire signed [`CalcTempBus]          temp_m1_6_10_r;
wire signed [`CalcTempBus]          temp_m1_6_10_i;
wire signed [`CalcTempBus]          temp_m1_6_11_r;
wire signed [`CalcTempBus]          temp_m1_6_11_i;
wire signed [`CalcTempBus]          temp_m1_6_12_r;
wire signed [`CalcTempBus]          temp_m1_6_12_i;
wire signed [`CalcTempBus]          temp_m1_6_13_r;
wire signed [`CalcTempBus]          temp_m1_6_13_i;
wire signed [`CalcTempBus]          temp_m1_6_14_r;
wire signed [`CalcTempBus]          temp_m1_6_14_i;
wire signed [`CalcTempBus]          temp_m1_6_15_r;
wire signed [`CalcTempBus]          temp_m1_6_15_i;
wire signed [`CalcTempBus]          temp_m1_6_16_r;
wire signed [`CalcTempBus]          temp_m1_6_16_i;
wire signed [`CalcTempBus]          temp_m1_6_17_r;
wire signed [`CalcTempBus]          temp_m1_6_17_i;
wire signed [`CalcTempBus]          temp_m1_6_18_r;
wire signed [`CalcTempBus]          temp_m1_6_18_i;
wire signed [`CalcTempBus]          temp_m1_6_19_r;
wire signed [`CalcTempBus]          temp_m1_6_19_i;
wire signed [`CalcTempBus]          temp_m1_6_20_r;
wire signed [`CalcTempBus]          temp_m1_6_20_i;
wire signed [`CalcTempBus]          temp_m1_6_21_r;
wire signed [`CalcTempBus]          temp_m1_6_21_i;
wire signed [`CalcTempBus]          temp_m1_6_22_r;
wire signed [`CalcTempBus]          temp_m1_6_22_i;
wire signed [`CalcTempBus]          temp_m1_6_23_r;
wire signed [`CalcTempBus]          temp_m1_6_23_i;
wire signed [`CalcTempBus]          temp_m1_6_24_r;
wire signed [`CalcTempBus]          temp_m1_6_24_i;
wire signed [`CalcTempBus]          temp_m1_6_25_r;
wire signed [`CalcTempBus]          temp_m1_6_25_i;
wire signed [`CalcTempBus]          temp_m1_6_26_r;
wire signed [`CalcTempBus]          temp_m1_6_26_i;
wire signed [`CalcTempBus]          temp_m1_6_27_r;
wire signed [`CalcTempBus]          temp_m1_6_27_i;
wire signed [`CalcTempBus]          temp_m1_6_28_r;
wire signed [`CalcTempBus]          temp_m1_6_28_i;
wire signed [`CalcTempBus]          temp_m1_6_29_r;
wire signed [`CalcTempBus]          temp_m1_6_29_i;
wire signed [`CalcTempBus]          temp_m1_6_30_r;
wire signed [`CalcTempBus]          temp_m1_6_30_i;
wire signed [`CalcTempBus]          temp_m1_6_31_r;
wire signed [`CalcTempBus]          temp_m1_6_31_i;
wire signed [`CalcTempBus]          temp_m1_6_32_r;
wire signed [`CalcTempBus]          temp_m1_6_32_i;
wire signed [`CalcTempBus]          temp_m1_7_1_r;
wire signed [`CalcTempBus]          temp_m1_7_1_i;
wire signed [`CalcTempBus]          temp_m1_7_2_r;
wire signed [`CalcTempBus]          temp_m1_7_2_i;
wire signed [`CalcTempBus]          temp_m1_7_3_r;
wire signed [`CalcTempBus]          temp_m1_7_3_i;
wire signed [`CalcTempBus]          temp_m1_7_4_r;
wire signed [`CalcTempBus]          temp_m1_7_4_i;
wire signed [`CalcTempBus]          temp_m1_7_5_r;
wire signed [`CalcTempBus]          temp_m1_7_5_i;
wire signed [`CalcTempBus]          temp_m1_7_6_r;
wire signed [`CalcTempBus]          temp_m1_7_6_i;
wire signed [`CalcTempBus]          temp_m1_7_7_r;
wire signed [`CalcTempBus]          temp_m1_7_7_i;
wire signed [`CalcTempBus]          temp_m1_7_8_r;
wire signed [`CalcTempBus]          temp_m1_7_8_i;
wire signed [`CalcTempBus]          temp_m1_7_9_r;
wire signed [`CalcTempBus]          temp_m1_7_9_i;
wire signed [`CalcTempBus]          temp_m1_7_10_r;
wire signed [`CalcTempBus]          temp_m1_7_10_i;
wire signed [`CalcTempBus]          temp_m1_7_11_r;
wire signed [`CalcTempBus]          temp_m1_7_11_i;
wire signed [`CalcTempBus]          temp_m1_7_12_r;
wire signed [`CalcTempBus]          temp_m1_7_12_i;
wire signed [`CalcTempBus]          temp_m1_7_13_r;
wire signed [`CalcTempBus]          temp_m1_7_13_i;
wire signed [`CalcTempBus]          temp_m1_7_14_r;
wire signed [`CalcTempBus]          temp_m1_7_14_i;
wire signed [`CalcTempBus]          temp_m1_7_15_r;
wire signed [`CalcTempBus]          temp_m1_7_15_i;
wire signed [`CalcTempBus]          temp_m1_7_16_r;
wire signed [`CalcTempBus]          temp_m1_7_16_i;
wire signed [`CalcTempBus]          temp_m1_7_17_r;
wire signed [`CalcTempBus]          temp_m1_7_17_i;
wire signed [`CalcTempBus]          temp_m1_7_18_r;
wire signed [`CalcTempBus]          temp_m1_7_18_i;
wire signed [`CalcTempBus]          temp_m1_7_19_r;
wire signed [`CalcTempBus]          temp_m1_7_19_i;
wire signed [`CalcTempBus]          temp_m1_7_20_r;
wire signed [`CalcTempBus]          temp_m1_7_20_i;
wire signed [`CalcTempBus]          temp_m1_7_21_r;
wire signed [`CalcTempBus]          temp_m1_7_21_i;
wire signed [`CalcTempBus]          temp_m1_7_22_r;
wire signed [`CalcTempBus]          temp_m1_7_22_i;
wire signed [`CalcTempBus]          temp_m1_7_23_r;
wire signed [`CalcTempBus]          temp_m1_7_23_i;
wire signed [`CalcTempBus]          temp_m1_7_24_r;
wire signed [`CalcTempBus]          temp_m1_7_24_i;
wire signed [`CalcTempBus]          temp_m1_7_25_r;
wire signed [`CalcTempBus]          temp_m1_7_25_i;
wire signed [`CalcTempBus]          temp_m1_7_26_r;
wire signed [`CalcTempBus]          temp_m1_7_26_i;
wire signed [`CalcTempBus]          temp_m1_7_27_r;
wire signed [`CalcTempBus]          temp_m1_7_27_i;
wire signed [`CalcTempBus]          temp_m1_7_28_r;
wire signed [`CalcTempBus]          temp_m1_7_28_i;
wire signed [`CalcTempBus]          temp_m1_7_29_r;
wire signed [`CalcTempBus]          temp_m1_7_29_i;
wire signed [`CalcTempBus]          temp_m1_7_30_r;
wire signed [`CalcTempBus]          temp_m1_7_30_i;
wire signed [`CalcTempBus]          temp_m1_7_31_r;
wire signed [`CalcTempBus]          temp_m1_7_31_i;
wire signed [`CalcTempBus]          temp_m1_7_32_r;
wire signed [`CalcTempBus]          temp_m1_7_32_i;
wire signed [`CalcTempBus]          temp_m1_8_1_r;
wire signed [`CalcTempBus]          temp_m1_8_1_i;
wire signed [`CalcTempBus]          temp_m1_8_2_r;
wire signed [`CalcTempBus]          temp_m1_8_2_i;
wire signed [`CalcTempBus]          temp_m1_8_3_r;
wire signed [`CalcTempBus]          temp_m1_8_3_i;
wire signed [`CalcTempBus]          temp_m1_8_4_r;
wire signed [`CalcTempBus]          temp_m1_8_4_i;
wire signed [`CalcTempBus]          temp_m1_8_5_r;
wire signed [`CalcTempBus]          temp_m1_8_5_i;
wire signed [`CalcTempBus]          temp_m1_8_6_r;
wire signed [`CalcTempBus]          temp_m1_8_6_i;
wire signed [`CalcTempBus]          temp_m1_8_7_r;
wire signed [`CalcTempBus]          temp_m1_8_7_i;
wire signed [`CalcTempBus]          temp_m1_8_8_r;
wire signed [`CalcTempBus]          temp_m1_8_8_i;
wire signed [`CalcTempBus]          temp_m1_8_9_r;
wire signed [`CalcTempBus]          temp_m1_8_9_i;
wire signed [`CalcTempBus]          temp_m1_8_10_r;
wire signed [`CalcTempBus]          temp_m1_8_10_i;
wire signed [`CalcTempBus]          temp_m1_8_11_r;
wire signed [`CalcTempBus]          temp_m1_8_11_i;
wire signed [`CalcTempBus]          temp_m1_8_12_r;
wire signed [`CalcTempBus]          temp_m1_8_12_i;
wire signed [`CalcTempBus]          temp_m1_8_13_r;
wire signed [`CalcTempBus]          temp_m1_8_13_i;
wire signed [`CalcTempBus]          temp_m1_8_14_r;
wire signed [`CalcTempBus]          temp_m1_8_14_i;
wire signed [`CalcTempBus]          temp_m1_8_15_r;
wire signed [`CalcTempBus]          temp_m1_8_15_i;
wire signed [`CalcTempBus]          temp_m1_8_16_r;
wire signed [`CalcTempBus]          temp_m1_8_16_i;
wire signed [`CalcTempBus]          temp_m1_8_17_r;
wire signed [`CalcTempBus]          temp_m1_8_17_i;
wire signed [`CalcTempBus]          temp_m1_8_18_r;
wire signed [`CalcTempBus]          temp_m1_8_18_i;
wire signed [`CalcTempBus]          temp_m1_8_19_r;
wire signed [`CalcTempBus]          temp_m1_8_19_i;
wire signed [`CalcTempBus]          temp_m1_8_20_r;
wire signed [`CalcTempBus]          temp_m1_8_20_i;
wire signed [`CalcTempBus]          temp_m1_8_21_r;
wire signed [`CalcTempBus]          temp_m1_8_21_i;
wire signed [`CalcTempBus]          temp_m1_8_22_r;
wire signed [`CalcTempBus]          temp_m1_8_22_i;
wire signed [`CalcTempBus]          temp_m1_8_23_r;
wire signed [`CalcTempBus]          temp_m1_8_23_i;
wire signed [`CalcTempBus]          temp_m1_8_24_r;
wire signed [`CalcTempBus]          temp_m1_8_24_i;
wire signed [`CalcTempBus]          temp_m1_8_25_r;
wire signed [`CalcTempBus]          temp_m1_8_25_i;
wire signed [`CalcTempBus]          temp_m1_8_26_r;
wire signed [`CalcTempBus]          temp_m1_8_26_i;
wire signed [`CalcTempBus]          temp_m1_8_27_r;
wire signed [`CalcTempBus]          temp_m1_8_27_i;
wire signed [`CalcTempBus]          temp_m1_8_28_r;
wire signed [`CalcTempBus]          temp_m1_8_28_i;
wire signed [`CalcTempBus]          temp_m1_8_29_r;
wire signed [`CalcTempBus]          temp_m1_8_29_i;
wire signed [`CalcTempBus]          temp_m1_8_30_r;
wire signed [`CalcTempBus]          temp_m1_8_30_i;
wire signed [`CalcTempBus]          temp_m1_8_31_r;
wire signed [`CalcTempBus]          temp_m1_8_31_i;
wire signed [`CalcTempBus]          temp_m1_8_32_r;
wire signed [`CalcTempBus]          temp_m1_8_32_i;
wire signed [`CalcTempBus]          temp_m1_9_1_r;
wire signed [`CalcTempBus]          temp_m1_9_1_i;
wire signed [`CalcTempBus]          temp_m1_9_2_r;
wire signed [`CalcTempBus]          temp_m1_9_2_i;
wire signed [`CalcTempBus]          temp_m1_9_3_r;
wire signed [`CalcTempBus]          temp_m1_9_3_i;
wire signed [`CalcTempBus]          temp_m1_9_4_r;
wire signed [`CalcTempBus]          temp_m1_9_4_i;
wire signed [`CalcTempBus]          temp_m1_9_5_r;
wire signed [`CalcTempBus]          temp_m1_9_5_i;
wire signed [`CalcTempBus]          temp_m1_9_6_r;
wire signed [`CalcTempBus]          temp_m1_9_6_i;
wire signed [`CalcTempBus]          temp_m1_9_7_r;
wire signed [`CalcTempBus]          temp_m1_9_7_i;
wire signed [`CalcTempBus]          temp_m1_9_8_r;
wire signed [`CalcTempBus]          temp_m1_9_8_i;
wire signed [`CalcTempBus]          temp_m1_9_9_r;
wire signed [`CalcTempBus]          temp_m1_9_9_i;
wire signed [`CalcTempBus]          temp_m1_9_10_r;
wire signed [`CalcTempBus]          temp_m1_9_10_i;
wire signed [`CalcTempBus]          temp_m1_9_11_r;
wire signed [`CalcTempBus]          temp_m1_9_11_i;
wire signed [`CalcTempBus]          temp_m1_9_12_r;
wire signed [`CalcTempBus]          temp_m1_9_12_i;
wire signed [`CalcTempBus]          temp_m1_9_13_r;
wire signed [`CalcTempBus]          temp_m1_9_13_i;
wire signed [`CalcTempBus]          temp_m1_9_14_r;
wire signed [`CalcTempBus]          temp_m1_9_14_i;
wire signed [`CalcTempBus]          temp_m1_9_15_r;
wire signed [`CalcTempBus]          temp_m1_9_15_i;
wire signed [`CalcTempBus]          temp_m1_9_16_r;
wire signed [`CalcTempBus]          temp_m1_9_16_i;
wire signed [`CalcTempBus]          temp_m1_9_17_r;
wire signed [`CalcTempBus]          temp_m1_9_17_i;
wire signed [`CalcTempBus]          temp_m1_9_18_r;
wire signed [`CalcTempBus]          temp_m1_9_18_i;
wire signed [`CalcTempBus]          temp_m1_9_19_r;
wire signed [`CalcTempBus]          temp_m1_9_19_i;
wire signed [`CalcTempBus]          temp_m1_9_20_r;
wire signed [`CalcTempBus]          temp_m1_9_20_i;
wire signed [`CalcTempBus]          temp_m1_9_21_r;
wire signed [`CalcTempBus]          temp_m1_9_21_i;
wire signed [`CalcTempBus]          temp_m1_9_22_r;
wire signed [`CalcTempBus]          temp_m1_9_22_i;
wire signed [`CalcTempBus]          temp_m1_9_23_r;
wire signed [`CalcTempBus]          temp_m1_9_23_i;
wire signed [`CalcTempBus]          temp_m1_9_24_r;
wire signed [`CalcTempBus]          temp_m1_9_24_i;
wire signed [`CalcTempBus]          temp_m1_9_25_r;
wire signed [`CalcTempBus]          temp_m1_9_25_i;
wire signed [`CalcTempBus]          temp_m1_9_26_r;
wire signed [`CalcTempBus]          temp_m1_9_26_i;
wire signed [`CalcTempBus]          temp_m1_9_27_r;
wire signed [`CalcTempBus]          temp_m1_9_27_i;
wire signed [`CalcTempBus]          temp_m1_9_28_r;
wire signed [`CalcTempBus]          temp_m1_9_28_i;
wire signed [`CalcTempBus]          temp_m1_9_29_r;
wire signed [`CalcTempBus]          temp_m1_9_29_i;
wire signed [`CalcTempBus]          temp_m1_9_30_r;
wire signed [`CalcTempBus]          temp_m1_9_30_i;
wire signed [`CalcTempBus]          temp_m1_9_31_r;
wire signed [`CalcTempBus]          temp_m1_9_31_i;
wire signed [`CalcTempBus]          temp_m1_9_32_r;
wire signed [`CalcTempBus]          temp_m1_9_32_i;
wire signed [`CalcTempBus]          temp_m1_10_1_r;
wire signed [`CalcTempBus]          temp_m1_10_1_i;
wire signed [`CalcTempBus]          temp_m1_10_2_r;
wire signed [`CalcTempBus]          temp_m1_10_2_i;
wire signed [`CalcTempBus]          temp_m1_10_3_r;
wire signed [`CalcTempBus]          temp_m1_10_3_i;
wire signed [`CalcTempBus]          temp_m1_10_4_r;
wire signed [`CalcTempBus]          temp_m1_10_4_i;
wire signed [`CalcTempBus]          temp_m1_10_5_r;
wire signed [`CalcTempBus]          temp_m1_10_5_i;
wire signed [`CalcTempBus]          temp_m1_10_6_r;
wire signed [`CalcTempBus]          temp_m1_10_6_i;
wire signed [`CalcTempBus]          temp_m1_10_7_r;
wire signed [`CalcTempBus]          temp_m1_10_7_i;
wire signed [`CalcTempBus]          temp_m1_10_8_r;
wire signed [`CalcTempBus]          temp_m1_10_8_i;
wire signed [`CalcTempBus]          temp_m1_10_9_r;
wire signed [`CalcTempBus]          temp_m1_10_9_i;
wire signed [`CalcTempBus]          temp_m1_10_10_r;
wire signed [`CalcTempBus]          temp_m1_10_10_i;
wire signed [`CalcTempBus]          temp_m1_10_11_r;
wire signed [`CalcTempBus]          temp_m1_10_11_i;
wire signed [`CalcTempBus]          temp_m1_10_12_r;
wire signed [`CalcTempBus]          temp_m1_10_12_i;
wire signed [`CalcTempBus]          temp_m1_10_13_r;
wire signed [`CalcTempBus]          temp_m1_10_13_i;
wire signed [`CalcTempBus]          temp_m1_10_14_r;
wire signed [`CalcTempBus]          temp_m1_10_14_i;
wire signed [`CalcTempBus]          temp_m1_10_15_r;
wire signed [`CalcTempBus]          temp_m1_10_15_i;
wire signed [`CalcTempBus]          temp_m1_10_16_r;
wire signed [`CalcTempBus]          temp_m1_10_16_i;
wire signed [`CalcTempBus]          temp_m1_10_17_r;
wire signed [`CalcTempBus]          temp_m1_10_17_i;
wire signed [`CalcTempBus]          temp_m1_10_18_r;
wire signed [`CalcTempBus]          temp_m1_10_18_i;
wire signed [`CalcTempBus]          temp_m1_10_19_r;
wire signed [`CalcTempBus]          temp_m1_10_19_i;
wire signed [`CalcTempBus]          temp_m1_10_20_r;
wire signed [`CalcTempBus]          temp_m1_10_20_i;
wire signed [`CalcTempBus]          temp_m1_10_21_r;
wire signed [`CalcTempBus]          temp_m1_10_21_i;
wire signed [`CalcTempBus]          temp_m1_10_22_r;
wire signed [`CalcTempBus]          temp_m1_10_22_i;
wire signed [`CalcTempBus]          temp_m1_10_23_r;
wire signed [`CalcTempBus]          temp_m1_10_23_i;
wire signed [`CalcTempBus]          temp_m1_10_24_r;
wire signed [`CalcTempBus]          temp_m1_10_24_i;
wire signed [`CalcTempBus]          temp_m1_10_25_r;
wire signed [`CalcTempBus]          temp_m1_10_25_i;
wire signed [`CalcTempBus]          temp_m1_10_26_r;
wire signed [`CalcTempBus]          temp_m1_10_26_i;
wire signed [`CalcTempBus]          temp_m1_10_27_r;
wire signed [`CalcTempBus]          temp_m1_10_27_i;
wire signed [`CalcTempBus]          temp_m1_10_28_r;
wire signed [`CalcTempBus]          temp_m1_10_28_i;
wire signed [`CalcTempBus]          temp_m1_10_29_r;
wire signed [`CalcTempBus]          temp_m1_10_29_i;
wire signed [`CalcTempBus]          temp_m1_10_30_r;
wire signed [`CalcTempBus]          temp_m1_10_30_i;
wire signed [`CalcTempBus]          temp_m1_10_31_r;
wire signed [`CalcTempBus]          temp_m1_10_31_i;
wire signed [`CalcTempBus]          temp_m1_10_32_r;
wire signed [`CalcTempBus]          temp_m1_10_32_i;
wire signed [`CalcTempBus]          temp_m1_11_1_r;
wire signed [`CalcTempBus]          temp_m1_11_1_i;
wire signed [`CalcTempBus]          temp_m1_11_2_r;
wire signed [`CalcTempBus]          temp_m1_11_2_i;
wire signed [`CalcTempBus]          temp_m1_11_3_r;
wire signed [`CalcTempBus]          temp_m1_11_3_i;
wire signed [`CalcTempBus]          temp_m1_11_4_r;
wire signed [`CalcTempBus]          temp_m1_11_4_i;
wire signed [`CalcTempBus]          temp_m1_11_5_r;
wire signed [`CalcTempBus]          temp_m1_11_5_i;
wire signed [`CalcTempBus]          temp_m1_11_6_r;
wire signed [`CalcTempBus]          temp_m1_11_6_i;
wire signed [`CalcTempBus]          temp_m1_11_7_r;
wire signed [`CalcTempBus]          temp_m1_11_7_i;
wire signed [`CalcTempBus]          temp_m1_11_8_r;
wire signed [`CalcTempBus]          temp_m1_11_8_i;
wire signed [`CalcTempBus]          temp_m1_11_9_r;
wire signed [`CalcTempBus]          temp_m1_11_9_i;
wire signed [`CalcTempBus]          temp_m1_11_10_r;
wire signed [`CalcTempBus]          temp_m1_11_10_i;
wire signed [`CalcTempBus]          temp_m1_11_11_r;
wire signed [`CalcTempBus]          temp_m1_11_11_i;
wire signed [`CalcTempBus]          temp_m1_11_12_r;
wire signed [`CalcTempBus]          temp_m1_11_12_i;
wire signed [`CalcTempBus]          temp_m1_11_13_r;
wire signed [`CalcTempBus]          temp_m1_11_13_i;
wire signed [`CalcTempBus]          temp_m1_11_14_r;
wire signed [`CalcTempBus]          temp_m1_11_14_i;
wire signed [`CalcTempBus]          temp_m1_11_15_r;
wire signed [`CalcTempBus]          temp_m1_11_15_i;
wire signed [`CalcTempBus]          temp_m1_11_16_r;
wire signed [`CalcTempBus]          temp_m1_11_16_i;
wire signed [`CalcTempBus]          temp_m1_11_17_r;
wire signed [`CalcTempBus]          temp_m1_11_17_i;
wire signed [`CalcTempBus]          temp_m1_11_18_r;
wire signed [`CalcTempBus]          temp_m1_11_18_i;
wire signed [`CalcTempBus]          temp_m1_11_19_r;
wire signed [`CalcTempBus]          temp_m1_11_19_i;
wire signed [`CalcTempBus]          temp_m1_11_20_r;
wire signed [`CalcTempBus]          temp_m1_11_20_i;
wire signed [`CalcTempBus]          temp_m1_11_21_r;
wire signed [`CalcTempBus]          temp_m1_11_21_i;
wire signed [`CalcTempBus]          temp_m1_11_22_r;
wire signed [`CalcTempBus]          temp_m1_11_22_i;
wire signed [`CalcTempBus]          temp_m1_11_23_r;
wire signed [`CalcTempBus]          temp_m1_11_23_i;
wire signed [`CalcTempBus]          temp_m1_11_24_r;
wire signed [`CalcTempBus]          temp_m1_11_24_i;
wire signed [`CalcTempBus]          temp_m1_11_25_r;
wire signed [`CalcTempBus]          temp_m1_11_25_i;
wire signed [`CalcTempBus]          temp_m1_11_26_r;
wire signed [`CalcTempBus]          temp_m1_11_26_i;
wire signed [`CalcTempBus]          temp_m1_11_27_r;
wire signed [`CalcTempBus]          temp_m1_11_27_i;
wire signed [`CalcTempBus]          temp_m1_11_28_r;
wire signed [`CalcTempBus]          temp_m1_11_28_i;
wire signed [`CalcTempBus]          temp_m1_11_29_r;
wire signed [`CalcTempBus]          temp_m1_11_29_i;
wire signed [`CalcTempBus]          temp_m1_11_30_r;
wire signed [`CalcTempBus]          temp_m1_11_30_i;
wire signed [`CalcTempBus]          temp_m1_11_31_r;
wire signed [`CalcTempBus]          temp_m1_11_31_i;
wire signed [`CalcTempBus]          temp_m1_11_32_r;
wire signed [`CalcTempBus]          temp_m1_11_32_i;
wire signed [`CalcTempBus]          temp_m1_12_1_r;
wire signed [`CalcTempBus]          temp_m1_12_1_i;
wire signed [`CalcTempBus]          temp_m1_12_2_r;
wire signed [`CalcTempBus]          temp_m1_12_2_i;
wire signed [`CalcTempBus]          temp_m1_12_3_r;
wire signed [`CalcTempBus]          temp_m1_12_3_i;
wire signed [`CalcTempBus]          temp_m1_12_4_r;
wire signed [`CalcTempBus]          temp_m1_12_4_i;
wire signed [`CalcTempBus]          temp_m1_12_5_r;
wire signed [`CalcTempBus]          temp_m1_12_5_i;
wire signed [`CalcTempBus]          temp_m1_12_6_r;
wire signed [`CalcTempBus]          temp_m1_12_6_i;
wire signed [`CalcTempBus]          temp_m1_12_7_r;
wire signed [`CalcTempBus]          temp_m1_12_7_i;
wire signed [`CalcTempBus]          temp_m1_12_8_r;
wire signed [`CalcTempBus]          temp_m1_12_8_i;
wire signed [`CalcTempBus]          temp_m1_12_9_r;
wire signed [`CalcTempBus]          temp_m1_12_9_i;
wire signed [`CalcTempBus]          temp_m1_12_10_r;
wire signed [`CalcTempBus]          temp_m1_12_10_i;
wire signed [`CalcTempBus]          temp_m1_12_11_r;
wire signed [`CalcTempBus]          temp_m1_12_11_i;
wire signed [`CalcTempBus]          temp_m1_12_12_r;
wire signed [`CalcTempBus]          temp_m1_12_12_i;
wire signed [`CalcTempBus]          temp_m1_12_13_r;
wire signed [`CalcTempBus]          temp_m1_12_13_i;
wire signed [`CalcTempBus]          temp_m1_12_14_r;
wire signed [`CalcTempBus]          temp_m1_12_14_i;
wire signed [`CalcTempBus]          temp_m1_12_15_r;
wire signed [`CalcTempBus]          temp_m1_12_15_i;
wire signed [`CalcTempBus]          temp_m1_12_16_r;
wire signed [`CalcTempBus]          temp_m1_12_16_i;
wire signed [`CalcTempBus]          temp_m1_12_17_r;
wire signed [`CalcTempBus]          temp_m1_12_17_i;
wire signed [`CalcTempBus]          temp_m1_12_18_r;
wire signed [`CalcTempBus]          temp_m1_12_18_i;
wire signed [`CalcTempBus]          temp_m1_12_19_r;
wire signed [`CalcTempBus]          temp_m1_12_19_i;
wire signed [`CalcTempBus]          temp_m1_12_20_r;
wire signed [`CalcTempBus]          temp_m1_12_20_i;
wire signed [`CalcTempBus]          temp_m1_12_21_r;
wire signed [`CalcTempBus]          temp_m1_12_21_i;
wire signed [`CalcTempBus]          temp_m1_12_22_r;
wire signed [`CalcTempBus]          temp_m1_12_22_i;
wire signed [`CalcTempBus]          temp_m1_12_23_r;
wire signed [`CalcTempBus]          temp_m1_12_23_i;
wire signed [`CalcTempBus]          temp_m1_12_24_r;
wire signed [`CalcTempBus]          temp_m1_12_24_i;
wire signed [`CalcTempBus]          temp_m1_12_25_r;
wire signed [`CalcTempBus]          temp_m1_12_25_i;
wire signed [`CalcTempBus]          temp_m1_12_26_r;
wire signed [`CalcTempBus]          temp_m1_12_26_i;
wire signed [`CalcTempBus]          temp_m1_12_27_r;
wire signed [`CalcTempBus]          temp_m1_12_27_i;
wire signed [`CalcTempBus]          temp_m1_12_28_r;
wire signed [`CalcTempBus]          temp_m1_12_28_i;
wire signed [`CalcTempBus]          temp_m1_12_29_r;
wire signed [`CalcTempBus]          temp_m1_12_29_i;
wire signed [`CalcTempBus]          temp_m1_12_30_r;
wire signed [`CalcTempBus]          temp_m1_12_30_i;
wire signed [`CalcTempBus]          temp_m1_12_31_r;
wire signed [`CalcTempBus]          temp_m1_12_31_i;
wire signed [`CalcTempBus]          temp_m1_12_32_r;
wire signed [`CalcTempBus]          temp_m1_12_32_i;
wire signed [`CalcTempBus]          temp_m1_13_1_r;
wire signed [`CalcTempBus]          temp_m1_13_1_i;
wire signed [`CalcTempBus]          temp_m1_13_2_r;
wire signed [`CalcTempBus]          temp_m1_13_2_i;
wire signed [`CalcTempBus]          temp_m1_13_3_r;
wire signed [`CalcTempBus]          temp_m1_13_3_i;
wire signed [`CalcTempBus]          temp_m1_13_4_r;
wire signed [`CalcTempBus]          temp_m1_13_4_i;
wire signed [`CalcTempBus]          temp_m1_13_5_r;
wire signed [`CalcTempBus]          temp_m1_13_5_i;
wire signed [`CalcTempBus]          temp_m1_13_6_r;
wire signed [`CalcTempBus]          temp_m1_13_6_i;
wire signed [`CalcTempBus]          temp_m1_13_7_r;
wire signed [`CalcTempBus]          temp_m1_13_7_i;
wire signed [`CalcTempBus]          temp_m1_13_8_r;
wire signed [`CalcTempBus]          temp_m1_13_8_i;
wire signed [`CalcTempBus]          temp_m1_13_9_r;
wire signed [`CalcTempBus]          temp_m1_13_9_i;
wire signed [`CalcTempBus]          temp_m1_13_10_r;
wire signed [`CalcTempBus]          temp_m1_13_10_i;
wire signed [`CalcTempBus]          temp_m1_13_11_r;
wire signed [`CalcTempBus]          temp_m1_13_11_i;
wire signed [`CalcTempBus]          temp_m1_13_12_r;
wire signed [`CalcTempBus]          temp_m1_13_12_i;
wire signed [`CalcTempBus]          temp_m1_13_13_r;
wire signed [`CalcTempBus]          temp_m1_13_13_i;
wire signed [`CalcTempBus]          temp_m1_13_14_r;
wire signed [`CalcTempBus]          temp_m1_13_14_i;
wire signed [`CalcTempBus]          temp_m1_13_15_r;
wire signed [`CalcTempBus]          temp_m1_13_15_i;
wire signed [`CalcTempBus]          temp_m1_13_16_r;
wire signed [`CalcTempBus]          temp_m1_13_16_i;
wire signed [`CalcTempBus]          temp_m1_13_17_r;
wire signed [`CalcTempBus]          temp_m1_13_17_i;
wire signed [`CalcTempBus]          temp_m1_13_18_r;
wire signed [`CalcTempBus]          temp_m1_13_18_i;
wire signed [`CalcTempBus]          temp_m1_13_19_r;
wire signed [`CalcTempBus]          temp_m1_13_19_i;
wire signed [`CalcTempBus]          temp_m1_13_20_r;
wire signed [`CalcTempBus]          temp_m1_13_20_i;
wire signed [`CalcTempBus]          temp_m1_13_21_r;
wire signed [`CalcTempBus]          temp_m1_13_21_i;
wire signed [`CalcTempBus]          temp_m1_13_22_r;
wire signed [`CalcTempBus]          temp_m1_13_22_i;
wire signed [`CalcTempBus]          temp_m1_13_23_r;
wire signed [`CalcTempBus]          temp_m1_13_23_i;
wire signed [`CalcTempBus]          temp_m1_13_24_r;
wire signed [`CalcTempBus]          temp_m1_13_24_i;
wire signed [`CalcTempBus]          temp_m1_13_25_r;
wire signed [`CalcTempBus]          temp_m1_13_25_i;
wire signed [`CalcTempBus]          temp_m1_13_26_r;
wire signed [`CalcTempBus]          temp_m1_13_26_i;
wire signed [`CalcTempBus]          temp_m1_13_27_r;
wire signed [`CalcTempBus]          temp_m1_13_27_i;
wire signed [`CalcTempBus]          temp_m1_13_28_r;
wire signed [`CalcTempBus]          temp_m1_13_28_i;
wire signed [`CalcTempBus]          temp_m1_13_29_r;
wire signed [`CalcTempBus]          temp_m1_13_29_i;
wire signed [`CalcTempBus]          temp_m1_13_30_r;
wire signed [`CalcTempBus]          temp_m1_13_30_i;
wire signed [`CalcTempBus]          temp_m1_13_31_r;
wire signed [`CalcTempBus]          temp_m1_13_31_i;
wire signed [`CalcTempBus]          temp_m1_13_32_r;
wire signed [`CalcTempBus]          temp_m1_13_32_i;
wire signed [`CalcTempBus]          temp_m1_14_1_r;
wire signed [`CalcTempBus]          temp_m1_14_1_i;
wire signed [`CalcTempBus]          temp_m1_14_2_r;
wire signed [`CalcTempBus]          temp_m1_14_2_i;
wire signed [`CalcTempBus]          temp_m1_14_3_r;
wire signed [`CalcTempBus]          temp_m1_14_3_i;
wire signed [`CalcTempBus]          temp_m1_14_4_r;
wire signed [`CalcTempBus]          temp_m1_14_4_i;
wire signed [`CalcTempBus]          temp_m1_14_5_r;
wire signed [`CalcTempBus]          temp_m1_14_5_i;
wire signed [`CalcTempBus]          temp_m1_14_6_r;
wire signed [`CalcTempBus]          temp_m1_14_6_i;
wire signed [`CalcTempBus]          temp_m1_14_7_r;
wire signed [`CalcTempBus]          temp_m1_14_7_i;
wire signed [`CalcTempBus]          temp_m1_14_8_r;
wire signed [`CalcTempBus]          temp_m1_14_8_i;
wire signed [`CalcTempBus]          temp_m1_14_9_r;
wire signed [`CalcTempBus]          temp_m1_14_9_i;
wire signed [`CalcTempBus]          temp_m1_14_10_r;
wire signed [`CalcTempBus]          temp_m1_14_10_i;
wire signed [`CalcTempBus]          temp_m1_14_11_r;
wire signed [`CalcTempBus]          temp_m1_14_11_i;
wire signed [`CalcTempBus]          temp_m1_14_12_r;
wire signed [`CalcTempBus]          temp_m1_14_12_i;
wire signed [`CalcTempBus]          temp_m1_14_13_r;
wire signed [`CalcTempBus]          temp_m1_14_13_i;
wire signed [`CalcTempBus]          temp_m1_14_14_r;
wire signed [`CalcTempBus]          temp_m1_14_14_i;
wire signed [`CalcTempBus]          temp_m1_14_15_r;
wire signed [`CalcTempBus]          temp_m1_14_15_i;
wire signed [`CalcTempBus]          temp_m1_14_16_r;
wire signed [`CalcTempBus]          temp_m1_14_16_i;
wire signed [`CalcTempBus]          temp_m1_14_17_r;
wire signed [`CalcTempBus]          temp_m1_14_17_i;
wire signed [`CalcTempBus]          temp_m1_14_18_r;
wire signed [`CalcTempBus]          temp_m1_14_18_i;
wire signed [`CalcTempBus]          temp_m1_14_19_r;
wire signed [`CalcTempBus]          temp_m1_14_19_i;
wire signed [`CalcTempBus]          temp_m1_14_20_r;
wire signed [`CalcTempBus]          temp_m1_14_20_i;
wire signed [`CalcTempBus]          temp_m1_14_21_r;
wire signed [`CalcTempBus]          temp_m1_14_21_i;
wire signed [`CalcTempBus]          temp_m1_14_22_r;
wire signed [`CalcTempBus]          temp_m1_14_22_i;
wire signed [`CalcTempBus]          temp_m1_14_23_r;
wire signed [`CalcTempBus]          temp_m1_14_23_i;
wire signed [`CalcTempBus]          temp_m1_14_24_r;
wire signed [`CalcTempBus]          temp_m1_14_24_i;
wire signed [`CalcTempBus]          temp_m1_14_25_r;
wire signed [`CalcTempBus]          temp_m1_14_25_i;
wire signed [`CalcTempBus]          temp_m1_14_26_r;
wire signed [`CalcTempBus]          temp_m1_14_26_i;
wire signed [`CalcTempBus]          temp_m1_14_27_r;
wire signed [`CalcTempBus]          temp_m1_14_27_i;
wire signed [`CalcTempBus]          temp_m1_14_28_r;
wire signed [`CalcTempBus]          temp_m1_14_28_i;
wire signed [`CalcTempBus]          temp_m1_14_29_r;
wire signed [`CalcTempBus]          temp_m1_14_29_i;
wire signed [`CalcTempBus]          temp_m1_14_30_r;
wire signed [`CalcTempBus]          temp_m1_14_30_i;
wire signed [`CalcTempBus]          temp_m1_14_31_r;
wire signed [`CalcTempBus]          temp_m1_14_31_i;
wire signed [`CalcTempBus]          temp_m1_14_32_r;
wire signed [`CalcTempBus]          temp_m1_14_32_i;
wire signed [`CalcTempBus]          temp_m1_15_1_r;
wire signed [`CalcTempBus]          temp_m1_15_1_i;
wire signed [`CalcTempBus]          temp_m1_15_2_r;
wire signed [`CalcTempBus]          temp_m1_15_2_i;
wire signed [`CalcTempBus]          temp_m1_15_3_r;
wire signed [`CalcTempBus]          temp_m1_15_3_i;
wire signed [`CalcTempBus]          temp_m1_15_4_r;
wire signed [`CalcTempBus]          temp_m1_15_4_i;
wire signed [`CalcTempBus]          temp_m1_15_5_r;
wire signed [`CalcTempBus]          temp_m1_15_5_i;
wire signed [`CalcTempBus]          temp_m1_15_6_r;
wire signed [`CalcTempBus]          temp_m1_15_6_i;
wire signed [`CalcTempBus]          temp_m1_15_7_r;
wire signed [`CalcTempBus]          temp_m1_15_7_i;
wire signed [`CalcTempBus]          temp_m1_15_8_r;
wire signed [`CalcTempBus]          temp_m1_15_8_i;
wire signed [`CalcTempBus]          temp_m1_15_9_r;
wire signed [`CalcTempBus]          temp_m1_15_9_i;
wire signed [`CalcTempBus]          temp_m1_15_10_r;
wire signed [`CalcTempBus]          temp_m1_15_10_i;
wire signed [`CalcTempBus]          temp_m1_15_11_r;
wire signed [`CalcTempBus]          temp_m1_15_11_i;
wire signed [`CalcTempBus]          temp_m1_15_12_r;
wire signed [`CalcTempBus]          temp_m1_15_12_i;
wire signed [`CalcTempBus]          temp_m1_15_13_r;
wire signed [`CalcTempBus]          temp_m1_15_13_i;
wire signed [`CalcTempBus]          temp_m1_15_14_r;
wire signed [`CalcTempBus]          temp_m1_15_14_i;
wire signed [`CalcTempBus]          temp_m1_15_15_r;
wire signed [`CalcTempBus]          temp_m1_15_15_i;
wire signed [`CalcTempBus]          temp_m1_15_16_r;
wire signed [`CalcTempBus]          temp_m1_15_16_i;
wire signed [`CalcTempBus]          temp_m1_15_17_r;
wire signed [`CalcTempBus]          temp_m1_15_17_i;
wire signed [`CalcTempBus]          temp_m1_15_18_r;
wire signed [`CalcTempBus]          temp_m1_15_18_i;
wire signed [`CalcTempBus]          temp_m1_15_19_r;
wire signed [`CalcTempBus]          temp_m1_15_19_i;
wire signed [`CalcTempBus]          temp_m1_15_20_r;
wire signed [`CalcTempBus]          temp_m1_15_20_i;
wire signed [`CalcTempBus]          temp_m1_15_21_r;
wire signed [`CalcTempBus]          temp_m1_15_21_i;
wire signed [`CalcTempBus]          temp_m1_15_22_r;
wire signed [`CalcTempBus]          temp_m1_15_22_i;
wire signed [`CalcTempBus]          temp_m1_15_23_r;
wire signed [`CalcTempBus]          temp_m1_15_23_i;
wire signed [`CalcTempBus]          temp_m1_15_24_r;
wire signed [`CalcTempBus]          temp_m1_15_24_i;
wire signed [`CalcTempBus]          temp_m1_15_25_r;
wire signed [`CalcTempBus]          temp_m1_15_25_i;
wire signed [`CalcTempBus]          temp_m1_15_26_r;
wire signed [`CalcTempBus]          temp_m1_15_26_i;
wire signed [`CalcTempBus]          temp_m1_15_27_r;
wire signed [`CalcTempBus]          temp_m1_15_27_i;
wire signed [`CalcTempBus]          temp_m1_15_28_r;
wire signed [`CalcTempBus]          temp_m1_15_28_i;
wire signed [`CalcTempBus]          temp_m1_15_29_r;
wire signed [`CalcTempBus]          temp_m1_15_29_i;
wire signed [`CalcTempBus]          temp_m1_15_30_r;
wire signed [`CalcTempBus]          temp_m1_15_30_i;
wire signed [`CalcTempBus]          temp_m1_15_31_r;
wire signed [`CalcTempBus]          temp_m1_15_31_i;
wire signed [`CalcTempBus]          temp_m1_15_32_r;
wire signed [`CalcTempBus]          temp_m1_15_32_i;
wire signed [`CalcTempBus]          temp_m1_16_1_r;
wire signed [`CalcTempBus]          temp_m1_16_1_i;
wire signed [`CalcTempBus]          temp_m1_16_2_r;
wire signed [`CalcTempBus]          temp_m1_16_2_i;
wire signed [`CalcTempBus]          temp_m1_16_3_r;
wire signed [`CalcTempBus]          temp_m1_16_3_i;
wire signed [`CalcTempBus]          temp_m1_16_4_r;
wire signed [`CalcTempBus]          temp_m1_16_4_i;
wire signed [`CalcTempBus]          temp_m1_16_5_r;
wire signed [`CalcTempBus]          temp_m1_16_5_i;
wire signed [`CalcTempBus]          temp_m1_16_6_r;
wire signed [`CalcTempBus]          temp_m1_16_6_i;
wire signed [`CalcTempBus]          temp_m1_16_7_r;
wire signed [`CalcTempBus]          temp_m1_16_7_i;
wire signed [`CalcTempBus]          temp_m1_16_8_r;
wire signed [`CalcTempBus]          temp_m1_16_8_i;
wire signed [`CalcTempBus]          temp_m1_16_9_r;
wire signed [`CalcTempBus]          temp_m1_16_9_i;
wire signed [`CalcTempBus]          temp_m1_16_10_r;
wire signed [`CalcTempBus]          temp_m1_16_10_i;
wire signed [`CalcTempBus]          temp_m1_16_11_r;
wire signed [`CalcTempBus]          temp_m1_16_11_i;
wire signed [`CalcTempBus]          temp_m1_16_12_r;
wire signed [`CalcTempBus]          temp_m1_16_12_i;
wire signed [`CalcTempBus]          temp_m1_16_13_r;
wire signed [`CalcTempBus]          temp_m1_16_13_i;
wire signed [`CalcTempBus]          temp_m1_16_14_r;
wire signed [`CalcTempBus]          temp_m1_16_14_i;
wire signed [`CalcTempBus]          temp_m1_16_15_r;
wire signed [`CalcTempBus]          temp_m1_16_15_i;
wire signed [`CalcTempBus]          temp_m1_16_16_r;
wire signed [`CalcTempBus]          temp_m1_16_16_i;
wire signed [`CalcTempBus]          temp_m1_16_17_r;
wire signed [`CalcTempBus]          temp_m1_16_17_i;
wire signed [`CalcTempBus]          temp_m1_16_18_r;
wire signed [`CalcTempBus]          temp_m1_16_18_i;
wire signed [`CalcTempBus]          temp_m1_16_19_r;
wire signed [`CalcTempBus]          temp_m1_16_19_i;
wire signed [`CalcTempBus]          temp_m1_16_20_r;
wire signed [`CalcTempBus]          temp_m1_16_20_i;
wire signed [`CalcTempBus]          temp_m1_16_21_r;
wire signed [`CalcTempBus]          temp_m1_16_21_i;
wire signed [`CalcTempBus]          temp_m1_16_22_r;
wire signed [`CalcTempBus]          temp_m1_16_22_i;
wire signed [`CalcTempBus]          temp_m1_16_23_r;
wire signed [`CalcTempBus]          temp_m1_16_23_i;
wire signed [`CalcTempBus]          temp_m1_16_24_r;
wire signed [`CalcTempBus]          temp_m1_16_24_i;
wire signed [`CalcTempBus]          temp_m1_16_25_r;
wire signed [`CalcTempBus]          temp_m1_16_25_i;
wire signed [`CalcTempBus]          temp_m1_16_26_r;
wire signed [`CalcTempBus]          temp_m1_16_26_i;
wire signed [`CalcTempBus]          temp_m1_16_27_r;
wire signed [`CalcTempBus]          temp_m1_16_27_i;
wire signed [`CalcTempBus]          temp_m1_16_28_r;
wire signed [`CalcTempBus]          temp_m1_16_28_i;
wire signed [`CalcTempBus]          temp_m1_16_29_r;
wire signed [`CalcTempBus]          temp_m1_16_29_i;
wire signed [`CalcTempBus]          temp_m1_16_30_r;
wire signed [`CalcTempBus]          temp_m1_16_30_i;
wire signed [`CalcTempBus]          temp_m1_16_31_r;
wire signed [`CalcTempBus]          temp_m1_16_31_i;
wire signed [`CalcTempBus]          temp_m1_16_32_r;
wire signed [`CalcTempBus]          temp_m1_16_32_i;
wire signed [`CalcTempBus]          temp_m1_17_1_r;
wire signed [`CalcTempBus]          temp_m1_17_1_i;
wire signed [`CalcTempBus]          temp_m1_17_2_r;
wire signed [`CalcTempBus]          temp_m1_17_2_i;
wire signed [`CalcTempBus]          temp_m1_17_3_r;
wire signed [`CalcTempBus]          temp_m1_17_3_i;
wire signed [`CalcTempBus]          temp_m1_17_4_r;
wire signed [`CalcTempBus]          temp_m1_17_4_i;
wire signed [`CalcTempBus]          temp_m1_17_5_r;
wire signed [`CalcTempBus]          temp_m1_17_5_i;
wire signed [`CalcTempBus]          temp_m1_17_6_r;
wire signed [`CalcTempBus]          temp_m1_17_6_i;
wire signed [`CalcTempBus]          temp_m1_17_7_r;
wire signed [`CalcTempBus]          temp_m1_17_7_i;
wire signed [`CalcTempBus]          temp_m1_17_8_r;
wire signed [`CalcTempBus]          temp_m1_17_8_i;
wire signed [`CalcTempBus]          temp_m1_17_9_r;
wire signed [`CalcTempBus]          temp_m1_17_9_i;
wire signed [`CalcTempBus]          temp_m1_17_10_r;
wire signed [`CalcTempBus]          temp_m1_17_10_i;
wire signed [`CalcTempBus]          temp_m1_17_11_r;
wire signed [`CalcTempBus]          temp_m1_17_11_i;
wire signed [`CalcTempBus]          temp_m1_17_12_r;
wire signed [`CalcTempBus]          temp_m1_17_12_i;
wire signed [`CalcTempBus]          temp_m1_17_13_r;
wire signed [`CalcTempBus]          temp_m1_17_13_i;
wire signed [`CalcTempBus]          temp_m1_17_14_r;
wire signed [`CalcTempBus]          temp_m1_17_14_i;
wire signed [`CalcTempBus]          temp_m1_17_15_r;
wire signed [`CalcTempBus]          temp_m1_17_15_i;
wire signed [`CalcTempBus]          temp_m1_17_16_r;
wire signed [`CalcTempBus]          temp_m1_17_16_i;
wire signed [`CalcTempBus]          temp_m1_17_17_r;
wire signed [`CalcTempBus]          temp_m1_17_17_i;
wire signed [`CalcTempBus]          temp_m1_17_18_r;
wire signed [`CalcTempBus]          temp_m1_17_18_i;
wire signed [`CalcTempBus]          temp_m1_17_19_r;
wire signed [`CalcTempBus]          temp_m1_17_19_i;
wire signed [`CalcTempBus]          temp_m1_17_20_r;
wire signed [`CalcTempBus]          temp_m1_17_20_i;
wire signed [`CalcTempBus]          temp_m1_17_21_r;
wire signed [`CalcTempBus]          temp_m1_17_21_i;
wire signed [`CalcTempBus]          temp_m1_17_22_r;
wire signed [`CalcTempBus]          temp_m1_17_22_i;
wire signed [`CalcTempBus]          temp_m1_17_23_r;
wire signed [`CalcTempBus]          temp_m1_17_23_i;
wire signed [`CalcTempBus]          temp_m1_17_24_r;
wire signed [`CalcTempBus]          temp_m1_17_24_i;
wire signed [`CalcTempBus]          temp_m1_17_25_r;
wire signed [`CalcTempBus]          temp_m1_17_25_i;
wire signed [`CalcTempBus]          temp_m1_17_26_r;
wire signed [`CalcTempBus]          temp_m1_17_26_i;
wire signed [`CalcTempBus]          temp_m1_17_27_r;
wire signed [`CalcTempBus]          temp_m1_17_27_i;
wire signed [`CalcTempBus]          temp_m1_17_28_r;
wire signed [`CalcTempBus]          temp_m1_17_28_i;
wire signed [`CalcTempBus]          temp_m1_17_29_r;
wire signed [`CalcTempBus]          temp_m1_17_29_i;
wire signed [`CalcTempBus]          temp_m1_17_30_r;
wire signed [`CalcTempBus]          temp_m1_17_30_i;
wire signed [`CalcTempBus]          temp_m1_17_31_r;
wire signed [`CalcTempBus]          temp_m1_17_31_i;
wire signed [`CalcTempBus]          temp_m1_17_32_r;
wire signed [`CalcTempBus]          temp_m1_17_32_i;
wire signed [`CalcTempBus]          temp_m1_18_1_r;
wire signed [`CalcTempBus]          temp_m1_18_1_i;
wire signed [`CalcTempBus]          temp_m1_18_2_r;
wire signed [`CalcTempBus]          temp_m1_18_2_i;
wire signed [`CalcTempBus]          temp_m1_18_3_r;
wire signed [`CalcTempBus]          temp_m1_18_3_i;
wire signed [`CalcTempBus]          temp_m1_18_4_r;
wire signed [`CalcTempBus]          temp_m1_18_4_i;
wire signed [`CalcTempBus]          temp_m1_18_5_r;
wire signed [`CalcTempBus]          temp_m1_18_5_i;
wire signed [`CalcTempBus]          temp_m1_18_6_r;
wire signed [`CalcTempBus]          temp_m1_18_6_i;
wire signed [`CalcTempBus]          temp_m1_18_7_r;
wire signed [`CalcTempBus]          temp_m1_18_7_i;
wire signed [`CalcTempBus]          temp_m1_18_8_r;
wire signed [`CalcTempBus]          temp_m1_18_8_i;
wire signed [`CalcTempBus]          temp_m1_18_9_r;
wire signed [`CalcTempBus]          temp_m1_18_9_i;
wire signed [`CalcTempBus]          temp_m1_18_10_r;
wire signed [`CalcTempBus]          temp_m1_18_10_i;
wire signed [`CalcTempBus]          temp_m1_18_11_r;
wire signed [`CalcTempBus]          temp_m1_18_11_i;
wire signed [`CalcTempBus]          temp_m1_18_12_r;
wire signed [`CalcTempBus]          temp_m1_18_12_i;
wire signed [`CalcTempBus]          temp_m1_18_13_r;
wire signed [`CalcTempBus]          temp_m1_18_13_i;
wire signed [`CalcTempBus]          temp_m1_18_14_r;
wire signed [`CalcTempBus]          temp_m1_18_14_i;
wire signed [`CalcTempBus]          temp_m1_18_15_r;
wire signed [`CalcTempBus]          temp_m1_18_15_i;
wire signed [`CalcTempBus]          temp_m1_18_16_r;
wire signed [`CalcTempBus]          temp_m1_18_16_i;
wire signed [`CalcTempBus]          temp_m1_18_17_r;
wire signed [`CalcTempBus]          temp_m1_18_17_i;
wire signed [`CalcTempBus]          temp_m1_18_18_r;
wire signed [`CalcTempBus]          temp_m1_18_18_i;
wire signed [`CalcTempBus]          temp_m1_18_19_r;
wire signed [`CalcTempBus]          temp_m1_18_19_i;
wire signed [`CalcTempBus]          temp_m1_18_20_r;
wire signed [`CalcTempBus]          temp_m1_18_20_i;
wire signed [`CalcTempBus]          temp_m1_18_21_r;
wire signed [`CalcTempBus]          temp_m1_18_21_i;
wire signed [`CalcTempBus]          temp_m1_18_22_r;
wire signed [`CalcTempBus]          temp_m1_18_22_i;
wire signed [`CalcTempBus]          temp_m1_18_23_r;
wire signed [`CalcTempBus]          temp_m1_18_23_i;
wire signed [`CalcTempBus]          temp_m1_18_24_r;
wire signed [`CalcTempBus]          temp_m1_18_24_i;
wire signed [`CalcTempBus]          temp_m1_18_25_r;
wire signed [`CalcTempBus]          temp_m1_18_25_i;
wire signed [`CalcTempBus]          temp_m1_18_26_r;
wire signed [`CalcTempBus]          temp_m1_18_26_i;
wire signed [`CalcTempBus]          temp_m1_18_27_r;
wire signed [`CalcTempBus]          temp_m1_18_27_i;
wire signed [`CalcTempBus]          temp_m1_18_28_r;
wire signed [`CalcTempBus]          temp_m1_18_28_i;
wire signed [`CalcTempBus]          temp_m1_18_29_r;
wire signed [`CalcTempBus]          temp_m1_18_29_i;
wire signed [`CalcTempBus]          temp_m1_18_30_r;
wire signed [`CalcTempBus]          temp_m1_18_30_i;
wire signed [`CalcTempBus]          temp_m1_18_31_r;
wire signed [`CalcTempBus]          temp_m1_18_31_i;
wire signed [`CalcTempBus]          temp_m1_18_32_r;
wire signed [`CalcTempBus]          temp_m1_18_32_i;
wire signed [`CalcTempBus]          temp_m1_19_1_r;
wire signed [`CalcTempBus]          temp_m1_19_1_i;
wire signed [`CalcTempBus]          temp_m1_19_2_r;
wire signed [`CalcTempBus]          temp_m1_19_2_i;
wire signed [`CalcTempBus]          temp_m1_19_3_r;
wire signed [`CalcTempBus]          temp_m1_19_3_i;
wire signed [`CalcTempBus]          temp_m1_19_4_r;
wire signed [`CalcTempBus]          temp_m1_19_4_i;
wire signed [`CalcTempBus]          temp_m1_19_5_r;
wire signed [`CalcTempBus]          temp_m1_19_5_i;
wire signed [`CalcTempBus]          temp_m1_19_6_r;
wire signed [`CalcTempBus]          temp_m1_19_6_i;
wire signed [`CalcTempBus]          temp_m1_19_7_r;
wire signed [`CalcTempBus]          temp_m1_19_7_i;
wire signed [`CalcTempBus]          temp_m1_19_8_r;
wire signed [`CalcTempBus]          temp_m1_19_8_i;
wire signed [`CalcTempBus]          temp_m1_19_9_r;
wire signed [`CalcTempBus]          temp_m1_19_9_i;
wire signed [`CalcTempBus]          temp_m1_19_10_r;
wire signed [`CalcTempBus]          temp_m1_19_10_i;
wire signed [`CalcTempBus]          temp_m1_19_11_r;
wire signed [`CalcTempBus]          temp_m1_19_11_i;
wire signed [`CalcTempBus]          temp_m1_19_12_r;
wire signed [`CalcTempBus]          temp_m1_19_12_i;
wire signed [`CalcTempBus]          temp_m1_19_13_r;
wire signed [`CalcTempBus]          temp_m1_19_13_i;
wire signed [`CalcTempBus]          temp_m1_19_14_r;
wire signed [`CalcTempBus]          temp_m1_19_14_i;
wire signed [`CalcTempBus]          temp_m1_19_15_r;
wire signed [`CalcTempBus]          temp_m1_19_15_i;
wire signed [`CalcTempBus]          temp_m1_19_16_r;
wire signed [`CalcTempBus]          temp_m1_19_16_i;
wire signed [`CalcTempBus]          temp_m1_19_17_r;
wire signed [`CalcTempBus]          temp_m1_19_17_i;
wire signed [`CalcTempBus]          temp_m1_19_18_r;
wire signed [`CalcTempBus]          temp_m1_19_18_i;
wire signed [`CalcTempBus]          temp_m1_19_19_r;
wire signed [`CalcTempBus]          temp_m1_19_19_i;
wire signed [`CalcTempBus]          temp_m1_19_20_r;
wire signed [`CalcTempBus]          temp_m1_19_20_i;
wire signed [`CalcTempBus]          temp_m1_19_21_r;
wire signed [`CalcTempBus]          temp_m1_19_21_i;
wire signed [`CalcTempBus]          temp_m1_19_22_r;
wire signed [`CalcTempBus]          temp_m1_19_22_i;
wire signed [`CalcTempBus]          temp_m1_19_23_r;
wire signed [`CalcTempBus]          temp_m1_19_23_i;
wire signed [`CalcTempBus]          temp_m1_19_24_r;
wire signed [`CalcTempBus]          temp_m1_19_24_i;
wire signed [`CalcTempBus]          temp_m1_19_25_r;
wire signed [`CalcTempBus]          temp_m1_19_25_i;
wire signed [`CalcTempBus]          temp_m1_19_26_r;
wire signed [`CalcTempBus]          temp_m1_19_26_i;
wire signed [`CalcTempBus]          temp_m1_19_27_r;
wire signed [`CalcTempBus]          temp_m1_19_27_i;
wire signed [`CalcTempBus]          temp_m1_19_28_r;
wire signed [`CalcTempBus]          temp_m1_19_28_i;
wire signed [`CalcTempBus]          temp_m1_19_29_r;
wire signed [`CalcTempBus]          temp_m1_19_29_i;
wire signed [`CalcTempBus]          temp_m1_19_30_r;
wire signed [`CalcTempBus]          temp_m1_19_30_i;
wire signed [`CalcTempBus]          temp_m1_19_31_r;
wire signed [`CalcTempBus]          temp_m1_19_31_i;
wire signed [`CalcTempBus]          temp_m1_19_32_r;
wire signed [`CalcTempBus]          temp_m1_19_32_i;
wire signed [`CalcTempBus]          temp_m1_20_1_r;
wire signed [`CalcTempBus]          temp_m1_20_1_i;
wire signed [`CalcTempBus]          temp_m1_20_2_r;
wire signed [`CalcTempBus]          temp_m1_20_2_i;
wire signed [`CalcTempBus]          temp_m1_20_3_r;
wire signed [`CalcTempBus]          temp_m1_20_3_i;
wire signed [`CalcTempBus]          temp_m1_20_4_r;
wire signed [`CalcTempBus]          temp_m1_20_4_i;
wire signed [`CalcTempBus]          temp_m1_20_5_r;
wire signed [`CalcTempBus]          temp_m1_20_5_i;
wire signed [`CalcTempBus]          temp_m1_20_6_r;
wire signed [`CalcTempBus]          temp_m1_20_6_i;
wire signed [`CalcTempBus]          temp_m1_20_7_r;
wire signed [`CalcTempBus]          temp_m1_20_7_i;
wire signed [`CalcTempBus]          temp_m1_20_8_r;
wire signed [`CalcTempBus]          temp_m1_20_8_i;
wire signed [`CalcTempBus]          temp_m1_20_9_r;
wire signed [`CalcTempBus]          temp_m1_20_9_i;
wire signed [`CalcTempBus]          temp_m1_20_10_r;
wire signed [`CalcTempBus]          temp_m1_20_10_i;
wire signed [`CalcTempBus]          temp_m1_20_11_r;
wire signed [`CalcTempBus]          temp_m1_20_11_i;
wire signed [`CalcTempBus]          temp_m1_20_12_r;
wire signed [`CalcTempBus]          temp_m1_20_12_i;
wire signed [`CalcTempBus]          temp_m1_20_13_r;
wire signed [`CalcTempBus]          temp_m1_20_13_i;
wire signed [`CalcTempBus]          temp_m1_20_14_r;
wire signed [`CalcTempBus]          temp_m1_20_14_i;
wire signed [`CalcTempBus]          temp_m1_20_15_r;
wire signed [`CalcTempBus]          temp_m1_20_15_i;
wire signed [`CalcTempBus]          temp_m1_20_16_r;
wire signed [`CalcTempBus]          temp_m1_20_16_i;
wire signed [`CalcTempBus]          temp_m1_20_17_r;
wire signed [`CalcTempBus]          temp_m1_20_17_i;
wire signed [`CalcTempBus]          temp_m1_20_18_r;
wire signed [`CalcTempBus]          temp_m1_20_18_i;
wire signed [`CalcTempBus]          temp_m1_20_19_r;
wire signed [`CalcTempBus]          temp_m1_20_19_i;
wire signed [`CalcTempBus]          temp_m1_20_20_r;
wire signed [`CalcTempBus]          temp_m1_20_20_i;
wire signed [`CalcTempBus]          temp_m1_20_21_r;
wire signed [`CalcTempBus]          temp_m1_20_21_i;
wire signed [`CalcTempBus]          temp_m1_20_22_r;
wire signed [`CalcTempBus]          temp_m1_20_22_i;
wire signed [`CalcTempBus]          temp_m1_20_23_r;
wire signed [`CalcTempBus]          temp_m1_20_23_i;
wire signed [`CalcTempBus]          temp_m1_20_24_r;
wire signed [`CalcTempBus]          temp_m1_20_24_i;
wire signed [`CalcTempBus]          temp_m1_20_25_r;
wire signed [`CalcTempBus]          temp_m1_20_25_i;
wire signed [`CalcTempBus]          temp_m1_20_26_r;
wire signed [`CalcTempBus]          temp_m1_20_26_i;
wire signed [`CalcTempBus]          temp_m1_20_27_r;
wire signed [`CalcTempBus]          temp_m1_20_27_i;
wire signed [`CalcTempBus]          temp_m1_20_28_r;
wire signed [`CalcTempBus]          temp_m1_20_28_i;
wire signed [`CalcTempBus]          temp_m1_20_29_r;
wire signed [`CalcTempBus]          temp_m1_20_29_i;
wire signed [`CalcTempBus]          temp_m1_20_30_r;
wire signed [`CalcTempBus]          temp_m1_20_30_i;
wire signed [`CalcTempBus]          temp_m1_20_31_r;
wire signed [`CalcTempBus]          temp_m1_20_31_i;
wire signed [`CalcTempBus]          temp_m1_20_32_r;
wire signed [`CalcTempBus]          temp_m1_20_32_i;
wire signed [`CalcTempBus]          temp_m1_21_1_r;
wire signed [`CalcTempBus]          temp_m1_21_1_i;
wire signed [`CalcTempBus]          temp_m1_21_2_r;
wire signed [`CalcTempBus]          temp_m1_21_2_i;
wire signed [`CalcTempBus]          temp_m1_21_3_r;
wire signed [`CalcTempBus]          temp_m1_21_3_i;
wire signed [`CalcTempBus]          temp_m1_21_4_r;
wire signed [`CalcTempBus]          temp_m1_21_4_i;
wire signed [`CalcTempBus]          temp_m1_21_5_r;
wire signed [`CalcTempBus]          temp_m1_21_5_i;
wire signed [`CalcTempBus]          temp_m1_21_6_r;
wire signed [`CalcTempBus]          temp_m1_21_6_i;
wire signed [`CalcTempBus]          temp_m1_21_7_r;
wire signed [`CalcTempBus]          temp_m1_21_7_i;
wire signed [`CalcTempBus]          temp_m1_21_8_r;
wire signed [`CalcTempBus]          temp_m1_21_8_i;
wire signed [`CalcTempBus]          temp_m1_21_9_r;
wire signed [`CalcTempBus]          temp_m1_21_9_i;
wire signed [`CalcTempBus]          temp_m1_21_10_r;
wire signed [`CalcTempBus]          temp_m1_21_10_i;
wire signed [`CalcTempBus]          temp_m1_21_11_r;
wire signed [`CalcTempBus]          temp_m1_21_11_i;
wire signed [`CalcTempBus]          temp_m1_21_12_r;
wire signed [`CalcTempBus]          temp_m1_21_12_i;
wire signed [`CalcTempBus]          temp_m1_21_13_r;
wire signed [`CalcTempBus]          temp_m1_21_13_i;
wire signed [`CalcTempBus]          temp_m1_21_14_r;
wire signed [`CalcTempBus]          temp_m1_21_14_i;
wire signed [`CalcTempBus]          temp_m1_21_15_r;
wire signed [`CalcTempBus]          temp_m1_21_15_i;
wire signed [`CalcTempBus]          temp_m1_21_16_r;
wire signed [`CalcTempBus]          temp_m1_21_16_i;
wire signed [`CalcTempBus]          temp_m1_21_17_r;
wire signed [`CalcTempBus]          temp_m1_21_17_i;
wire signed [`CalcTempBus]          temp_m1_21_18_r;
wire signed [`CalcTempBus]          temp_m1_21_18_i;
wire signed [`CalcTempBus]          temp_m1_21_19_r;
wire signed [`CalcTempBus]          temp_m1_21_19_i;
wire signed [`CalcTempBus]          temp_m1_21_20_r;
wire signed [`CalcTempBus]          temp_m1_21_20_i;
wire signed [`CalcTempBus]          temp_m1_21_21_r;
wire signed [`CalcTempBus]          temp_m1_21_21_i;
wire signed [`CalcTempBus]          temp_m1_21_22_r;
wire signed [`CalcTempBus]          temp_m1_21_22_i;
wire signed [`CalcTempBus]          temp_m1_21_23_r;
wire signed [`CalcTempBus]          temp_m1_21_23_i;
wire signed [`CalcTempBus]          temp_m1_21_24_r;
wire signed [`CalcTempBus]          temp_m1_21_24_i;
wire signed [`CalcTempBus]          temp_m1_21_25_r;
wire signed [`CalcTempBus]          temp_m1_21_25_i;
wire signed [`CalcTempBus]          temp_m1_21_26_r;
wire signed [`CalcTempBus]          temp_m1_21_26_i;
wire signed [`CalcTempBus]          temp_m1_21_27_r;
wire signed [`CalcTempBus]          temp_m1_21_27_i;
wire signed [`CalcTempBus]          temp_m1_21_28_r;
wire signed [`CalcTempBus]          temp_m1_21_28_i;
wire signed [`CalcTempBus]          temp_m1_21_29_r;
wire signed [`CalcTempBus]          temp_m1_21_29_i;
wire signed [`CalcTempBus]          temp_m1_21_30_r;
wire signed [`CalcTempBus]          temp_m1_21_30_i;
wire signed [`CalcTempBus]          temp_m1_21_31_r;
wire signed [`CalcTempBus]          temp_m1_21_31_i;
wire signed [`CalcTempBus]          temp_m1_21_32_r;
wire signed [`CalcTempBus]          temp_m1_21_32_i;
wire signed [`CalcTempBus]          temp_m1_22_1_r;
wire signed [`CalcTempBus]          temp_m1_22_1_i;
wire signed [`CalcTempBus]          temp_m1_22_2_r;
wire signed [`CalcTempBus]          temp_m1_22_2_i;
wire signed [`CalcTempBus]          temp_m1_22_3_r;
wire signed [`CalcTempBus]          temp_m1_22_3_i;
wire signed [`CalcTempBus]          temp_m1_22_4_r;
wire signed [`CalcTempBus]          temp_m1_22_4_i;
wire signed [`CalcTempBus]          temp_m1_22_5_r;
wire signed [`CalcTempBus]          temp_m1_22_5_i;
wire signed [`CalcTempBus]          temp_m1_22_6_r;
wire signed [`CalcTempBus]          temp_m1_22_6_i;
wire signed [`CalcTempBus]          temp_m1_22_7_r;
wire signed [`CalcTempBus]          temp_m1_22_7_i;
wire signed [`CalcTempBus]          temp_m1_22_8_r;
wire signed [`CalcTempBus]          temp_m1_22_8_i;
wire signed [`CalcTempBus]          temp_m1_22_9_r;
wire signed [`CalcTempBus]          temp_m1_22_9_i;
wire signed [`CalcTempBus]          temp_m1_22_10_r;
wire signed [`CalcTempBus]          temp_m1_22_10_i;
wire signed [`CalcTempBus]          temp_m1_22_11_r;
wire signed [`CalcTempBus]          temp_m1_22_11_i;
wire signed [`CalcTempBus]          temp_m1_22_12_r;
wire signed [`CalcTempBus]          temp_m1_22_12_i;
wire signed [`CalcTempBus]          temp_m1_22_13_r;
wire signed [`CalcTempBus]          temp_m1_22_13_i;
wire signed [`CalcTempBus]          temp_m1_22_14_r;
wire signed [`CalcTempBus]          temp_m1_22_14_i;
wire signed [`CalcTempBus]          temp_m1_22_15_r;
wire signed [`CalcTempBus]          temp_m1_22_15_i;
wire signed [`CalcTempBus]          temp_m1_22_16_r;
wire signed [`CalcTempBus]          temp_m1_22_16_i;
wire signed [`CalcTempBus]          temp_m1_22_17_r;
wire signed [`CalcTempBus]          temp_m1_22_17_i;
wire signed [`CalcTempBus]          temp_m1_22_18_r;
wire signed [`CalcTempBus]          temp_m1_22_18_i;
wire signed [`CalcTempBus]          temp_m1_22_19_r;
wire signed [`CalcTempBus]          temp_m1_22_19_i;
wire signed [`CalcTempBus]          temp_m1_22_20_r;
wire signed [`CalcTempBus]          temp_m1_22_20_i;
wire signed [`CalcTempBus]          temp_m1_22_21_r;
wire signed [`CalcTempBus]          temp_m1_22_21_i;
wire signed [`CalcTempBus]          temp_m1_22_22_r;
wire signed [`CalcTempBus]          temp_m1_22_22_i;
wire signed [`CalcTempBus]          temp_m1_22_23_r;
wire signed [`CalcTempBus]          temp_m1_22_23_i;
wire signed [`CalcTempBus]          temp_m1_22_24_r;
wire signed [`CalcTempBus]          temp_m1_22_24_i;
wire signed [`CalcTempBus]          temp_m1_22_25_r;
wire signed [`CalcTempBus]          temp_m1_22_25_i;
wire signed [`CalcTempBus]          temp_m1_22_26_r;
wire signed [`CalcTempBus]          temp_m1_22_26_i;
wire signed [`CalcTempBus]          temp_m1_22_27_r;
wire signed [`CalcTempBus]          temp_m1_22_27_i;
wire signed [`CalcTempBus]          temp_m1_22_28_r;
wire signed [`CalcTempBus]          temp_m1_22_28_i;
wire signed [`CalcTempBus]          temp_m1_22_29_r;
wire signed [`CalcTempBus]          temp_m1_22_29_i;
wire signed [`CalcTempBus]          temp_m1_22_30_r;
wire signed [`CalcTempBus]          temp_m1_22_30_i;
wire signed [`CalcTempBus]          temp_m1_22_31_r;
wire signed [`CalcTempBus]          temp_m1_22_31_i;
wire signed [`CalcTempBus]          temp_m1_22_32_r;
wire signed [`CalcTempBus]          temp_m1_22_32_i;
wire signed [`CalcTempBus]          temp_m1_23_1_r;
wire signed [`CalcTempBus]          temp_m1_23_1_i;
wire signed [`CalcTempBus]          temp_m1_23_2_r;
wire signed [`CalcTempBus]          temp_m1_23_2_i;
wire signed [`CalcTempBus]          temp_m1_23_3_r;
wire signed [`CalcTempBus]          temp_m1_23_3_i;
wire signed [`CalcTempBus]          temp_m1_23_4_r;
wire signed [`CalcTempBus]          temp_m1_23_4_i;
wire signed [`CalcTempBus]          temp_m1_23_5_r;
wire signed [`CalcTempBus]          temp_m1_23_5_i;
wire signed [`CalcTempBus]          temp_m1_23_6_r;
wire signed [`CalcTempBus]          temp_m1_23_6_i;
wire signed [`CalcTempBus]          temp_m1_23_7_r;
wire signed [`CalcTempBus]          temp_m1_23_7_i;
wire signed [`CalcTempBus]          temp_m1_23_8_r;
wire signed [`CalcTempBus]          temp_m1_23_8_i;
wire signed [`CalcTempBus]          temp_m1_23_9_r;
wire signed [`CalcTempBus]          temp_m1_23_9_i;
wire signed [`CalcTempBus]          temp_m1_23_10_r;
wire signed [`CalcTempBus]          temp_m1_23_10_i;
wire signed [`CalcTempBus]          temp_m1_23_11_r;
wire signed [`CalcTempBus]          temp_m1_23_11_i;
wire signed [`CalcTempBus]          temp_m1_23_12_r;
wire signed [`CalcTempBus]          temp_m1_23_12_i;
wire signed [`CalcTempBus]          temp_m1_23_13_r;
wire signed [`CalcTempBus]          temp_m1_23_13_i;
wire signed [`CalcTempBus]          temp_m1_23_14_r;
wire signed [`CalcTempBus]          temp_m1_23_14_i;
wire signed [`CalcTempBus]          temp_m1_23_15_r;
wire signed [`CalcTempBus]          temp_m1_23_15_i;
wire signed [`CalcTempBus]          temp_m1_23_16_r;
wire signed [`CalcTempBus]          temp_m1_23_16_i;
wire signed [`CalcTempBus]          temp_m1_23_17_r;
wire signed [`CalcTempBus]          temp_m1_23_17_i;
wire signed [`CalcTempBus]          temp_m1_23_18_r;
wire signed [`CalcTempBus]          temp_m1_23_18_i;
wire signed [`CalcTempBus]          temp_m1_23_19_r;
wire signed [`CalcTempBus]          temp_m1_23_19_i;
wire signed [`CalcTempBus]          temp_m1_23_20_r;
wire signed [`CalcTempBus]          temp_m1_23_20_i;
wire signed [`CalcTempBus]          temp_m1_23_21_r;
wire signed [`CalcTempBus]          temp_m1_23_21_i;
wire signed [`CalcTempBus]          temp_m1_23_22_r;
wire signed [`CalcTempBus]          temp_m1_23_22_i;
wire signed [`CalcTempBus]          temp_m1_23_23_r;
wire signed [`CalcTempBus]          temp_m1_23_23_i;
wire signed [`CalcTempBus]          temp_m1_23_24_r;
wire signed [`CalcTempBus]          temp_m1_23_24_i;
wire signed [`CalcTempBus]          temp_m1_23_25_r;
wire signed [`CalcTempBus]          temp_m1_23_25_i;
wire signed [`CalcTempBus]          temp_m1_23_26_r;
wire signed [`CalcTempBus]          temp_m1_23_26_i;
wire signed [`CalcTempBus]          temp_m1_23_27_r;
wire signed [`CalcTempBus]          temp_m1_23_27_i;
wire signed [`CalcTempBus]          temp_m1_23_28_r;
wire signed [`CalcTempBus]          temp_m1_23_28_i;
wire signed [`CalcTempBus]          temp_m1_23_29_r;
wire signed [`CalcTempBus]          temp_m1_23_29_i;
wire signed [`CalcTempBus]          temp_m1_23_30_r;
wire signed [`CalcTempBus]          temp_m1_23_30_i;
wire signed [`CalcTempBus]          temp_m1_23_31_r;
wire signed [`CalcTempBus]          temp_m1_23_31_i;
wire signed [`CalcTempBus]          temp_m1_23_32_r;
wire signed [`CalcTempBus]          temp_m1_23_32_i;
wire signed [`CalcTempBus]          temp_m1_24_1_r;
wire signed [`CalcTempBus]          temp_m1_24_1_i;
wire signed [`CalcTempBus]          temp_m1_24_2_r;
wire signed [`CalcTempBus]          temp_m1_24_2_i;
wire signed [`CalcTempBus]          temp_m1_24_3_r;
wire signed [`CalcTempBus]          temp_m1_24_3_i;
wire signed [`CalcTempBus]          temp_m1_24_4_r;
wire signed [`CalcTempBus]          temp_m1_24_4_i;
wire signed [`CalcTempBus]          temp_m1_24_5_r;
wire signed [`CalcTempBus]          temp_m1_24_5_i;
wire signed [`CalcTempBus]          temp_m1_24_6_r;
wire signed [`CalcTempBus]          temp_m1_24_6_i;
wire signed [`CalcTempBus]          temp_m1_24_7_r;
wire signed [`CalcTempBus]          temp_m1_24_7_i;
wire signed [`CalcTempBus]          temp_m1_24_8_r;
wire signed [`CalcTempBus]          temp_m1_24_8_i;
wire signed [`CalcTempBus]          temp_m1_24_9_r;
wire signed [`CalcTempBus]          temp_m1_24_9_i;
wire signed [`CalcTempBus]          temp_m1_24_10_r;
wire signed [`CalcTempBus]          temp_m1_24_10_i;
wire signed [`CalcTempBus]          temp_m1_24_11_r;
wire signed [`CalcTempBus]          temp_m1_24_11_i;
wire signed [`CalcTempBus]          temp_m1_24_12_r;
wire signed [`CalcTempBus]          temp_m1_24_12_i;
wire signed [`CalcTempBus]          temp_m1_24_13_r;
wire signed [`CalcTempBus]          temp_m1_24_13_i;
wire signed [`CalcTempBus]          temp_m1_24_14_r;
wire signed [`CalcTempBus]          temp_m1_24_14_i;
wire signed [`CalcTempBus]          temp_m1_24_15_r;
wire signed [`CalcTempBus]          temp_m1_24_15_i;
wire signed [`CalcTempBus]          temp_m1_24_16_r;
wire signed [`CalcTempBus]          temp_m1_24_16_i;
wire signed [`CalcTempBus]          temp_m1_24_17_r;
wire signed [`CalcTempBus]          temp_m1_24_17_i;
wire signed [`CalcTempBus]          temp_m1_24_18_r;
wire signed [`CalcTempBus]          temp_m1_24_18_i;
wire signed [`CalcTempBus]          temp_m1_24_19_r;
wire signed [`CalcTempBus]          temp_m1_24_19_i;
wire signed [`CalcTempBus]          temp_m1_24_20_r;
wire signed [`CalcTempBus]          temp_m1_24_20_i;
wire signed [`CalcTempBus]          temp_m1_24_21_r;
wire signed [`CalcTempBus]          temp_m1_24_21_i;
wire signed [`CalcTempBus]          temp_m1_24_22_r;
wire signed [`CalcTempBus]          temp_m1_24_22_i;
wire signed [`CalcTempBus]          temp_m1_24_23_r;
wire signed [`CalcTempBus]          temp_m1_24_23_i;
wire signed [`CalcTempBus]          temp_m1_24_24_r;
wire signed [`CalcTempBus]          temp_m1_24_24_i;
wire signed [`CalcTempBus]          temp_m1_24_25_r;
wire signed [`CalcTempBus]          temp_m1_24_25_i;
wire signed [`CalcTempBus]          temp_m1_24_26_r;
wire signed [`CalcTempBus]          temp_m1_24_26_i;
wire signed [`CalcTempBus]          temp_m1_24_27_r;
wire signed [`CalcTempBus]          temp_m1_24_27_i;
wire signed [`CalcTempBus]          temp_m1_24_28_r;
wire signed [`CalcTempBus]          temp_m1_24_28_i;
wire signed [`CalcTempBus]          temp_m1_24_29_r;
wire signed [`CalcTempBus]          temp_m1_24_29_i;
wire signed [`CalcTempBus]          temp_m1_24_30_r;
wire signed [`CalcTempBus]          temp_m1_24_30_i;
wire signed [`CalcTempBus]          temp_m1_24_31_r;
wire signed [`CalcTempBus]          temp_m1_24_31_i;
wire signed [`CalcTempBus]          temp_m1_24_32_r;
wire signed [`CalcTempBus]          temp_m1_24_32_i;
wire signed [`CalcTempBus]          temp_m1_25_1_r;
wire signed [`CalcTempBus]          temp_m1_25_1_i;
wire signed [`CalcTempBus]          temp_m1_25_2_r;
wire signed [`CalcTempBus]          temp_m1_25_2_i;
wire signed [`CalcTempBus]          temp_m1_25_3_r;
wire signed [`CalcTempBus]          temp_m1_25_3_i;
wire signed [`CalcTempBus]          temp_m1_25_4_r;
wire signed [`CalcTempBus]          temp_m1_25_4_i;
wire signed [`CalcTempBus]          temp_m1_25_5_r;
wire signed [`CalcTempBus]          temp_m1_25_5_i;
wire signed [`CalcTempBus]          temp_m1_25_6_r;
wire signed [`CalcTempBus]          temp_m1_25_6_i;
wire signed [`CalcTempBus]          temp_m1_25_7_r;
wire signed [`CalcTempBus]          temp_m1_25_7_i;
wire signed [`CalcTempBus]          temp_m1_25_8_r;
wire signed [`CalcTempBus]          temp_m1_25_8_i;
wire signed [`CalcTempBus]          temp_m1_25_9_r;
wire signed [`CalcTempBus]          temp_m1_25_9_i;
wire signed [`CalcTempBus]          temp_m1_25_10_r;
wire signed [`CalcTempBus]          temp_m1_25_10_i;
wire signed [`CalcTempBus]          temp_m1_25_11_r;
wire signed [`CalcTempBus]          temp_m1_25_11_i;
wire signed [`CalcTempBus]          temp_m1_25_12_r;
wire signed [`CalcTempBus]          temp_m1_25_12_i;
wire signed [`CalcTempBus]          temp_m1_25_13_r;
wire signed [`CalcTempBus]          temp_m1_25_13_i;
wire signed [`CalcTempBus]          temp_m1_25_14_r;
wire signed [`CalcTempBus]          temp_m1_25_14_i;
wire signed [`CalcTempBus]          temp_m1_25_15_r;
wire signed [`CalcTempBus]          temp_m1_25_15_i;
wire signed [`CalcTempBus]          temp_m1_25_16_r;
wire signed [`CalcTempBus]          temp_m1_25_16_i;
wire signed [`CalcTempBus]          temp_m1_25_17_r;
wire signed [`CalcTempBus]          temp_m1_25_17_i;
wire signed [`CalcTempBus]          temp_m1_25_18_r;
wire signed [`CalcTempBus]          temp_m1_25_18_i;
wire signed [`CalcTempBus]          temp_m1_25_19_r;
wire signed [`CalcTempBus]          temp_m1_25_19_i;
wire signed [`CalcTempBus]          temp_m1_25_20_r;
wire signed [`CalcTempBus]          temp_m1_25_20_i;
wire signed [`CalcTempBus]          temp_m1_25_21_r;
wire signed [`CalcTempBus]          temp_m1_25_21_i;
wire signed [`CalcTempBus]          temp_m1_25_22_r;
wire signed [`CalcTempBus]          temp_m1_25_22_i;
wire signed [`CalcTempBus]          temp_m1_25_23_r;
wire signed [`CalcTempBus]          temp_m1_25_23_i;
wire signed [`CalcTempBus]          temp_m1_25_24_r;
wire signed [`CalcTempBus]          temp_m1_25_24_i;
wire signed [`CalcTempBus]          temp_m1_25_25_r;
wire signed [`CalcTempBus]          temp_m1_25_25_i;
wire signed [`CalcTempBus]          temp_m1_25_26_r;
wire signed [`CalcTempBus]          temp_m1_25_26_i;
wire signed [`CalcTempBus]          temp_m1_25_27_r;
wire signed [`CalcTempBus]          temp_m1_25_27_i;
wire signed [`CalcTempBus]          temp_m1_25_28_r;
wire signed [`CalcTempBus]          temp_m1_25_28_i;
wire signed [`CalcTempBus]          temp_m1_25_29_r;
wire signed [`CalcTempBus]          temp_m1_25_29_i;
wire signed [`CalcTempBus]          temp_m1_25_30_r;
wire signed [`CalcTempBus]          temp_m1_25_30_i;
wire signed [`CalcTempBus]          temp_m1_25_31_r;
wire signed [`CalcTempBus]          temp_m1_25_31_i;
wire signed [`CalcTempBus]          temp_m1_25_32_r;
wire signed [`CalcTempBus]          temp_m1_25_32_i;
wire signed [`CalcTempBus]          temp_m1_26_1_r;
wire signed [`CalcTempBus]          temp_m1_26_1_i;
wire signed [`CalcTempBus]          temp_m1_26_2_r;
wire signed [`CalcTempBus]          temp_m1_26_2_i;
wire signed [`CalcTempBus]          temp_m1_26_3_r;
wire signed [`CalcTempBus]          temp_m1_26_3_i;
wire signed [`CalcTempBus]          temp_m1_26_4_r;
wire signed [`CalcTempBus]          temp_m1_26_4_i;
wire signed [`CalcTempBus]          temp_m1_26_5_r;
wire signed [`CalcTempBus]          temp_m1_26_5_i;
wire signed [`CalcTempBus]          temp_m1_26_6_r;
wire signed [`CalcTempBus]          temp_m1_26_6_i;
wire signed [`CalcTempBus]          temp_m1_26_7_r;
wire signed [`CalcTempBus]          temp_m1_26_7_i;
wire signed [`CalcTempBus]          temp_m1_26_8_r;
wire signed [`CalcTempBus]          temp_m1_26_8_i;
wire signed [`CalcTempBus]          temp_m1_26_9_r;
wire signed [`CalcTempBus]          temp_m1_26_9_i;
wire signed [`CalcTempBus]          temp_m1_26_10_r;
wire signed [`CalcTempBus]          temp_m1_26_10_i;
wire signed [`CalcTempBus]          temp_m1_26_11_r;
wire signed [`CalcTempBus]          temp_m1_26_11_i;
wire signed [`CalcTempBus]          temp_m1_26_12_r;
wire signed [`CalcTempBus]          temp_m1_26_12_i;
wire signed [`CalcTempBus]          temp_m1_26_13_r;
wire signed [`CalcTempBus]          temp_m1_26_13_i;
wire signed [`CalcTempBus]          temp_m1_26_14_r;
wire signed [`CalcTempBus]          temp_m1_26_14_i;
wire signed [`CalcTempBus]          temp_m1_26_15_r;
wire signed [`CalcTempBus]          temp_m1_26_15_i;
wire signed [`CalcTempBus]          temp_m1_26_16_r;
wire signed [`CalcTempBus]          temp_m1_26_16_i;
wire signed [`CalcTempBus]          temp_m1_26_17_r;
wire signed [`CalcTempBus]          temp_m1_26_17_i;
wire signed [`CalcTempBus]          temp_m1_26_18_r;
wire signed [`CalcTempBus]          temp_m1_26_18_i;
wire signed [`CalcTempBus]          temp_m1_26_19_r;
wire signed [`CalcTempBus]          temp_m1_26_19_i;
wire signed [`CalcTempBus]          temp_m1_26_20_r;
wire signed [`CalcTempBus]          temp_m1_26_20_i;
wire signed [`CalcTempBus]          temp_m1_26_21_r;
wire signed [`CalcTempBus]          temp_m1_26_21_i;
wire signed [`CalcTempBus]          temp_m1_26_22_r;
wire signed [`CalcTempBus]          temp_m1_26_22_i;
wire signed [`CalcTempBus]          temp_m1_26_23_r;
wire signed [`CalcTempBus]          temp_m1_26_23_i;
wire signed [`CalcTempBus]          temp_m1_26_24_r;
wire signed [`CalcTempBus]          temp_m1_26_24_i;
wire signed [`CalcTempBus]          temp_m1_26_25_r;
wire signed [`CalcTempBus]          temp_m1_26_25_i;
wire signed [`CalcTempBus]          temp_m1_26_26_r;
wire signed [`CalcTempBus]          temp_m1_26_26_i;
wire signed [`CalcTempBus]          temp_m1_26_27_r;
wire signed [`CalcTempBus]          temp_m1_26_27_i;
wire signed [`CalcTempBus]          temp_m1_26_28_r;
wire signed [`CalcTempBus]          temp_m1_26_28_i;
wire signed [`CalcTempBus]          temp_m1_26_29_r;
wire signed [`CalcTempBus]          temp_m1_26_29_i;
wire signed [`CalcTempBus]          temp_m1_26_30_r;
wire signed [`CalcTempBus]          temp_m1_26_30_i;
wire signed [`CalcTempBus]          temp_m1_26_31_r;
wire signed [`CalcTempBus]          temp_m1_26_31_i;
wire signed [`CalcTempBus]          temp_m1_26_32_r;
wire signed [`CalcTempBus]          temp_m1_26_32_i;
wire signed [`CalcTempBus]          temp_m1_27_1_r;
wire signed [`CalcTempBus]          temp_m1_27_1_i;
wire signed [`CalcTempBus]          temp_m1_27_2_r;
wire signed [`CalcTempBus]          temp_m1_27_2_i;
wire signed [`CalcTempBus]          temp_m1_27_3_r;
wire signed [`CalcTempBus]          temp_m1_27_3_i;
wire signed [`CalcTempBus]          temp_m1_27_4_r;
wire signed [`CalcTempBus]          temp_m1_27_4_i;
wire signed [`CalcTempBus]          temp_m1_27_5_r;
wire signed [`CalcTempBus]          temp_m1_27_5_i;
wire signed [`CalcTempBus]          temp_m1_27_6_r;
wire signed [`CalcTempBus]          temp_m1_27_6_i;
wire signed [`CalcTempBus]          temp_m1_27_7_r;
wire signed [`CalcTempBus]          temp_m1_27_7_i;
wire signed [`CalcTempBus]          temp_m1_27_8_r;
wire signed [`CalcTempBus]          temp_m1_27_8_i;
wire signed [`CalcTempBus]          temp_m1_27_9_r;
wire signed [`CalcTempBus]          temp_m1_27_9_i;
wire signed [`CalcTempBus]          temp_m1_27_10_r;
wire signed [`CalcTempBus]          temp_m1_27_10_i;
wire signed [`CalcTempBus]          temp_m1_27_11_r;
wire signed [`CalcTempBus]          temp_m1_27_11_i;
wire signed [`CalcTempBus]          temp_m1_27_12_r;
wire signed [`CalcTempBus]          temp_m1_27_12_i;
wire signed [`CalcTempBus]          temp_m1_27_13_r;
wire signed [`CalcTempBus]          temp_m1_27_13_i;
wire signed [`CalcTempBus]          temp_m1_27_14_r;
wire signed [`CalcTempBus]          temp_m1_27_14_i;
wire signed [`CalcTempBus]          temp_m1_27_15_r;
wire signed [`CalcTempBus]          temp_m1_27_15_i;
wire signed [`CalcTempBus]          temp_m1_27_16_r;
wire signed [`CalcTempBus]          temp_m1_27_16_i;
wire signed [`CalcTempBus]          temp_m1_27_17_r;
wire signed [`CalcTempBus]          temp_m1_27_17_i;
wire signed [`CalcTempBus]          temp_m1_27_18_r;
wire signed [`CalcTempBus]          temp_m1_27_18_i;
wire signed [`CalcTempBus]          temp_m1_27_19_r;
wire signed [`CalcTempBus]          temp_m1_27_19_i;
wire signed [`CalcTempBus]          temp_m1_27_20_r;
wire signed [`CalcTempBus]          temp_m1_27_20_i;
wire signed [`CalcTempBus]          temp_m1_27_21_r;
wire signed [`CalcTempBus]          temp_m1_27_21_i;
wire signed [`CalcTempBus]          temp_m1_27_22_r;
wire signed [`CalcTempBus]          temp_m1_27_22_i;
wire signed [`CalcTempBus]          temp_m1_27_23_r;
wire signed [`CalcTempBus]          temp_m1_27_23_i;
wire signed [`CalcTempBus]          temp_m1_27_24_r;
wire signed [`CalcTempBus]          temp_m1_27_24_i;
wire signed [`CalcTempBus]          temp_m1_27_25_r;
wire signed [`CalcTempBus]          temp_m1_27_25_i;
wire signed [`CalcTempBus]          temp_m1_27_26_r;
wire signed [`CalcTempBus]          temp_m1_27_26_i;
wire signed [`CalcTempBus]          temp_m1_27_27_r;
wire signed [`CalcTempBus]          temp_m1_27_27_i;
wire signed [`CalcTempBus]          temp_m1_27_28_r;
wire signed [`CalcTempBus]          temp_m1_27_28_i;
wire signed [`CalcTempBus]          temp_m1_27_29_r;
wire signed [`CalcTempBus]          temp_m1_27_29_i;
wire signed [`CalcTempBus]          temp_m1_27_30_r;
wire signed [`CalcTempBus]          temp_m1_27_30_i;
wire signed [`CalcTempBus]          temp_m1_27_31_r;
wire signed [`CalcTempBus]          temp_m1_27_31_i;
wire signed [`CalcTempBus]          temp_m1_27_32_r;
wire signed [`CalcTempBus]          temp_m1_27_32_i;
wire signed [`CalcTempBus]          temp_m1_28_1_r;
wire signed [`CalcTempBus]          temp_m1_28_1_i;
wire signed [`CalcTempBus]          temp_m1_28_2_r;
wire signed [`CalcTempBus]          temp_m1_28_2_i;
wire signed [`CalcTempBus]          temp_m1_28_3_r;
wire signed [`CalcTempBus]          temp_m1_28_3_i;
wire signed [`CalcTempBus]          temp_m1_28_4_r;
wire signed [`CalcTempBus]          temp_m1_28_4_i;
wire signed [`CalcTempBus]          temp_m1_28_5_r;
wire signed [`CalcTempBus]          temp_m1_28_5_i;
wire signed [`CalcTempBus]          temp_m1_28_6_r;
wire signed [`CalcTempBus]          temp_m1_28_6_i;
wire signed [`CalcTempBus]          temp_m1_28_7_r;
wire signed [`CalcTempBus]          temp_m1_28_7_i;
wire signed [`CalcTempBus]          temp_m1_28_8_r;
wire signed [`CalcTempBus]          temp_m1_28_8_i;
wire signed [`CalcTempBus]          temp_m1_28_9_r;
wire signed [`CalcTempBus]          temp_m1_28_9_i;
wire signed [`CalcTempBus]          temp_m1_28_10_r;
wire signed [`CalcTempBus]          temp_m1_28_10_i;
wire signed [`CalcTempBus]          temp_m1_28_11_r;
wire signed [`CalcTempBus]          temp_m1_28_11_i;
wire signed [`CalcTempBus]          temp_m1_28_12_r;
wire signed [`CalcTempBus]          temp_m1_28_12_i;
wire signed [`CalcTempBus]          temp_m1_28_13_r;
wire signed [`CalcTempBus]          temp_m1_28_13_i;
wire signed [`CalcTempBus]          temp_m1_28_14_r;
wire signed [`CalcTempBus]          temp_m1_28_14_i;
wire signed [`CalcTempBus]          temp_m1_28_15_r;
wire signed [`CalcTempBus]          temp_m1_28_15_i;
wire signed [`CalcTempBus]          temp_m1_28_16_r;
wire signed [`CalcTempBus]          temp_m1_28_16_i;
wire signed [`CalcTempBus]          temp_m1_28_17_r;
wire signed [`CalcTempBus]          temp_m1_28_17_i;
wire signed [`CalcTempBus]          temp_m1_28_18_r;
wire signed [`CalcTempBus]          temp_m1_28_18_i;
wire signed [`CalcTempBus]          temp_m1_28_19_r;
wire signed [`CalcTempBus]          temp_m1_28_19_i;
wire signed [`CalcTempBus]          temp_m1_28_20_r;
wire signed [`CalcTempBus]          temp_m1_28_20_i;
wire signed [`CalcTempBus]          temp_m1_28_21_r;
wire signed [`CalcTempBus]          temp_m1_28_21_i;
wire signed [`CalcTempBus]          temp_m1_28_22_r;
wire signed [`CalcTempBus]          temp_m1_28_22_i;
wire signed [`CalcTempBus]          temp_m1_28_23_r;
wire signed [`CalcTempBus]          temp_m1_28_23_i;
wire signed [`CalcTempBus]          temp_m1_28_24_r;
wire signed [`CalcTempBus]          temp_m1_28_24_i;
wire signed [`CalcTempBus]          temp_m1_28_25_r;
wire signed [`CalcTempBus]          temp_m1_28_25_i;
wire signed [`CalcTempBus]          temp_m1_28_26_r;
wire signed [`CalcTempBus]          temp_m1_28_26_i;
wire signed [`CalcTempBus]          temp_m1_28_27_r;
wire signed [`CalcTempBus]          temp_m1_28_27_i;
wire signed [`CalcTempBus]          temp_m1_28_28_r;
wire signed [`CalcTempBus]          temp_m1_28_28_i;
wire signed [`CalcTempBus]          temp_m1_28_29_r;
wire signed [`CalcTempBus]          temp_m1_28_29_i;
wire signed [`CalcTempBus]          temp_m1_28_30_r;
wire signed [`CalcTempBus]          temp_m1_28_30_i;
wire signed [`CalcTempBus]          temp_m1_28_31_r;
wire signed [`CalcTempBus]          temp_m1_28_31_i;
wire signed [`CalcTempBus]          temp_m1_28_32_r;
wire signed [`CalcTempBus]          temp_m1_28_32_i;
wire signed [`CalcTempBus]          temp_m1_29_1_r;
wire signed [`CalcTempBus]          temp_m1_29_1_i;
wire signed [`CalcTempBus]          temp_m1_29_2_r;
wire signed [`CalcTempBus]          temp_m1_29_2_i;
wire signed [`CalcTempBus]          temp_m1_29_3_r;
wire signed [`CalcTempBus]          temp_m1_29_3_i;
wire signed [`CalcTempBus]          temp_m1_29_4_r;
wire signed [`CalcTempBus]          temp_m1_29_4_i;
wire signed [`CalcTempBus]          temp_m1_29_5_r;
wire signed [`CalcTempBus]          temp_m1_29_5_i;
wire signed [`CalcTempBus]          temp_m1_29_6_r;
wire signed [`CalcTempBus]          temp_m1_29_6_i;
wire signed [`CalcTempBus]          temp_m1_29_7_r;
wire signed [`CalcTempBus]          temp_m1_29_7_i;
wire signed [`CalcTempBus]          temp_m1_29_8_r;
wire signed [`CalcTempBus]          temp_m1_29_8_i;
wire signed [`CalcTempBus]          temp_m1_29_9_r;
wire signed [`CalcTempBus]          temp_m1_29_9_i;
wire signed [`CalcTempBus]          temp_m1_29_10_r;
wire signed [`CalcTempBus]          temp_m1_29_10_i;
wire signed [`CalcTempBus]          temp_m1_29_11_r;
wire signed [`CalcTempBus]          temp_m1_29_11_i;
wire signed [`CalcTempBus]          temp_m1_29_12_r;
wire signed [`CalcTempBus]          temp_m1_29_12_i;
wire signed [`CalcTempBus]          temp_m1_29_13_r;
wire signed [`CalcTempBus]          temp_m1_29_13_i;
wire signed [`CalcTempBus]          temp_m1_29_14_r;
wire signed [`CalcTempBus]          temp_m1_29_14_i;
wire signed [`CalcTempBus]          temp_m1_29_15_r;
wire signed [`CalcTempBus]          temp_m1_29_15_i;
wire signed [`CalcTempBus]          temp_m1_29_16_r;
wire signed [`CalcTempBus]          temp_m1_29_16_i;
wire signed [`CalcTempBus]          temp_m1_29_17_r;
wire signed [`CalcTempBus]          temp_m1_29_17_i;
wire signed [`CalcTempBus]          temp_m1_29_18_r;
wire signed [`CalcTempBus]          temp_m1_29_18_i;
wire signed [`CalcTempBus]          temp_m1_29_19_r;
wire signed [`CalcTempBus]          temp_m1_29_19_i;
wire signed [`CalcTempBus]          temp_m1_29_20_r;
wire signed [`CalcTempBus]          temp_m1_29_20_i;
wire signed [`CalcTempBus]          temp_m1_29_21_r;
wire signed [`CalcTempBus]          temp_m1_29_21_i;
wire signed [`CalcTempBus]          temp_m1_29_22_r;
wire signed [`CalcTempBus]          temp_m1_29_22_i;
wire signed [`CalcTempBus]          temp_m1_29_23_r;
wire signed [`CalcTempBus]          temp_m1_29_23_i;
wire signed [`CalcTempBus]          temp_m1_29_24_r;
wire signed [`CalcTempBus]          temp_m1_29_24_i;
wire signed [`CalcTempBus]          temp_m1_29_25_r;
wire signed [`CalcTempBus]          temp_m1_29_25_i;
wire signed [`CalcTempBus]          temp_m1_29_26_r;
wire signed [`CalcTempBus]          temp_m1_29_26_i;
wire signed [`CalcTempBus]          temp_m1_29_27_r;
wire signed [`CalcTempBus]          temp_m1_29_27_i;
wire signed [`CalcTempBus]          temp_m1_29_28_r;
wire signed [`CalcTempBus]          temp_m1_29_28_i;
wire signed [`CalcTempBus]          temp_m1_29_29_r;
wire signed [`CalcTempBus]          temp_m1_29_29_i;
wire signed [`CalcTempBus]          temp_m1_29_30_r;
wire signed [`CalcTempBus]          temp_m1_29_30_i;
wire signed [`CalcTempBus]          temp_m1_29_31_r;
wire signed [`CalcTempBus]          temp_m1_29_31_i;
wire signed [`CalcTempBus]          temp_m1_29_32_r;
wire signed [`CalcTempBus]          temp_m1_29_32_i;
wire signed [`CalcTempBus]          temp_m1_30_1_r;
wire signed [`CalcTempBus]          temp_m1_30_1_i;
wire signed [`CalcTempBus]          temp_m1_30_2_r;
wire signed [`CalcTempBus]          temp_m1_30_2_i;
wire signed [`CalcTempBus]          temp_m1_30_3_r;
wire signed [`CalcTempBus]          temp_m1_30_3_i;
wire signed [`CalcTempBus]          temp_m1_30_4_r;
wire signed [`CalcTempBus]          temp_m1_30_4_i;
wire signed [`CalcTempBus]          temp_m1_30_5_r;
wire signed [`CalcTempBus]          temp_m1_30_5_i;
wire signed [`CalcTempBus]          temp_m1_30_6_r;
wire signed [`CalcTempBus]          temp_m1_30_6_i;
wire signed [`CalcTempBus]          temp_m1_30_7_r;
wire signed [`CalcTempBus]          temp_m1_30_7_i;
wire signed [`CalcTempBus]          temp_m1_30_8_r;
wire signed [`CalcTempBus]          temp_m1_30_8_i;
wire signed [`CalcTempBus]          temp_m1_30_9_r;
wire signed [`CalcTempBus]          temp_m1_30_9_i;
wire signed [`CalcTempBus]          temp_m1_30_10_r;
wire signed [`CalcTempBus]          temp_m1_30_10_i;
wire signed [`CalcTempBus]          temp_m1_30_11_r;
wire signed [`CalcTempBus]          temp_m1_30_11_i;
wire signed [`CalcTempBus]          temp_m1_30_12_r;
wire signed [`CalcTempBus]          temp_m1_30_12_i;
wire signed [`CalcTempBus]          temp_m1_30_13_r;
wire signed [`CalcTempBus]          temp_m1_30_13_i;
wire signed [`CalcTempBus]          temp_m1_30_14_r;
wire signed [`CalcTempBus]          temp_m1_30_14_i;
wire signed [`CalcTempBus]          temp_m1_30_15_r;
wire signed [`CalcTempBus]          temp_m1_30_15_i;
wire signed [`CalcTempBus]          temp_m1_30_16_r;
wire signed [`CalcTempBus]          temp_m1_30_16_i;
wire signed [`CalcTempBus]          temp_m1_30_17_r;
wire signed [`CalcTempBus]          temp_m1_30_17_i;
wire signed [`CalcTempBus]          temp_m1_30_18_r;
wire signed [`CalcTempBus]          temp_m1_30_18_i;
wire signed [`CalcTempBus]          temp_m1_30_19_r;
wire signed [`CalcTempBus]          temp_m1_30_19_i;
wire signed [`CalcTempBus]          temp_m1_30_20_r;
wire signed [`CalcTempBus]          temp_m1_30_20_i;
wire signed [`CalcTempBus]          temp_m1_30_21_r;
wire signed [`CalcTempBus]          temp_m1_30_21_i;
wire signed [`CalcTempBus]          temp_m1_30_22_r;
wire signed [`CalcTempBus]          temp_m1_30_22_i;
wire signed [`CalcTempBus]          temp_m1_30_23_r;
wire signed [`CalcTempBus]          temp_m1_30_23_i;
wire signed [`CalcTempBus]          temp_m1_30_24_r;
wire signed [`CalcTempBus]          temp_m1_30_24_i;
wire signed [`CalcTempBus]          temp_m1_30_25_r;
wire signed [`CalcTempBus]          temp_m1_30_25_i;
wire signed [`CalcTempBus]          temp_m1_30_26_r;
wire signed [`CalcTempBus]          temp_m1_30_26_i;
wire signed [`CalcTempBus]          temp_m1_30_27_r;
wire signed [`CalcTempBus]          temp_m1_30_27_i;
wire signed [`CalcTempBus]          temp_m1_30_28_r;
wire signed [`CalcTempBus]          temp_m1_30_28_i;
wire signed [`CalcTempBus]          temp_m1_30_29_r;
wire signed [`CalcTempBus]          temp_m1_30_29_i;
wire signed [`CalcTempBus]          temp_m1_30_30_r;
wire signed [`CalcTempBus]          temp_m1_30_30_i;
wire signed [`CalcTempBus]          temp_m1_30_31_r;
wire signed [`CalcTempBus]          temp_m1_30_31_i;
wire signed [`CalcTempBus]          temp_m1_30_32_r;
wire signed [`CalcTempBus]          temp_m1_30_32_i;
wire signed [`CalcTempBus]          temp_m1_31_1_r;
wire signed [`CalcTempBus]          temp_m1_31_1_i;
wire signed [`CalcTempBus]          temp_m1_31_2_r;
wire signed [`CalcTempBus]          temp_m1_31_2_i;
wire signed [`CalcTempBus]          temp_m1_31_3_r;
wire signed [`CalcTempBus]          temp_m1_31_3_i;
wire signed [`CalcTempBus]          temp_m1_31_4_r;
wire signed [`CalcTempBus]          temp_m1_31_4_i;
wire signed [`CalcTempBus]          temp_m1_31_5_r;
wire signed [`CalcTempBus]          temp_m1_31_5_i;
wire signed [`CalcTempBus]          temp_m1_31_6_r;
wire signed [`CalcTempBus]          temp_m1_31_6_i;
wire signed [`CalcTempBus]          temp_m1_31_7_r;
wire signed [`CalcTempBus]          temp_m1_31_7_i;
wire signed [`CalcTempBus]          temp_m1_31_8_r;
wire signed [`CalcTempBus]          temp_m1_31_8_i;
wire signed [`CalcTempBus]          temp_m1_31_9_r;
wire signed [`CalcTempBus]          temp_m1_31_9_i;
wire signed [`CalcTempBus]          temp_m1_31_10_r;
wire signed [`CalcTempBus]          temp_m1_31_10_i;
wire signed [`CalcTempBus]          temp_m1_31_11_r;
wire signed [`CalcTempBus]          temp_m1_31_11_i;
wire signed [`CalcTempBus]          temp_m1_31_12_r;
wire signed [`CalcTempBus]          temp_m1_31_12_i;
wire signed [`CalcTempBus]          temp_m1_31_13_r;
wire signed [`CalcTempBus]          temp_m1_31_13_i;
wire signed [`CalcTempBus]          temp_m1_31_14_r;
wire signed [`CalcTempBus]          temp_m1_31_14_i;
wire signed [`CalcTempBus]          temp_m1_31_15_r;
wire signed [`CalcTempBus]          temp_m1_31_15_i;
wire signed [`CalcTempBus]          temp_m1_31_16_r;
wire signed [`CalcTempBus]          temp_m1_31_16_i;
wire signed [`CalcTempBus]          temp_m1_31_17_r;
wire signed [`CalcTempBus]          temp_m1_31_17_i;
wire signed [`CalcTempBus]          temp_m1_31_18_r;
wire signed [`CalcTempBus]          temp_m1_31_18_i;
wire signed [`CalcTempBus]          temp_m1_31_19_r;
wire signed [`CalcTempBus]          temp_m1_31_19_i;
wire signed [`CalcTempBus]          temp_m1_31_20_r;
wire signed [`CalcTempBus]          temp_m1_31_20_i;
wire signed [`CalcTempBus]          temp_m1_31_21_r;
wire signed [`CalcTempBus]          temp_m1_31_21_i;
wire signed [`CalcTempBus]          temp_m1_31_22_r;
wire signed [`CalcTempBus]          temp_m1_31_22_i;
wire signed [`CalcTempBus]          temp_m1_31_23_r;
wire signed [`CalcTempBus]          temp_m1_31_23_i;
wire signed [`CalcTempBus]          temp_m1_31_24_r;
wire signed [`CalcTempBus]          temp_m1_31_24_i;
wire signed [`CalcTempBus]          temp_m1_31_25_r;
wire signed [`CalcTempBus]          temp_m1_31_25_i;
wire signed [`CalcTempBus]          temp_m1_31_26_r;
wire signed [`CalcTempBus]          temp_m1_31_26_i;
wire signed [`CalcTempBus]          temp_m1_31_27_r;
wire signed [`CalcTempBus]          temp_m1_31_27_i;
wire signed [`CalcTempBus]          temp_m1_31_28_r;
wire signed [`CalcTempBus]          temp_m1_31_28_i;
wire signed [`CalcTempBus]          temp_m1_31_29_r;
wire signed [`CalcTempBus]          temp_m1_31_29_i;
wire signed [`CalcTempBus]          temp_m1_31_30_r;
wire signed [`CalcTempBus]          temp_m1_31_30_i;
wire signed [`CalcTempBus]          temp_m1_31_31_r;
wire signed [`CalcTempBus]          temp_m1_31_31_i;
wire signed [`CalcTempBus]          temp_m1_31_32_r;
wire signed [`CalcTempBus]          temp_m1_31_32_i;
wire signed [`CalcTempBus]          temp_m1_32_1_r;
wire signed [`CalcTempBus]          temp_m1_32_1_i;
wire signed [`CalcTempBus]          temp_m1_32_2_r;
wire signed [`CalcTempBus]          temp_m1_32_2_i;
wire signed [`CalcTempBus]          temp_m1_32_3_r;
wire signed [`CalcTempBus]          temp_m1_32_3_i;
wire signed [`CalcTempBus]          temp_m1_32_4_r;
wire signed [`CalcTempBus]          temp_m1_32_4_i;
wire signed [`CalcTempBus]          temp_m1_32_5_r;
wire signed [`CalcTempBus]          temp_m1_32_5_i;
wire signed [`CalcTempBus]          temp_m1_32_6_r;
wire signed [`CalcTempBus]          temp_m1_32_6_i;
wire signed [`CalcTempBus]          temp_m1_32_7_r;
wire signed [`CalcTempBus]          temp_m1_32_7_i;
wire signed [`CalcTempBus]          temp_m1_32_8_r;
wire signed [`CalcTempBus]          temp_m1_32_8_i;
wire signed [`CalcTempBus]          temp_m1_32_9_r;
wire signed [`CalcTempBus]          temp_m1_32_9_i;
wire signed [`CalcTempBus]          temp_m1_32_10_r;
wire signed [`CalcTempBus]          temp_m1_32_10_i;
wire signed [`CalcTempBus]          temp_m1_32_11_r;
wire signed [`CalcTempBus]          temp_m1_32_11_i;
wire signed [`CalcTempBus]          temp_m1_32_12_r;
wire signed [`CalcTempBus]          temp_m1_32_12_i;
wire signed [`CalcTempBus]          temp_m1_32_13_r;
wire signed [`CalcTempBus]          temp_m1_32_13_i;
wire signed [`CalcTempBus]          temp_m1_32_14_r;
wire signed [`CalcTempBus]          temp_m1_32_14_i;
wire signed [`CalcTempBus]          temp_m1_32_15_r;
wire signed [`CalcTempBus]          temp_m1_32_15_i;
wire signed [`CalcTempBus]          temp_m1_32_16_r;
wire signed [`CalcTempBus]          temp_m1_32_16_i;
wire signed [`CalcTempBus]          temp_m1_32_17_r;
wire signed [`CalcTempBus]          temp_m1_32_17_i;
wire signed [`CalcTempBus]          temp_m1_32_18_r;
wire signed [`CalcTempBus]          temp_m1_32_18_i;
wire signed [`CalcTempBus]          temp_m1_32_19_r;
wire signed [`CalcTempBus]          temp_m1_32_19_i;
wire signed [`CalcTempBus]          temp_m1_32_20_r;
wire signed [`CalcTempBus]          temp_m1_32_20_i;
wire signed [`CalcTempBus]          temp_m1_32_21_r;
wire signed [`CalcTempBus]          temp_m1_32_21_i;
wire signed [`CalcTempBus]          temp_m1_32_22_r;
wire signed [`CalcTempBus]          temp_m1_32_22_i;
wire signed [`CalcTempBus]          temp_m1_32_23_r;
wire signed [`CalcTempBus]          temp_m1_32_23_i;
wire signed [`CalcTempBus]          temp_m1_32_24_r;
wire signed [`CalcTempBus]          temp_m1_32_24_i;
wire signed [`CalcTempBus]          temp_m1_32_25_r;
wire signed [`CalcTempBus]          temp_m1_32_25_i;
wire signed [`CalcTempBus]          temp_m1_32_26_r;
wire signed [`CalcTempBus]          temp_m1_32_26_i;
wire signed [`CalcTempBus]          temp_m1_32_27_r;
wire signed [`CalcTempBus]          temp_m1_32_27_i;
wire signed [`CalcTempBus]          temp_m1_32_28_r;
wire signed [`CalcTempBus]          temp_m1_32_28_i;
wire signed [`CalcTempBus]          temp_m1_32_29_r;
wire signed [`CalcTempBus]          temp_m1_32_29_i;
wire signed [`CalcTempBus]          temp_m1_32_30_r;
wire signed [`CalcTempBus]          temp_m1_32_30_i;
wire signed [`CalcTempBus]          temp_m1_32_31_r;
wire signed [`CalcTempBus]          temp_m1_32_31_i;
wire signed [`CalcTempBus]          temp_m1_32_32_r;
wire signed [`CalcTempBus]          temp_m1_32_32_i;
wire signed [`CalcTempBus]          temp_m2_1_1_r;
wire signed [`CalcTempBus]          temp_m2_1_1_i;
wire signed [`CalcTempBus]          temp_m2_1_2_r;
wire signed [`CalcTempBus]          temp_m2_1_2_i;
wire signed [`CalcTempBus]          temp_m2_1_3_r;
wire signed [`CalcTempBus]          temp_m2_1_3_i;
wire signed [`CalcTempBus]          temp_m2_1_4_r;
wire signed [`CalcTempBus]          temp_m2_1_4_i;
wire signed [`CalcTempBus]          temp_m2_1_5_r;
wire signed [`CalcTempBus]          temp_m2_1_5_i;
wire signed [`CalcTempBus]          temp_m2_1_6_r;
wire signed [`CalcTempBus]          temp_m2_1_6_i;
wire signed [`CalcTempBus]          temp_m2_1_7_r;
wire signed [`CalcTempBus]          temp_m2_1_7_i;
wire signed [`CalcTempBus]          temp_m2_1_8_r;
wire signed [`CalcTempBus]          temp_m2_1_8_i;
wire signed [`CalcTempBus]          temp_m2_1_9_r;
wire signed [`CalcTempBus]          temp_m2_1_9_i;
wire signed [`CalcTempBus]          temp_m2_1_10_r;
wire signed [`CalcTempBus]          temp_m2_1_10_i;
wire signed [`CalcTempBus]          temp_m2_1_11_r;
wire signed [`CalcTempBus]          temp_m2_1_11_i;
wire signed [`CalcTempBus]          temp_m2_1_12_r;
wire signed [`CalcTempBus]          temp_m2_1_12_i;
wire signed [`CalcTempBus]          temp_m2_1_13_r;
wire signed [`CalcTempBus]          temp_m2_1_13_i;
wire signed [`CalcTempBus]          temp_m2_1_14_r;
wire signed [`CalcTempBus]          temp_m2_1_14_i;
wire signed [`CalcTempBus]          temp_m2_1_15_r;
wire signed [`CalcTempBus]          temp_m2_1_15_i;
wire signed [`CalcTempBus]          temp_m2_1_16_r;
wire signed [`CalcTempBus]          temp_m2_1_16_i;
wire signed [`CalcTempBus]          temp_m2_1_17_r;
wire signed [`CalcTempBus]          temp_m2_1_17_i;
wire signed [`CalcTempBus]          temp_m2_1_18_r;
wire signed [`CalcTempBus]          temp_m2_1_18_i;
wire signed [`CalcTempBus]          temp_m2_1_19_r;
wire signed [`CalcTempBus]          temp_m2_1_19_i;
wire signed [`CalcTempBus]          temp_m2_1_20_r;
wire signed [`CalcTempBus]          temp_m2_1_20_i;
wire signed [`CalcTempBus]          temp_m2_1_21_r;
wire signed [`CalcTempBus]          temp_m2_1_21_i;
wire signed [`CalcTempBus]          temp_m2_1_22_r;
wire signed [`CalcTempBus]          temp_m2_1_22_i;
wire signed [`CalcTempBus]          temp_m2_1_23_r;
wire signed [`CalcTempBus]          temp_m2_1_23_i;
wire signed [`CalcTempBus]          temp_m2_1_24_r;
wire signed [`CalcTempBus]          temp_m2_1_24_i;
wire signed [`CalcTempBus]          temp_m2_1_25_r;
wire signed [`CalcTempBus]          temp_m2_1_25_i;
wire signed [`CalcTempBus]          temp_m2_1_26_r;
wire signed [`CalcTempBus]          temp_m2_1_26_i;
wire signed [`CalcTempBus]          temp_m2_1_27_r;
wire signed [`CalcTempBus]          temp_m2_1_27_i;
wire signed [`CalcTempBus]          temp_m2_1_28_r;
wire signed [`CalcTempBus]          temp_m2_1_28_i;
wire signed [`CalcTempBus]          temp_m2_1_29_r;
wire signed [`CalcTempBus]          temp_m2_1_29_i;
wire signed [`CalcTempBus]          temp_m2_1_30_r;
wire signed [`CalcTempBus]          temp_m2_1_30_i;
wire signed [`CalcTempBus]          temp_m2_1_31_r;
wire signed [`CalcTempBus]          temp_m2_1_31_i;
wire signed [`CalcTempBus]          temp_m2_1_32_r;
wire signed [`CalcTempBus]          temp_m2_1_32_i;
wire signed [`CalcTempBus]          temp_m2_2_1_r;
wire signed [`CalcTempBus]          temp_m2_2_1_i;
wire signed [`CalcTempBus]          temp_m2_2_2_r;
wire signed [`CalcTempBus]          temp_m2_2_2_i;
wire signed [`CalcTempBus]          temp_m2_2_3_r;
wire signed [`CalcTempBus]          temp_m2_2_3_i;
wire signed [`CalcTempBus]          temp_m2_2_4_r;
wire signed [`CalcTempBus]          temp_m2_2_4_i;
wire signed [`CalcTempBus]          temp_m2_2_5_r;
wire signed [`CalcTempBus]          temp_m2_2_5_i;
wire signed [`CalcTempBus]          temp_m2_2_6_r;
wire signed [`CalcTempBus]          temp_m2_2_6_i;
wire signed [`CalcTempBus]          temp_m2_2_7_r;
wire signed [`CalcTempBus]          temp_m2_2_7_i;
wire signed [`CalcTempBus]          temp_m2_2_8_r;
wire signed [`CalcTempBus]          temp_m2_2_8_i;
wire signed [`CalcTempBus]          temp_m2_2_9_r;
wire signed [`CalcTempBus]          temp_m2_2_9_i;
wire signed [`CalcTempBus]          temp_m2_2_10_r;
wire signed [`CalcTempBus]          temp_m2_2_10_i;
wire signed [`CalcTempBus]          temp_m2_2_11_r;
wire signed [`CalcTempBus]          temp_m2_2_11_i;
wire signed [`CalcTempBus]          temp_m2_2_12_r;
wire signed [`CalcTempBus]          temp_m2_2_12_i;
wire signed [`CalcTempBus]          temp_m2_2_13_r;
wire signed [`CalcTempBus]          temp_m2_2_13_i;
wire signed [`CalcTempBus]          temp_m2_2_14_r;
wire signed [`CalcTempBus]          temp_m2_2_14_i;
wire signed [`CalcTempBus]          temp_m2_2_15_r;
wire signed [`CalcTempBus]          temp_m2_2_15_i;
wire signed [`CalcTempBus]          temp_m2_2_16_r;
wire signed [`CalcTempBus]          temp_m2_2_16_i;
wire signed [`CalcTempBus]          temp_m2_2_17_r;
wire signed [`CalcTempBus]          temp_m2_2_17_i;
wire signed [`CalcTempBus]          temp_m2_2_18_r;
wire signed [`CalcTempBus]          temp_m2_2_18_i;
wire signed [`CalcTempBus]          temp_m2_2_19_r;
wire signed [`CalcTempBus]          temp_m2_2_19_i;
wire signed [`CalcTempBus]          temp_m2_2_20_r;
wire signed [`CalcTempBus]          temp_m2_2_20_i;
wire signed [`CalcTempBus]          temp_m2_2_21_r;
wire signed [`CalcTempBus]          temp_m2_2_21_i;
wire signed [`CalcTempBus]          temp_m2_2_22_r;
wire signed [`CalcTempBus]          temp_m2_2_22_i;
wire signed [`CalcTempBus]          temp_m2_2_23_r;
wire signed [`CalcTempBus]          temp_m2_2_23_i;
wire signed [`CalcTempBus]          temp_m2_2_24_r;
wire signed [`CalcTempBus]          temp_m2_2_24_i;
wire signed [`CalcTempBus]          temp_m2_2_25_r;
wire signed [`CalcTempBus]          temp_m2_2_25_i;
wire signed [`CalcTempBus]          temp_m2_2_26_r;
wire signed [`CalcTempBus]          temp_m2_2_26_i;
wire signed [`CalcTempBus]          temp_m2_2_27_r;
wire signed [`CalcTempBus]          temp_m2_2_27_i;
wire signed [`CalcTempBus]          temp_m2_2_28_r;
wire signed [`CalcTempBus]          temp_m2_2_28_i;
wire signed [`CalcTempBus]          temp_m2_2_29_r;
wire signed [`CalcTempBus]          temp_m2_2_29_i;
wire signed [`CalcTempBus]          temp_m2_2_30_r;
wire signed [`CalcTempBus]          temp_m2_2_30_i;
wire signed [`CalcTempBus]          temp_m2_2_31_r;
wire signed [`CalcTempBus]          temp_m2_2_31_i;
wire signed [`CalcTempBus]          temp_m2_2_32_r;
wire signed [`CalcTempBus]          temp_m2_2_32_i;
wire signed [`CalcTempBus]          temp_m2_3_1_r;
wire signed [`CalcTempBus]          temp_m2_3_1_i;
wire signed [`CalcTempBus]          temp_m2_3_2_r;
wire signed [`CalcTempBus]          temp_m2_3_2_i;
wire signed [`CalcTempBus]          temp_m2_3_3_r;
wire signed [`CalcTempBus]          temp_m2_3_3_i;
wire signed [`CalcTempBus]          temp_m2_3_4_r;
wire signed [`CalcTempBus]          temp_m2_3_4_i;
wire signed [`CalcTempBus]          temp_m2_3_5_r;
wire signed [`CalcTempBus]          temp_m2_3_5_i;
wire signed [`CalcTempBus]          temp_m2_3_6_r;
wire signed [`CalcTempBus]          temp_m2_3_6_i;
wire signed [`CalcTempBus]          temp_m2_3_7_r;
wire signed [`CalcTempBus]          temp_m2_3_7_i;
wire signed [`CalcTempBus]          temp_m2_3_8_r;
wire signed [`CalcTempBus]          temp_m2_3_8_i;
wire signed [`CalcTempBus]          temp_m2_3_9_r;
wire signed [`CalcTempBus]          temp_m2_3_9_i;
wire signed [`CalcTempBus]          temp_m2_3_10_r;
wire signed [`CalcTempBus]          temp_m2_3_10_i;
wire signed [`CalcTempBus]          temp_m2_3_11_r;
wire signed [`CalcTempBus]          temp_m2_3_11_i;
wire signed [`CalcTempBus]          temp_m2_3_12_r;
wire signed [`CalcTempBus]          temp_m2_3_12_i;
wire signed [`CalcTempBus]          temp_m2_3_13_r;
wire signed [`CalcTempBus]          temp_m2_3_13_i;
wire signed [`CalcTempBus]          temp_m2_3_14_r;
wire signed [`CalcTempBus]          temp_m2_3_14_i;
wire signed [`CalcTempBus]          temp_m2_3_15_r;
wire signed [`CalcTempBus]          temp_m2_3_15_i;
wire signed [`CalcTempBus]          temp_m2_3_16_r;
wire signed [`CalcTempBus]          temp_m2_3_16_i;
wire signed [`CalcTempBus]          temp_m2_3_17_r;
wire signed [`CalcTempBus]          temp_m2_3_17_i;
wire signed [`CalcTempBus]          temp_m2_3_18_r;
wire signed [`CalcTempBus]          temp_m2_3_18_i;
wire signed [`CalcTempBus]          temp_m2_3_19_r;
wire signed [`CalcTempBus]          temp_m2_3_19_i;
wire signed [`CalcTempBus]          temp_m2_3_20_r;
wire signed [`CalcTempBus]          temp_m2_3_20_i;
wire signed [`CalcTempBus]          temp_m2_3_21_r;
wire signed [`CalcTempBus]          temp_m2_3_21_i;
wire signed [`CalcTempBus]          temp_m2_3_22_r;
wire signed [`CalcTempBus]          temp_m2_3_22_i;
wire signed [`CalcTempBus]          temp_m2_3_23_r;
wire signed [`CalcTempBus]          temp_m2_3_23_i;
wire signed [`CalcTempBus]          temp_m2_3_24_r;
wire signed [`CalcTempBus]          temp_m2_3_24_i;
wire signed [`CalcTempBus]          temp_m2_3_25_r;
wire signed [`CalcTempBus]          temp_m2_3_25_i;
wire signed [`CalcTempBus]          temp_m2_3_26_r;
wire signed [`CalcTempBus]          temp_m2_3_26_i;
wire signed [`CalcTempBus]          temp_m2_3_27_r;
wire signed [`CalcTempBus]          temp_m2_3_27_i;
wire signed [`CalcTempBus]          temp_m2_3_28_r;
wire signed [`CalcTempBus]          temp_m2_3_28_i;
wire signed [`CalcTempBus]          temp_m2_3_29_r;
wire signed [`CalcTempBus]          temp_m2_3_29_i;
wire signed [`CalcTempBus]          temp_m2_3_30_r;
wire signed [`CalcTempBus]          temp_m2_3_30_i;
wire signed [`CalcTempBus]          temp_m2_3_31_r;
wire signed [`CalcTempBus]          temp_m2_3_31_i;
wire signed [`CalcTempBus]          temp_m2_3_32_r;
wire signed [`CalcTempBus]          temp_m2_3_32_i;
wire signed [`CalcTempBus]          temp_m2_4_1_r;
wire signed [`CalcTempBus]          temp_m2_4_1_i;
wire signed [`CalcTempBus]          temp_m2_4_2_r;
wire signed [`CalcTempBus]          temp_m2_4_2_i;
wire signed [`CalcTempBus]          temp_m2_4_3_r;
wire signed [`CalcTempBus]          temp_m2_4_3_i;
wire signed [`CalcTempBus]          temp_m2_4_4_r;
wire signed [`CalcTempBus]          temp_m2_4_4_i;
wire signed [`CalcTempBus]          temp_m2_4_5_r;
wire signed [`CalcTempBus]          temp_m2_4_5_i;
wire signed [`CalcTempBus]          temp_m2_4_6_r;
wire signed [`CalcTempBus]          temp_m2_4_6_i;
wire signed [`CalcTempBus]          temp_m2_4_7_r;
wire signed [`CalcTempBus]          temp_m2_4_7_i;
wire signed [`CalcTempBus]          temp_m2_4_8_r;
wire signed [`CalcTempBus]          temp_m2_4_8_i;
wire signed [`CalcTempBus]          temp_m2_4_9_r;
wire signed [`CalcTempBus]          temp_m2_4_9_i;
wire signed [`CalcTempBus]          temp_m2_4_10_r;
wire signed [`CalcTempBus]          temp_m2_4_10_i;
wire signed [`CalcTempBus]          temp_m2_4_11_r;
wire signed [`CalcTempBus]          temp_m2_4_11_i;
wire signed [`CalcTempBus]          temp_m2_4_12_r;
wire signed [`CalcTempBus]          temp_m2_4_12_i;
wire signed [`CalcTempBus]          temp_m2_4_13_r;
wire signed [`CalcTempBus]          temp_m2_4_13_i;
wire signed [`CalcTempBus]          temp_m2_4_14_r;
wire signed [`CalcTempBus]          temp_m2_4_14_i;
wire signed [`CalcTempBus]          temp_m2_4_15_r;
wire signed [`CalcTempBus]          temp_m2_4_15_i;
wire signed [`CalcTempBus]          temp_m2_4_16_r;
wire signed [`CalcTempBus]          temp_m2_4_16_i;
wire signed [`CalcTempBus]          temp_m2_4_17_r;
wire signed [`CalcTempBus]          temp_m2_4_17_i;
wire signed [`CalcTempBus]          temp_m2_4_18_r;
wire signed [`CalcTempBus]          temp_m2_4_18_i;
wire signed [`CalcTempBus]          temp_m2_4_19_r;
wire signed [`CalcTempBus]          temp_m2_4_19_i;
wire signed [`CalcTempBus]          temp_m2_4_20_r;
wire signed [`CalcTempBus]          temp_m2_4_20_i;
wire signed [`CalcTempBus]          temp_m2_4_21_r;
wire signed [`CalcTempBus]          temp_m2_4_21_i;
wire signed [`CalcTempBus]          temp_m2_4_22_r;
wire signed [`CalcTempBus]          temp_m2_4_22_i;
wire signed [`CalcTempBus]          temp_m2_4_23_r;
wire signed [`CalcTempBus]          temp_m2_4_23_i;
wire signed [`CalcTempBus]          temp_m2_4_24_r;
wire signed [`CalcTempBus]          temp_m2_4_24_i;
wire signed [`CalcTempBus]          temp_m2_4_25_r;
wire signed [`CalcTempBus]          temp_m2_4_25_i;
wire signed [`CalcTempBus]          temp_m2_4_26_r;
wire signed [`CalcTempBus]          temp_m2_4_26_i;
wire signed [`CalcTempBus]          temp_m2_4_27_r;
wire signed [`CalcTempBus]          temp_m2_4_27_i;
wire signed [`CalcTempBus]          temp_m2_4_28_r;
wire signed [`CalcTempBus]          temp_m2_4_28_i;
wire signed [`CalcTempBus]          temp_m2_4_29_r;
wire signed [`CalcTempBus]          temp_m2_4_29_i;
wire signed [`CalcTempBus]          temp_m2_4_30_r;
wire signed [`CalcTempBus]          temp_m2_4_30_i;
wire signed [`CalcTempBus]          temp_m2_4_31_r;
wire signed [`CalcTempBus]          temp_m2_4_31_i;
wire signed [`CalcTempBus]          temp_m2_4_32_r;
wire signed [`CalcTempBus]          temp_m2_4_32_i;
wire signed [`CalcTempBus]          temp_m2_5_1_r;
wire signed [`CalcTempBus]          temp_m2_5_1_i;
wire signed [`CalcTempBus]          temp_m2_5_2_r;
wire signed [`CalcTempBus]          temp_m2_5_2_i;
wire signed [`CalcTempBus]          temp_m2_5_3_r;
wire signed [`CalcTempBus]          temp_m2_5_3_i;
wire signed [`CalcTempBus]          temp_m2_5_4_r;
wire signed [`CalcTempBus]          temp_m2_5_4_i;
wire signed [`CalcTempBus]          temp_m2_5_5_r;
wire signed [`CalcTempBus]          temp_m2_5_5_i;
wire signed [`CalcTempBus]          temp_m2_5_6_r;
wire signed [`CalcTempBus]          temp_m2_5_6_i;
wire signed [`CalcTempBus]          temp_m2_5_7_r;
wire signed [`CalcTempBus]          temp_m2_5_7_i;
wire signed [`CalcTempBus]          temp_m2_5_8_r;
wire signed [`CalcTempBus]          temp_m2_5_8_i;
wire signed [`CalcTempBus]          temp_m2_5_9_r;
wire signed [`CalcTempBus]          temp_m2_5_9_i;
wire signed [`CalcTempBus]          temp_m2_5_10_r;
wire signed [`CalcTempBus]          temp_m2_5_10_i;
wire signed [`CalcTempBus]          temp_m2_5_11_r;
wire signed [`CalcTempBus]          temp_m2_5_11_i;
wire signed [`CalcTempBus]          temp_m2_5_12_r;
wire signed [`CalcTempBus]          temp_m2_5_12_i;
wire signed [`CalcTempBus]          temp_m2_5_13_r;
wire signed [`CalcTempBus]          temp_m2_5_13_i;
wire signed [`CalcTempBus]          temp_m2_5_14_r;
wire signed [`CalcTempBus]          temp_m2_5_14_i;
wire signed [`CalcTempBus]          temp_m2_5_15_r;
wire signed [`CalcTempBus]          temp_m2_5_15_i;
wire signed [`CalcTempBus]          temp_m2_5_16_r;
wire signed [`CalcTempBus]          temp_m2_5_16_i;
wire signed [`CalcTempBus]          temp_m2_5_17_r;
wire signed [`CalcTempBus]          temp_m2_5_17_i;
wire signed [`CalcTempBus]          temp_m2_5_18_r;
wire signed [`CalcTempBus]          temp_m2_5_18_i;
wire signed [`CalcTempBus]          temp_m2_5_19_r;
wire signed [`CalcTempBus]          temp_m2_5_19_i;
wire signed [`CalcTempBus]          temp_m2_5_20_r;
wire signed [`CalcTempBus]          temp_m2_5_20_i;
wire signed [`CalcTempBus]          temp_m2_5_21_r;
wire signed [`CalcTempBus]          temp_m2_5_21_i;
wire signed [`CalcTempBus]          temp_m2_5_22_r;
wire signed [`CalcTempBus]          temp_m2_5_22_i;
wire signed [`CalcTempBus]          temp_m2_5_23_r;
wire signed [`CalcTempBus]          temp_m2_5_23_i;
wire signed [`CalcTempBus]          temp_m2_5_24_r;
wire signed [`CalcTempBus]          temp_m2_5_24_i;
wire signed [`CalcTempBus]          temp_m2_5_25_r;
wire signed [`CalcTempBus]          temp_m2_5_25_i;
wire signed [`CalcTempBus]          temp_m2_5_26_r;
wire signed [`CalcTempBus]          temp_m2_5_26_i;
wire signed [`CalcTempBus]          temp_m2_5_27_r;
wire signed [`CalcTempBus]          temp_m2_5_27_i;
wire signed [`CalcTempBus]          temp_m2_5_28_r;
wire signed [`CalcTempBus]          temp_m2_5_28_i;
wire signed [`CalcTempBus]          temp_m2_5_29_r;
wire signed [`CalcTempBus]          temp_m2_5_29_i;
wire signed [`CalcTempBus]          temp_m2_5_30_r;
wire signed [`CalcTempBus]          temp_m2_5_30_i;
wire signed [`CalcTempBus]          temp_m2_5_31_r;
wire signed [`CalcTempBus]          temp_m2_5_31_i;
wire signed [`CalcTempBus]          temp_m2_5_32_r;
wire signed [`CalcTempBus]          temp_m2_5_32_i;
wire signed [`CalcTempBus]          temp_m2_6_1_r;
wire signed [`CalcTempBus]          temp_m2_6_1_i;
wire signed [`CalcTempBus]          temp_m2_6_2_r;
wire signed [`CalcTempBus]          temp_m2_6_2_i;
wire signed [`CalcTempBus]          temp_m2_6_3_r;
wire signed [`CalcTempBus]          temp_m2_6_3_i;
wire signed [`CalcTempBus]          temp_m2_6_4_r;
wire signed [`CalcTempBus]          temp_m2_6_4_i;
wire signed [`CalcTempBus]          temp_m2_6_5_r;
wire signed [`CalcTempBus]          temp_m2_6_5_i;
wire signed [`CalcTempBus]          temp_m2_6_6_r;
wire signed [`CalcTempBus]          temp_m2_6_6_i;
wire signed [`CalcTempBus]          temp_m2_6_7_r;
wire signed [`CalcTempBus]          temp_m2_6_7_i;
wire signed [`CalcTempBus]          temp_m2_6_8_r;
wire signed [`CalcTempBus]          temp_m2_6_8_i;
wire signed [`CalcTempBus]          temp_m2_6_9_r;
wire signed [`CalcTempBus]          temp_m2_6_9_i;
wire signed [`CalcTempBus]          temp_m2_6_10_r;
wire signed [`CalcTempBus]          temp_m2_6_10_i;
wire signed [`CalcTempBus]          temp_m2_6_11_r;
wire signed [`CalcTempBus]          temp_m2_6_11_i;
wire signed [`CalcTempBus]          temp_m2_6_12_r;
wire signed [`CalcTempBus]          temp_m2_6_12_i;
wire signed [`CalcTempBus]          temp_m2_6_13_r;
wire signed [`CalcTempBus]          temp_m2_6_13_i;
wire signed [`CalcTempBus]          temp_m2_6_14_r;
wire signed [`CalcTempBus]          temp_m2_6_14_i;
wire signed [`CalcTempBus]          temp_m2_6_15_r;
wire signed [`CalcTempBus]          temp_m2_6_15_i;
wire signed [`CalcTempBus]          temp_m2_6_16_r;
wire signed [`CalcTempBus]          temp_m2_6_16_i;
wire signed [`CalcTempBus]          temp_m2_6_17_r;
wire signed [`CalcTempBus]          temp_m2_6_17_i;
wire signed [`CalcTempBus]          temp_m2_6_18_r;
wire signed [`CalcTempBus]          temp_m2_6_18_i;
wire signed [`CalcTempBus]          temp_m2_6_19_r;
wire signed [`CalcTempBus]          temp_m2_6_19_i;
wire signed [`CalcTempBus]          temp_m2_6_20_r;
wire signed [`CalcTempBus]          temp_m2_6_20_i;
wire signed [`CalcTempBus]          temp_m2_6_21_r;
wire signed [`CalcTempBus]          temp_m2_6_21_i;
wire signed [`CalcTempBus]          temp_m2_6_22_r;
wire signed [`CalcTempBus]          temp_m2_6_22_i;
wire signed [`CalcTempBus]          temp_m2_6_23_r;
wire signed [`CalcTempBus]          temp_m2_6_23_i;
wire signed [`CalcTempBus]          temp_m2_6_24_r;
wire signed [`CalcTempBus]          temp_m2_6_24_i;
wire signed [`CalcTempBus]          temp_m2_6_25_r;
wire signed [`CalcTempBus]          temp_m2_6_25_i;
wire signed [`CalcTempBus]          temp_m2_6_26_r;
wire signed [`CalcTempBus]          temp_m2_6_26_i;
wire signed [`CalcTempBus]          temp_m2_6_27_r;
wire signed [`CalcTempBus]          temp_m2_6_27_i;
wire signed [`CalcTempBus]          temp_m2_6_28_r;
wire signed [`CalcTempBus]          temp_m2_6_28_i;
wire signed [`CalcTempBus]          temp_m2_6_29_r;
wire signed [`CalcTempBus]          temp_m2_6_29_i;
wire signed [`CalcTempBus]          temp_m2_6_30_r;
wire signed [`CalcTempBus]          temp_m2_6_30_i;
wire signed [`CalcTempBus]          temp_m2_6_31_r;
wire signed [`CalcTempBus]          temp_m2_6_31_i;
wire signed [`CalcTempBus]          temp_m2_6_32_r;
wire signed [`CalcTempBus]          temp_m2_6_32_i;
wire signed [`CalcTempBus]          temp_m2_7_1_r;
wire signed [`CalcTempBus]          temp_m2_7_1_i;
wire signed [`CalcTempBus]          temp_m2_7_2_r;
wire signed [`CalcTempBus]          temp_m2_7_2_i;
wire signed [`CalcTempBus]          temp_m2_7_3_r;
wire signed [`CalcTempBus]          temp_m2_7_3_i;
wire signed [`CalcTempBus]          temp_m2_7_4_r;
wire signed [`CalcTempBus]          temp_m2_7_4_i;
wire signed [`CalcTempBus]          temp_m2_7_5_r;
wire signed [`CalcTempBus]          temp_m2_7_5_i;
wire signed [`CalcTempBus]          temp_m2_7_6_r;
wire signed [`CalcTempBus]          temp_m2_7_6_i;
wire signed [`CalcTempBus]          temp_m2_7_7_r;
wire signed [`CalcTempBus]          temp_m2_7_7_i;
wire signed [`CalcTempBus]          temp_m2_7_8_r;
wire signed [`CalcTempBus]          temp_m2_7_8_i;
wire signed [`CalcTempBus]          temp_m2_7_9_r;
wire signed [`CalcTempBus]          temp_m2_7_9_i;
wire signed [`CalcTempBus]          temp_m2_7_10_r;
wire signed [`CalcTempBus]          temp_m2_7_10_i;
wire signed [`CalcTempBus]          temp_m2_7_11_r;
wire signed [`CalcTempBus]          temp_m2_7_11_i;
wire signed [`CalcTempBus]          temp_m2_7_12_r;
wire signed [`CalcTempBus]          temp_m2_7_12_i;
wire signed [`CalcTempBus]          temp_m2_7_13_r;
wire signed [`CalcTempBus]          temp_m2_7_13_i;
wire signed [`CalcTempBus]          temp_m2_7_14_r;
wire signed [`CalcTempBus]          temp_m2_7_14_i;
wire signed [`CalcTempBus]          temp_m2_7_15_r;
wire signed [`CalcTempBus]          temp_m2_7_15_i;
wire signed [`CalcTempBus]          temp_m2_7_16_r;
wire signed [`CalcTempBus]          temp_m2_7_16_i;
wire signed [`CalcTempBus]          temp_m2_7_17_r;
wire signed [`CalcTempBus]          temp_m2_7_17_i;
wire signed [`CalcTempBus]          temp_m2_7_18_r;
wire signed [`CalcTempBus]          temp_m2_7_18_i;
wire signed [`CalcTempBus]          temp_m2_7_19_r;
wire signed [`CalcTempBus]          temp_m2_7_19_i;
wire signed [`CalcTempBus]          temp_m2_7_20_r;
wire signed [`CalcTempBus]          temp_m2_7_20_i;
wire signed [`CalcTempBus]          temp_m2_7_21_r;
wire signed [`CalcTempBus]          temp_m2_7_21_i;
wire signed [`CalcTempBus]          temp_m2_7_22_r;
wire signed [`CalcTempBus]          temp_m2_7_22_i;
wire signed [`CalcTempBus]          temp_m2_7_23_r;
wire signed [`CalcTempBus]          temp_m2_7_23_i;
wire signed [`CalcTempBus]          temp_m2_7_24_r;
wire signed [`CalcTempBus]          temp_m2_7_24_i;
wire signed [`CalcTempBus]          temp_m2_7_25_r;
wire signed [`CalcTempBus]          temp_m2_7_25_i;
wire signed [`CalcTempBus]          temp_m2_7_26_r;
wire signed [`CalcTempBus]          temp_m2_7_26_i;
wire signed [`CalcTempBus]          temp_m2_7_27_r;
wire signed [`CalcTempBus]          temp_m2_7_27_i;
wire signed [`CalcTempBus]          temp_m2_7_28_r;
wire signed [`CalcTempBus]          temp_m2_7_28_i;
wire signed [`CalcTempBus]          temp_m2_7_29_r;
wire signed [`CalcTempBus]          temp_m2_7_29_i;
wire signed [`CalcTempBus]          temp_m2_7_30_r;
wire signed [`CalcTempBus]          temp_m2_7_30_i;
wire signed [`CalcTempBus]          temp_m2_7_31_r;
wire signed [`CalcTempBus]          temp_m2_7_31_i;
wire signed [`CalcTempBus]          temp_m2_7_32_r;
wire signed [`CalcTempBus]          temp_m2_7_32_i;
wire signed [`CalcTempBus]          temp_m2_8_1_r;
wire signed [`CalcTempBus]          temp_m2_8_1_i;
wire signed [`CalcTempBus]          temp_m2_8_2_r;
wire signed [`CalcTempBus]          temp_m2_8_2_i;
wire signed [`CalcTempBus]          temp_m2_8_3_r;
wire signed [`CalcTempBus]          temp_m2_8_3_i;
wire signed [`CalcTempBus]          temp_m2_8_4_r;
wire signed [`CalcTempBus]          temp_m2_8_4_i;
wire signed [`CalcTempBus]          temp_m2_8_5_r;
wire signed [`CalcTempBus]          temp_m2_8_5_i;
wire signed [`CalcTempBus]          temp_m2_8_6_r;
wire signed [`CalcTempBus]          temp_m2_8_6_i;
wire signed [`CalcTempBus]          temp_m2_8_7_r;
wire signed [`CalcTempBus]          temp_m2_8_7_i;
wire signed [`CalcTempBus]          temp_m2_8_8_r;
wire signed [`CalcTempBus]          temp_m2_8_8_i;
wire signed [`CalcTempBus]          temp_m2_8_9_r;
wire signed [`CalcTempBus]          temp_m2_8_9_i;
wire signed [`CalcTempBus]          temp_m2_8_10_r;
wire signed [`CalcTempBus]          temp_m2_8_10_i;
wire signed [`CalcTempBus]          temp_m2_8_11_r;
wire signed [`CalcTempBus]          temp_m2_8_11_i;
wire signed [`CalcTempBus]          temp_m2_8_12_r;
wire signed [`CalcTempBus]          temp_m2_8_12_i;
wire signed [`CalcTempBus]          temp_m2_8_13_r;
wire signed [`CalcTempBus]          temp_m2_8_13_i;
wire signed [`CalcTempBus]          temp_m2_8_14_r;
wire signed [`CalcTempBus]          temp_m2_8_14_i;
wire signed [`CalcTempBus]          temp_m2_8_15_r;
wire signed [`CalcTempBus]          temp_m2_8_15_i;
wire signed [`CalcTempBus]          temp_m2_8_16_r;
wire signed [`CalcTempBus]          temp_m2_8_16_i;
wire signed [`CalcTempBus]          temp_m2_8_17_r;
wire signed [`CalcTempBus]          temp_m2_8_17_i;
wire signed [`CalcTempBus]          temp_m2_8_18_r;
wire signed [`CalcTempBus]          temp_m2_8_18_i;
wire signed [`CalcTempBus]          temp_m2_8_19_r;
wire signed [`CalcTempBus]          temp_m2_8_19_i;
wire signed [`CalcTempBus]          temp_m2_8_20_r;
wire signed [`CalcTempBus]          temp_m2_8_20_i;
wire signed [`CalcTempBus]          temp_m2_8_21_r;
wire signed [`CalcTempBus]          temp_m2_8_21_i;
wire signed [`CalcTempBus]          temp_m2_8_22_r;
wire signed [`CalcTempBus]          temp_m2_8_22_i;
wire signed [`CalcTempBus]          temp_m2_8_23_r;
wire signed [`CalcTempBus]          temp_m2_8_23_i;
wire signed [`CalcTempBus]          temp_m2_8_24_r;
wire signed [`CalcTempBus]          temp_m2_8_24_i;
wire signed [`CalcTempBus]          temp_m2_8_25_r;
wire signed [`CalcTempBus]          temp_m2_8_25_i;
wire signed [`CalcTempBus]          temp_m2_8_26_r;
wire signed [`CalcTempBus]          temp_m2_8_26_i;
wire signed [`CalcTempBus]          temp_m2_8_27_r;
wire signed [`CalcTempBus]          temp_m2_8_27_i;
wire signed [`CalcTempBus]          temp_m2_8_28_r;
wire signed [`CalcTempBus]          temp_m2_8_28_i;
wire signed [`CalcTempBus]          temp_m2_8_29_r;
wire signed [`CalcTempBus]          temp_m2_8_29_i;
wire signed [`CalcTempBus]          temp_m2_8_30_r;
wire signed [`CalcTempBus]          temp_m2_8_30_i;
wire signed [`CalcTempBus]          temp_m2_8_31_r;
wire signed [`CalcTempBus]          temp_m2_8_31_i;
wire signed [`CalcTempBus]          temp_m2_8_32_r;
wire signed [`CalcTempBus]          temp_m2_8_32_i;
wire signed [`CalcTempBus]          temp_m2_9_1_r;
wire signed [`CalcTempBus]          temp_m2_9_1_i;
wire signed [`CalcTempBus]          temp_m2_9_2_r;
wire signed [`CalcTempBus]          temp_m2_9_2_i;
wire signed [`CalcTempBus]          temp_m2_9_3_r;
wire signed [`CalcTempBus]          temp_m2_9_3_i;
wire signed [`CalcTempBus]          temp_m2_9_4_r;
wire signed [`CalcTempBus]          temp_m2_9_4_i;
wire signed [`CalcTempBus]          temp_m2_9_5_r;
wire signed [`CalcTempBus]          temp_m2_9_5_i;
wire signed [`CalcTempBus]          temp_m2_9_6_r;
wire signed [`CalcTempBus]          temp_m2_9_6_i;
wire signed [`CalcTempBus]          temp_m2_9_7_r;
wire signed [`CalcTempBus]          temp_m2_9_7_i;
wire signed [`CalcTempBus]          temp_m2_9_8_r;
wire signed [`CalcTempBus]          temp_m2_9_8_i;
wire signed [`CalcTempBus]          temp_m2_9_9_r;
wire signed [`CalcTempBus]          temp_m2_9_9_i;
wire signed [`CalcTempBus]          temp_m2_9_10_r;
wire signed [`CalcTempBus]          temp_m2_9_10_i;
wire signed [`CalcTempBus]          temp_m2_9_11_r;
wire signed [`CalcTempBus]          temp_m2_9_11_i;
wire signed [`CalcTempBus]          temp_m2_9_12_r;
wire signed [`CalcTempBus]          temp_m2_9_12_i;
wire signed [`CalcTempBus]          temp_m2_9_13_r;
wire signed [`CalcTempBus]          temp_m2_9_13_i;
wire signed [`CalcTempBus]          temp_m2_9_14_r;
wire signed [`CalcTempBus]          temp_m2_9_14_i;
wire signed [`CalcTempBus]          temp_m2_9_15_r;
wire signed [`CalcTempBus]          temp_m2_9_15_i;
wire signed [`CalcTempBus]          temp_m2_9_16_r;
wire signed [`CalcTempBus]          temp_m2_9_16_i;
wire signed [`CalcTempBus]          temp_m2_9_17_r;
wire signed [`CalcTempBus]          temp_m2_9_17_i;
wire signed [`CalcTempBus]          temp_m2_9_18_r;
wire signed [`CalcTempBus]          temp_m2_9_18_i;
wire signed [`CalcTempBus]          temp_m2_9_19_r;
wire signed [`CalcTempBus]          temp_m2_9_19_i;
wire signed [`CalcTempBus]          temp_m2_9_20_r;
wire signed [`CalcTempBus]          temp_m2_9_20_i;
wire signed [`CalcTempBus]          temp_m2_9_21_r;
wire signed [`CalcTempBus]          temp_m2_9_21_i;
wire signed [`CalcTempBus]          temp_m2_9_22_r;
wire signed [`CalcTempBus]          temp_m2_9_22_i;
wire signed [`CalcTempBus]          temp_m2_9_23_r;
wire signed [`CalcTempBus]          temp_m2_9_23_i;
wire signed [`CalcTempBus]          temp_m2_9_24_r;
wire signed [`CalcTempBus]          temp_m2_9_24_i;
wire signed [`CalcTempBus]          temp_m2_9_25_r;
wire signed [`CalcTempBus]          temp_m2_9_25_i;
wire signed [`CalcTempBus]          temp_m2_9_26_r;
wire signed [`CalcTempBus]          temp_m2_9_26_i;
wire signed [`CalcTempBus]          temp_m2_9_27_r;
wire signed [`CalcTempBus]          temp_m2_9_27_i;
wire signed [`CalcTempBus]          temp_m2_9_28_r;
wire signed [`CalcTempBus]          temp_m2_9_28_i;
wire signed [`CalcTempBus]          temp_m2_9_29_r;
wire signed [`CalcTempBus]          temp_m2_9_29_i;
wire signed [`CalcTempBus]          temp_m2_9_30_r;
wire signed [`CalcTempBus]          temp_m2_9_30_i;
wire signed [`CalcTempBus]          temp_m2_9_31_r;
wire signed [`CalcTempBus]          temp_m2_9_31_i;
wire signed [`CalcTempBus]          temp_m2_9_32_r;
wire signed [`CalcTempBus]          temp_m2_9_32_i;
wire signed [`CalcTempBus]          temp_m2_10_1_r;
wire signed [`CalcTempBus]          temp_m2_10_1_i;
wire signed [`CalcTempBus]          temp_m2_10_2_r;
wire signed [`CalcTempBus]          temp_m2_10_2_i;
wire signed [`CalcTempBus]          temp_m2_10_3_r;
wire signed [`CalcTempBus]          temp_m2_10_3_i;
wire signed [`CalcTempBus]          temp_m2_10_4_r;
wire signed [`CalcTempBus]          temp_m2_10_4_i;
wire signed [`CalcTempBus]          temp_m2_10_5_r;
wire signed [`CalcTempBus]          temp_m2_10_5_i;
wire signed [`CalcTempBus]          temp_m2_10_6_r;
wire signed [`CalcTempBus]          temp_m2_10_6_i;
wire signed [`CalcTempBus]          temp_m2_10_7_r;
wire signed [`CalcTempBus]          temp_m2_10_7_i;
wire signed [`CalcTempBus]          temp_m2_10_8_r;
wire signed [`CalcTempBus]          temp_m2_10_8_i;
wire signed [`CalcTempBus]          temp_m2_10_9_r;
wire signed [`CalcTempBus]          temp_m2_10_9_i;
wire signed [`CalcTempBus]          temp_m2_10_10_r;
wire signed [`CalcTempBus]          temp_m2_10_10_i;
wire signed [`CalcTempBus]          temp_m2_10_11_r;
wire signed [`CalcTempBus]          temp_m2_10_11_i;
wire signed [`CalcTempBus]          temp_m2_10_12_r;
wire signed [`CalcTempBus]          temp_m2_10_12_i;
wire signed [`CalcTempBus]          temp_m2_10_13_r;
wire signed [`CalcTempBus]          temp_m2_10_13_i;
wire signed [`CalcTempBus]          temp_m2_10_14_r;
wire signed [`CalcTempBus]          temp_m2_10_14_i;
wire signed [`CalcTempBus]          temp_m2_10_15_r;
wire signed [`CalcTempBus]          temp_m2_10_15_i;
wire signed [`CalcTempBus]          temp_m2_10_16_r;
wire signed [`CalcTempBus]          temp_m2_10_16_i;
wire signed [`CalcTempBus]          temp_m2_10_17_r;
wire signed [`CalcTempBus]          temp_m2_10_17_i;
wire signed [`CalcTempBus]          temp_m2_10_18_r;
wire signed [`CalcTempBus]          temp_m2_10_18_i;
wire signed [`CalcTempBus]          temp_m2_10_19_r;
wire signed [`CalcTempBus]          temp_m2_10_19_i;
wire signed [`CalcTempBus]          temp_m2_10_20_r;
wire signed [`CalcTempBus]          temp_m2_10_20_i;
wire signed [`CalcTempBus]          temp_m2_10_21_r;
wire signed [`CalcTempBus]          temp_m2_10_21_i;
wire signed [`CalcTempBus]          temp_m2_10_22_r;
wire signed [`CalcTempBus]          temp_m2_10_22_i;
wire signed [`CalcTempBus]          temp_m2_10_23_r;
wire signed [`CalcTempBus]          temp_m2_10_23_i;
wire signed [`CalcTempBus]          temp_m2_10_24_r;
wire signed [`CalcTempBus]          temp_m2_10_24_i;
wire signed [`CalcTempBus]          temp_m2_10_25_r;
wire signed [`CalcTempBus]          temp_m2_10_25_i;
wire signed [`CalcTempBus]          temp_m2_10_26_r;
wire signed [`CalcTempBus]          temp_m2_10_26_i;
wire signed [`CalcTempBus]          temp_m2_10_27_r;
wire signed [`CalcTempBus]          temp_m2_10_27_i;
wire signed [`CalcTempBus]          temp_m2_10_28_r;
wire signed [`CalcTempBus]          temp_m2_10_28_i;
wire signed [`CalcTempBus]          temp_m2_10_29_r;
wire signed [`CalcTempBus]          temp_m2_10_29_i;
wire signed [`CalcTempBus]          temp_m2_10_30_r;
wire signed [`CalcTempBus]          temp_m2_10_30_i;
wire signed [`CalcTempBus]          temp_m2_10_31_r;
wire signed [`CalcTempBus]          temp_m2_10_31_i;
wire signed [`CalcTempBus]          temp_m2_10_32_r;
wire signed [`CalcTempBus]          temp_m2_10_32_i;
wire signed [`CalcTempBus]          temp_m2_11_1_r;
wire signed [`CalcTempBus]          temp_m2_11_1_i;
wire signed [`CalcTempBus]          temp_m2_11_2_r;
wire signed [`CalcTempBus]          temp_m2_11_2_i;
wire signed [`CalcTempBus]          temp_m2_11_3_r;
wire signed [`CalcTempBus]          temp_m2_11_3_i;
wire signed [`CalcTempBus]          temp_m2_11_4_r;
wire signed [`CalcTempBus]          temp_m2_11_4_i;
wire signed [`CalcTempBus]          temp_m2_11_5_r;
wire signed [`CalcTempBus]          temp_m2_11_5_i;
wire signed [`CalcTempBus]          temp_m2_11_6_r;
wire signed [`CalcTempBus]          temp_m2_11_6_i;
wire signed [`CalcTempBus]          temp_m2_11_7_r;
wire signed [`CalcTempBus]          temp_m2_11_7_i;
wire signed [`CalcTempBus]          temp_m2_11_8_r;
wire signed [`CalcTempBus]          temp_m2_11_8_i;
wire signed [`CalcTempBus]          temp_m2_11_9_r;
wire signed [`CalcTempBus]          temp_m2_11_9_i;
wire signed [`CalcTempBus]          temp_m2_11_10_r;
wire signed [`CalcTempBus]          temp_m2_11_10_i;
wire signed [`CalcTempBus]          temp_m2_11_11_r;
wire signed [`CalcTempBus]          temp_m2_11_11_i;
wire signed [`CalcTempBus]          temp_m2_11_12_r;
wire signed [`CalcTempBus]          temp_m2_11_12_i;
wire signed [`CalcTempBus]          temp_m2_11_13_r;
wire signed [`CalcTempBus]          temp_m2_11_13_i;
wire signed [`CalcTempBus]          temp_m2_11_14_r;
wire signed [`CalcTempBus]          temp_m2_11_14_i;
wire signed [`CalcTempBus]          temp_m2_11_15_r;
wire signed [`CalcTempBus]          temp_m2_11_15_i;
wire signed [`CalcTempBus]          temp_m2_11_16_r;
wire signed [`CalcTempBus]          temp_m2_11_16_i;
wire signed [`CalcTempBus]          temp_m2_11_17_r;
wire signed [`CalcTempBus]          temp_m2_11_17_i;
wire signed [`CalcTempBus]          temp_m2_11_18_r;
wire signed [`CalcTempBus]          temp_m2_11_18_i;
wire signed [`CalcTempBus]          temp_m2_11_19_r;
wire signed [`CalcTempBus]          temp_m2_11_19_i;
wire signed [`CalcTempBus]          temp_m2_11_20_r;
wire signed [`CalcTempBus]          temp_m2_11_20_i;
wire signed [`CalcTempBus]          temp_m2_11_21_r;
wire signed [`CalcTempBus]          temp_m2_11_21_i;
wire signed [`CalcTempBus]          temp_m2_11_22_r;
wire signed [`CalcTempBus]          temp_m2_11_22_i;
wire signed [`CalcTempBus]          temp_m2_11_23_r;
wire signed [`CalcTempBus]          temp_m2_11_23_i;
wire signed [`CalcTempBus]          temp_m2_11_24_r;
wire signed [`CalcTempBus]          temp_m2_11_24_i;
wire signed [`CalcTempBus]          temp_m2_11_25_r;
wire signed [`CalcTempBus]          temp_m2_11_25_i;
wire signed [`CalcTempBus]          temp_m2_11_26_r;
wire signed [`CalcTempBus]          temp_m2_11_26_i;
wire signed [`CalcTempBus]          temp_m2_11_27_r;
wire signed [`CalcTempBus]          temp_m2_11_27_i;
wire signed [`CalcTempBus]          temp_m2_11_28_r;
wire signed [`CalcTempBus]          temp_m2_11_28_i;
wire signed [`CalcTempBus]          temp_m2_11_29_r;
wire signed [`CalcTempBus]          temp_m2_11_29_i;
wire signed [`CalcTempBus]          temp_m2_11_30_r;
wire signed [`CalcTempBus]          temp_m2_11_30_i;
wire signed [`CalcTempBus]          temp_m2_11_31_r;
wire signed [`CalcTempBus]          temp_m2_11_31_i;
wire signed [`CalcTempBus]          temp_m2_11_32_r;
wire signed [`CalcTempBus]          temp_m2_11_32_i;
wire signed [`CalcTempBus]          temp_m2_12_1_r;
wire signed [`CalcTempBus]          temp_m2_12_1_i;
wire signed [`CalcTempBus]          temp_m2_12_2_r;
wire signed [`CalcTempBus]          temp_m2_12_2_i;
wire signed [`CalcTempBus]          temp_m2_12_3_r;
wire signed [`CalcTempBus]          temp_m2_12_3_i;
wire signed [`CalcTempBus]          temp_m2_12_4_r;
wire signed [`CalcTempBus]          temp_m2_12_4_i;
wire signed [`CalcTempBus]          temp_m2_12_5_r;
wire signed [`CalcTempBus]          temp_m2_12_5_i;
wire signed [`CalcTempBus]          temp_m2_12_6_r;
wire signed [`CalcTempBus]          temp_m2_12_6_i;
wire signed [`CalcTempBus]          temp_m2_12_7_r;
wire signed [`CalcTempBus]          temp_m2_12_7_i;
wire signed [`CalcTempBus]          temp_m2_12_8_r;
wire signed [`CalcTempBus]          temp_m2_12_8_i;
wire signed [`CalcTempBus]          temp_m2_12_9_r;
wire signed [`CalcTempBus]          temp_m2_12_9_i;
wire signed [`CalcTempBus]          temp_m2_12_10_r;
wire signed [`CalcTempBus]          temp_m2_12_10_i;
wire signed [`CalcTempBus]          temp_m2_12_11_r;
wire signed [`CalcTempBus]          temp_m2_12_11_i;
wire signed [`CalcTempBus]          temp_m2_12_12_r;
wire signed [`CalcTempBus]          temp_m2_12_12_i;
wire signed [`CalcTempBus]          temp_m2_12_13_r;
wire signed [`CalcTempBus]          temp_m2_12_13_i;
wire signed [`CalcTempBus]          temp_m2_12_14_r;
wire signed [`CalcTempBus]          temp_m2_12_14_i;
wire signed [`CalcTempBus]          temp_m2_12_15_r;
wire signed [`CalcTempBus]          temp_m2_12_15_i;
wire signed [`CalcTempBus]          temp_m2_12_16_r;
wire signed [`CalcTempBus]          temp_m2_12_16_i;
wire signed [`CalcTempBus]          temp_m2_12_17_r;
wire signed [`CalcTempBus]          temp_m2_12_17_i;
wire signed [`CalcTempBus]          temp_m2_12_18_r;
wire signed [`CalcTempBus]          temp_m2_12_18_i;
wire signed [`CalcTempBus]          temp_m2_12_19_r;
wire signed [`CalcTempBus]          temp_m2_12_19_i;
wire signed [`CalcTempBus]          temp_m2_12_20_r;
wire signed [`CalcTempBus]          temp_m2_12_20_i;
wire signed [`CalcTempBus]          temp_m2_12_21_r;
wire signed [`CalcTempBus]          temp_m2_12_21_i;
wire signed [`CalcTempBus]          temp_m2_12_22_r;
wire signed [`CalcTempBus]          temp_m2_12_22_i;
wire signed [`CalcTempBus]          temp_m2_12_23_r;
wire signed [`CalcTempBus]          temp_m2_12_23_i;
wire signed [`CalcTempBus]          temp_m2_12_24_r;
wire signed [`CalcTempBus]          temp_m2_12_24_i;
wire signed [`CalcTempBus]          temp_m2_12_25_r;
wire signed [`CalcTempBus]          temp_m2_12_25_i;
wire signed [`CalcTempBus]          temp_m2_12_26_r;
wire signed [`CalcTempBus]          temp_m2_12_26_i;
wire signed [`CalcTempBus]          temp_m2_12_27_r;
wire signed [`CalcTempBus]          temp_m2_12_27_i;
wire signed [`CalcTempBus]          temp_m2_12_28_r;
wire signed [`CalcTempBus]          temp_m2_12_28_i;
wire signed [`CalcTempBus]          temp_m2_12_29_r;
wire signed [`CalcTempBus]          temp_m2_12_29_i;
wire signed [`CalcTempBus]          temp_m2_12_30_r;
wire signed [`CalcTempBus]          temp_m2_12_30_i;
wire signed [`CalcTempBus]          temp_m2_12_31_r;
wire signed [`CalcTempBus]          temp_m2_12_31_i;
wire signed [`CalcTempBus]          temp_m2_12_32_r;
wire signed [`CalcTempBus]          temp_m2_12_32_i;
wire signed [`CalcTempBus]          temp_m2_13_1_r;
wire signed [`CalcTempBus]          temp_m2_13_1_i;
wire signed [`CalcTempBus]          temp_m2_13_2_r;
wire signed [`CalcTempBus]          temp_m2_13_2_i;
wire signed [`CalcTempBus]          temp_m2_13_3_r;
wire signed [`CalcTempBus]          temp_m2_13_3_i;
wire signed [`CalcTempBus]          temp_m2_13_4_r;
wire signed [`CalcTempBus]          temp_m2_13_4_i;
wire signed [`CalcTempBus]          temp_m2_13_5_r;
wire signed [`CalcTempBus]          temp_m2_13_5_i;
wire signed [`CalcTempBus]          temp_m2_13_6_r;
wire signed [`CalcTempBus]          temp_m2_13_6_i;
wire signed [`CalcTempBus]          temp_m2_13_7_r;
wire signed [`CalcTempBus]          temp_m2_13_7_i;
wire signed [`CalcTempBus]          temp_m2_13_8_r;
wire signed [`CalcTempBus]          temp_m2_13_8_i;
wire signed [`CalcTempBus]          temp_m2_13_9_r;
wire signed [`CalcTempBus]          temp_m2_13_9_i;
wire signed [`CalcTempBus]          temp_m2_13_10_r;
wire signed [`CalcTempBus]          temp_m2_13_10_i;
wire signed [`CalcTempBus]          temp_m2_13_11_r;
wire signed [`CalcTempBus]          temp_m2_13_11_i;
wire signed [`CalcTempBus]          temp_m2_13_12_r;
wire signed [`CalcTempBus]          temp_m2_13_12_i;
wire signed [`CalcTempBus]          temp_m2_13_13_r;
wire signed [`CalcTempBus]          temp_m2_13_13_i;
wire signed [`CalcTempBus]          temp_m2_13_14_r;
wire signed [`CalcTempBus]          temp_m2_13_14_i;
wire signed [`CalcTempBus]          temp_m2_13_15_r;
wire signed [`CalcTempBus]          temp_m2_13_15_i;
wire signed [`CalcTempBus]          temp_m2_13_16_r;
wire signed [`CalcTempBus]          temp_m2_13_16_i;
wire signed [`CalcTempBus]          temp_m2_13_17_r;
wire signed [`CalcTempBus]          temp_m2_13_17_i;
wire signed [`CalcTempBus]          temp_m2_13_18_r;
wire signed [`CalcTempBus]          temp_m2_13_18_i;
wire signed [`CalcTempBus]          temp_m2_13_19_r;
wire signed [`CalcTempBus]          temp_m2_13_19_i;
wire signed [`CalcTempBus]          temp_m2_13_20_r;
wire signed [`CalcTempBus]          temp_m2_13_20_i;
wire signed [`CalcTempBus]          temp_m2_13_21_r;
wire signed [`CalcTempBus]          temp_m2_13_21_i;
wire signed [`CalcTempBus]          temp_m2_13_22_r;
wire signed [`CalcTempBus]          temp_m2_13_22_i;
wire signed [`CalcTempBus]          temp_m2_13_23_r;
wire signed [`CalcTempBus]          temp_m2_13_23_i;
wire signed [`CalcTempBus]          temp_m2_13_24_r;
wire signed [`CalcTempBus]          temp_m2_13_24_i;
wire signed [`CalcTempBus]          temp_m2_13_25_r;
wire signed [`CalcTempBus]          temp_m2_13_25_i;
wire signed [`CalcTempBus]          temp_m2_13_26_r;
wire signed [`CalcTempBus]          temp_m2_13_26_i;
wire signed [`CalcTempBus]          temp_m2_13_27_r;
wire signed [`CalcTempBus]          temp_m2_13_27_i;
wire signed [`CalcTempBus]          temp_m2_13_28_r;
wire signed [`CalcTempBus]          temp_m2_13_28_i;
wire signed [`CalcTempBus]          temp_m2_13_29_r;
wire signed [`CalcTempBus]          temp_m2_13_29_i;
wire signed [`CalcTempBus]          temp_m2_13_30_r;
wire signed [`CalcTempBus]          temp_m2_13_30_i;
wire signed [`CalcTempBus]          temp_m2_13_31_r;
wire signed [`CalcTempBus]          temp_m2_13_31_i;
wire signed [`CalcTempBus]          temp_m2_13_32_r;
wire signed [`CalcTempBus]          temp_m2_13_32_i;
wire signed [`CalcTempBus]          temp_m2_14_1_r;
wire signed [`CalcTempBus]          temp_m2_14_1_i;
wire signed [`CalcTempBus]          temp_m2_14_2_r;
wire signed [`CalcTempBus]          temp_m2_14_2_i;
wire signed [`CalcTempBus]          temp_m2_14_3_r;
wire signed [`CalcTempBus]          temp_m2_14_3_i;
wire signed [`CalcTempBus]          temp_m2_14_4_r;
wire signed [`CalcTempBus]          temp_m2_14_4_i;
wire signed [`CalcTempBus]          temp_m2_14_5_r;
wire signed [`CalcTempBus]          temp_m2_14_5_i;
wire signed [`CalcTempBus]          temp_m2_14_6_r;
wire signed [`CalcTempBus]          temp_m2_14_6_i;
wire signed [`CalcTempBus]          temp_m2_14_7_r;
wire signed [`CalcTempBus]          temp_m2_14_7_i;
wire signed [`CalcTempBus]          temp_m2_14_8_r;
wire signed [`CalcTempBus]          temp_m2_14_8_i;
wire signed [`CalcTempBus]          temp_m2_14_9_r;
wire signed [`CalcTempBus]          temp_m2_14_9_i;
wire signed [`CalcTempBus]          temp_m2_14_10_r;
wire signed [`CalcTempBus]          temp_m2_14_10_i;
wire signed [`CalcTempBus]          temp_m2_14_11_r;
wire signed [`CalcTempBus]          temp_m2_14_11_i;
wire signed [`CalcTempBus]          temp_m2_14_12_r;
wire signed [`CalcTempBus]          temp_m2_14_12_i;
wire signed [`CalcTempBus]          temp_m2_14_13_r;
wire signed [`CalcTempBus]          temp_m2_14_13_i;
wire signed [`CalcTempBus]          temp_m2_14_14_r;
wire signed [`CalcTempBus]          temp_m2_14_14_i;
wire signed [`CalcTempBus]          temp_m2_14_15_r;
wire signed [`CalcTempBus]          temp_m2_14_15_i;
wire signed [`CalcTempBus]          temp_m2_14_16_r;
wire signed [`CalcTempBus]          temp_m2_14_16_i;
wire signed [`CalcTempBus]          temp_m2_14_17_r;
wire signed [`CalcTempBus]          temp_m2_14_17_i;
wire signed [`CalcTempBus]          temp_m2_14_18_r;
wire signed [`CalcTempBus]          temp_m2_14_18_i;
wire signed [`CalcTempBus]          temp_m2_14_19_r;
wire signed [`CalcTempBus]          temp_m2_14_19_i;
wire signed [`CalcTempBus]          temp_m2_14_20_r;
wire signed [`CalcTempBus]          temp_m2_14_20_i;
wire signed [`CalcTempBus]          temp_m2_14_21_r;
wire signed [`CalcTempBus]          temp_m2_14_21_i;
wire signed [`CalcTempBus]          temp_m2_14_22_r;
wire signed [`CalcTempBus]          temp_m2_14_22_i;
wire signed [`CalcTempBus]          temp_m2_14_23_r;
wire signed [`CalcTempBus]          temp_m2_14_23_i;
wire signed [`CalcTempBus]          temp_m2_14_24_r;
wire signed [`CalcTempBus]          temp_m2_14_24_i;
wire signed [`CalcTempBus]          temp_m2_14_25_r;
wire signed [`CalcTempBus]          temp_m2_14_25_i;
wire signed [`CalcTempBus]          temp_m2_14_26_r;
wire signed [`CalcTempBus]          temp_m2_14_26_i;
wire signed [`CalcTempBus]          temp_m2_14_27_r;
wire signed [`CalcTempBus]          temp_m2_14_27_i;
wire signed [`CalcTempBus]          temp_m2_14_28_r;
wire signed [`CalcTempBus]          temp_m2_14_28_i;
wire signed [`CalcTempBus]          temp_m2_14_29_r;
wire signed [`CalcTempBus]          temp_m2_14_29_i;
wire signed [`CalcTempBus]          temp_m2_14_30_r;
wire signed [`CalcTempBus]          temp_m2_14_30_i;
wire signed [`CalcTempBus]          temp_m2_14_31_r;
wire signed [`CalcTempBus]          temp_m2_14_31_i;
wire signed [`CalcTempBus]          temp_m2_14_32_r;
wire signed [`CalcTempBus]          temp_m2_14_32_i;
wire signed [`CalcTempBus]          temp_m2_15_1_r;
wire signed [`CalcTempBus]          temp_m2_15_1_i;
wire signed [`CalcTempBus]          temp_m2_15_2_r;
wire signed [`CalcTempBus]          temp_m2_15_2_i;
wire signed [`CalcTempBus]          temp_m2_15_3_r;
wire signed [`CalcTempBus]          temp_m2_15_3_i;
wire signed [`CalcTempBus]          temp_m2_15_4_r;
wire signed [`CalcTempBus]          temp_m2_15_4_i;
wire signed [`CalcTempBus]          temp_m2_15_5_r;
wire signed [`CalcTempBus]          temp_m2_15_5_i;
wire signed [`CalcTempBus]          temp_m2_15_6_r;
wire signed [`CalcTempBus]          temp_m2_15_6_i;
wire signed [`CalcTempBus]          temp_m2_15_7_r;
wire signed [`CalcTempBus]          temp_m2_15_7_i;
wire signed [`CalcTempBus]          temp_m2_15_8_r;
wire signed [`CalcTempBus]          temp_m2_15_8_i;
wire signed [`CalcTempBus]          temp_m2_15_9_r;
wire signed [`CalcTempBus]          temp_m2_15_9_i;
wire signed [`CalcTempBus]          temp_m2_15_10_r;
wire signed [`CalcTempBus]          temp_m2_15_10_i;
wire signed [`CalcTempBus]          temp_m2_15_11_r;
wire signed [`CalcTempBus]          temp_m2_15_11_i;
wire signed [`CalcTempBus]          temp_m2_15_12_r;
wire signed [`CalcTempBus]          temp_m2_15_12_i;
wire signed [`CalcTempBus]          temp_m2_15_13_r;
wire signed [`CalcTempBus]          temp_m2_15_13_i;
wire signed [`CalcTempBus]          temp_m2_15_14_r;
wire signed [`CalcTempBus]          temp_m2_15_14_i;
wire signed [`CalcTempBus]          temp_m2_15_15_r;
wire signed [`CalcTempBus]          temp_m2_15_15_i;
wire signed [`CalcTempBus]          temp_m2_15_16_r;
wire signed [`CalcTempBus]          temp_m2_15_16_i;
wire signed [`CalcTempBus]          temp_m2_15_17_r;
wire signed [`CalcTempBus]          temp_m2_15_17_i;
wire signed [`CalcTempBus]          temp_m2_15_18_r;
wire signed [`CalcTempBus]          temp_m2_15_18_i;
wire signed [`CalcTempBus]          temp_m2_15_19_r;
wire signed [`CalcTempBus]          temp_m2_15_19_i;
wire signed [`CalcTempBus]          temp_m2_15_20_r;
wire signed [`CalcTempBus]          temp_m2_15_20_i;
wire signed [`CalcTempBus]          temp_m2_15_21_r;
wire signed [`CalcTempBus]          temp_m2_15_21_i;
wire signed [`CalcTempBus]          temp_m2_15_22_r;
wire signed [`CalcTempBus]          temp_m2_15_22_i;
wire signed [`CalcTempBus]          temp_m2_15_23_r;
wire signed [`CalcTempBus]          temp_m2_15_23_i;
wire signed [`CalcTempBus]          temp_m2_15_24_r;
wire signed [`CalcTempBus]          temp_m2_15_24_i;
wire signed [`CalcTempBus]          temp_m2_15_25_r;
wire signed [`CalcTempBus]          temp_m2_15_25_i;
wire signed [`CalcTempBus]          temp_m2_15_26_r;
wire signed [`CalcTempBus]          temp_m2_15_26_i;
wire signed [`CalcTempBus]          temp_m2_15_27_r;
wire signed [`CalcTempBus]          temp_m2_15_27_i;
wire signed [`CalcTempBus]          temp_m2_15_28_r;
wire signed [`CalcTempBus]          temp_m2_15_28_i;
wire signed [`CalcTempBus]          temp_m2_15_29_r;
wire signed [`CalcTempBus]          temp_m2_15_29_i;
wire signed [`CalcTempBus]          temp_m2_15_30_r;
wire signed [`CalcTempBus]          temp_m2_15_30_i;
wire signed [`CalcTempBus]          temp_m2_15_31_r;
wire signed [`CalcTempBus]          temp_m2_15_31_i;
wire signed [`CalcTempBus]          temp_m2_15_32_r;
wire signed [`CalcTempBus]          temp_m2_15_32_i;
wire signed [`CalcTempBus]          temp_m2_16_1_r;
wire signed [`CalcTempBus]          temp_m2_16_1_i;
wire signed [`CalcTempBus]          temp_m2_16_2_r;
wire signed [`CalcTempBus]          temp_m2_16_2_i;
wire signed [`CalcTempBus]          temp_m2_16_3_r;
wire signed [`CalcTempBus]          temp_m2_16_3_i;
wire signed [`CalcTempBus]          temp_m2_16_4_r;
wire signed [`CalcTempBus]          temp_m2_16_4_i;
wire signed [`CalcTempBus]          temp_m2_16_5_r;
wire signed [`CalcTempBus]          temp_m2_16_5_i;
wire signed [`CalcTempBus]          temp_m2_16_6_r;
wire signed [`CalcTempBus]          temp_m2_16_6_i;
wire signed [`CalcTempBus]          temp_m2_16_7_r;
wire signed [`CalcTempBus]          temp_m2_16_7_i;
wire signed [`CalcTempBus]          temp_m2_16_8_r;
wire signed [`CalcTempBus]          temp_m2_16_8_i;
wire signed [`CalcTempBus]          temp_m2_16_9_r;
wire signed [`CalcTempBus]          temp_m2_16_9_i;
wire signed [`CalcTempBus]          temp_m2_16_10_r;
wire signed [`CalcTempBus]          temp_m2_16_10_i;
wire signed [`CalcTempBus]          temp_m2_16_11_r;
wire signed [`CalcTempBus]          temp_m2_16_11_i;
wire signed [`CalcTempBus]          temp_m2_16_12_r;
wire signed [`CalcTempBus]          temp_m2_16_12_i;
wire signed [`CalcTempBus]          temp_m2_16_13_r;
wire signed [`CalcTempBus]          temp_m2_16_13_i;
wire signed [`CalcTempBus]          temp_m2_16_14_r;
wire signed [`CalcTempBus]          temp_m2_16_14_i;
wire signed [`CalcTempBus]          temp_m2_16_15_r;
wire signed [`CalcTempBus]          temp_m2_16_15_i;
wire signed [`CalcTempBus]          temp_m2_16_16_r;
wire signed [`CalcTempBus]          temp_m2_16_16_i;
wire signed [`CalcTempBus]          temp_m2_16_17_r;
wire signed [`CalcTempBus]          temp_m2_16_17_i;
wire signed [`CalcTempBus]          temp_m2_16_18_r;
wire signed [`CalcTempBus]          temp_m2_16_18_i;
wire signed [`CalcTempBus]          temp_m2_16_19_r;
wire signed [`CalcTempBus]          temp_m2_16_19_i;
wire signed [`CalcTempBus]          temp_m2_16_20_r;
wire signed [`CalcTempBus]          temp_m2_16_20_i;
wire signed [`CalcTempBus]          temp_m2_16_21_r;
wire signed [`CalcTempBus]          temp_m2_16_21_i;
wire signed [`CalcTempBus]          temp_m2_16_22_r;
wire signed [`CalcTempBus]          temp_m2_16_22_i;
wire signed [`CalcTempBus]          temp_m2_16_23_r;
wire signed [`CalcTempBus]          temp_m2_16_23_i;
wire signed [`CalcTempBus]          temp_m2_16_24_r;
wire signed [`CalcTempBus]          temp_m2_16_24_i;
wire signed [`CalcTempBus]          temp_m2_16_25_r;
wire signed [`CalcTempBus]          temp_m2_16_25_i;
wire signed [`CalcTempBus]          temp_m2_16_26_r;
wire signed [`CalcTempBus]          temp_m2_16_26_i;
wire signed [`CalcTempBus]          temp_m2_16_27_r;
wire signed [`CalcTempBus]          temp_m2_16_27_i;
wire signed [`CalcTempBus]          temp_m2_16_28_r;
wire signed [`CalcTempBus]          temp_m2_16_28_i;
wire signed [`CalcTempBus]          temp_m2_16_29_r;
wire signed [`CalcTempBus]          temp_m2_16_29_i;
wire signed [`CalcTempBus]          temp_m2_16_30_r;
wire signed [`CalcTempBus]          temp_m2_16_30_i;
wire signed [`CalcTempBus]          temp_m2_16_31_r;
wire signed [`CalcTempBus]          temp_m2_16_31_i;
wire signed [`CalcTempBus]          temp_m2_16_32_r;
wire signed [`CalcTempBus]          temp_m2_16_32_i;
wire signed [`CalcTempBus]          temp_m2_17_1_r;
wire signed [`CalcTempBus]          temp_m2_17_1_i;
wire signed [`CalcTempBus]          temp_m2_17_2_r;
wire signed [`CalcTempBus]          temp_m2_17_2_i;
wire signed [`CalcTempBus]          temp_m2_17_3_r;
wire signed [`CalcTempBus]          temp_m2_17_3_i;
wire signed [`CalcTempBus]          temp_m2_17_4_r;
wire signed [`CalcTempBus]          temp_m2_17_4_i;
wire signed [`CalcTempBus]          temp_m2_17_5_r;
wire signed [`CalcTempBus]          temp_m2_17_5_i;
wire signed [`CalcTempBus]          temp_m2_17_6_r;
wire signed [`CalcTempBus]          temp_m2_17_6_i;
wire signed [`CalcTempBus]          temp_m2_17_7_r;
wire signed [`CalcTempBus]          temp_m2_17_7_i;
wire signed [`CalcTempBus]          temp_m2_17_8_r;
wire signed [`CalcTempBus]          temp_m2_17_8_i;
wire signed [`CalcTempBus]          temp_m2_17_9_r;
wire signed [`CalcTempBus]          temp_m2_17_9_i;
wire signed [`CalcTempBus]          temp_m2_17_10_r;
wire signed [`CalcTempBus]          temp_m2_17_10_i;
wire signed [`CalcTempBus]          temp_m2_17_11_r;
wire signed [`CalcTempBus]          temp_m2_17_11_i;
wire signed [`CalcTempBus]          temp_m2_17_12_r;
wire signed [`CalcTempBus]          temp_m2_17_12_i;
wire signed [`CalcTempBus]          temp_m2_17_13_r;
wire signed [`CalcTempBus]          temp_m2_17_13_i;
wire signed [`CalcTempBus]          temp_m2_17_14_r;
wire signed [`CalcTempBus]          temp_m2_17_14_i;
wire signed [`CalcTempBus]          temp_m2_17_15_r;
wire signed [`CalcTempBus]          temp_m2_17_15_i;
wire signed [`CalcTempBus]          temp_m2_17_16_r;
wire signed [`CalcTempBus]          temp_m2_17_16_i;
wire signed [`CalcTempBus]          temp_m2_17_17_r;
wire signed [`CalcTempBus]          temp_m2_17_17_i;
wire signed [`CalcTempBus]          temp_m2_17_18_r;
wire signed [`CalcTempBus]          temp_m2_17_18_i;
wire signed [`CalcTempBus]          temp_m2_17_19_r;
wire signed [`CalcTempBus]          temp_m2_17_19_i;
wire signed [`CalcTempBus]          temp_m2_17_20_r;
wire signed [`CalcTempBus]          temp_m2_17_20_i;
wire signed [`CalcTempBus]          temp_m2_17_21_r;
wire signed [`CalcTempBus]          temp_m2_17_21_i;
wire signed [`CalcTempBus]          temp_m2_17_22_r;
wire signed [`CalcTempBus]          temp_m2_17_22_i;
wire signed [`CalcTempBus]          temp_m2_17_23_r;
wire signed [`CalcTempBus]          temp_m2_17_23_i;
wire signed [`CalcTempBus]          temp_m2_17_24_r;
wire signed [`CalcTempBus]          temp_m2_17_24_i;
wire signed [`CalcTempBus]          temp_m2_17_25_r;
wire signed [`CalcTempBus]          temp_m2_17_25_i;
wire signed [`CalcTempBus]          temp_m2_17_26_r;
wire signed [`CalcTempBus]          temp_m2_17_26_i;
wire signed [`CalcTempBus]          temp_m2_17_27_r;
wire signed [`CalcTempBus]          temp_m2_17_27_i;
wire signed [`CalcTempBus]          temp_m2_17_28_r;
wire signed [`CalcTempBus]          temp_m2_17_28_i;
wire signed [`CalcTempBus]          temp_m2_17_29_r;
wire signed [`CalcTempBus]          temp_m2_17_29_i;
wire signed [`CalcTempBus]          temp_m2_17_30_r;
wire signed [`CalcTempBus]          temp_m2_17_30_i;
wire signed [`CalcTempBus]          temp_m2_17_31_r;
wire signed [`CalcTempBus]          temp_m2_17_31_i;
wire signed [`CalcTempBus]          temp_m2_17_32_r;
wire signed [`CalcTempBus]          temp_m2_17_32_i;
wire signed [`CalcTempBus]          temp_m2_18_1_r;
wire signed [`CalcTempBus]          temp_m2_18_1_i;
wire signed [`CalcTempBus]          temp_m2_18_2_r;
wire signed [`CalcTempBus]          temp_m2_18_2_i;
wire signed [`CalcTempBus]          temp_m2_18_3_r;
wire signed [`CalcTempBus]          temp_m2_18_3_i;
wire signed [`CalcTempBus]          temp_m2_18_4_r;
wire signed [`CalcTempBus]          temp_m2_18_4_i;
wire signed [`CalcTempBus]          temp_m2_18_5_r;
wire signed [`CalcTempBus]          temp_m2_18_5_i;
wire signed [`CalcTempBus]          temp_m2_18_6_r;
wire signed [`CalcTempBus]          temp_m2_18_6_i;
wire signed [`CalcTempBus]          temp_m2_18_7_r;
wire signed [`CalcTempBus]          temp_m2_18_7_i;
wire signed [`CalcTempBus]          temp_m2_18_8_r;
wire signed [`CalcTempBus]          temp_m2_18_8_i;
wire signed [`CalcTempBus]          temp_m2_18_9_r;
wire signed [`CalcTempBus]          temp_m2_18_9_i;
wire signed [`CalcTempBus]          temp_m2_18_10_r;
wire signed [`CalcTempBus]          temp_m2_18_10_i;
wire signed [`CalcTempBus]          temp_m2_18_11_r;
wire signed [`CalcTempBus]          temp_m2_18_11_i;
wire signed [`CalcTempBus]          temp_m2_18_12_r;
wire signed [`CalcTempBus]          temp_m2_18_12_i;
wire signed [`CalcTempBus]          temp_m2_18_13_r;
wire signed [`CalcTempBus]          temp_m2_18_13_i;
wire signed [`CalcTempBus]          temp_m2_18_14_r;
wire signed [`CalcTempBus]          temp_m2_18_14_i;
wire signed [`CalcTempBus]          temp_m2_18_15_r;
wire signed [`CalcTempBus]          temp_m2_18_15_i;
wire signed [`CalcTempBus]          temp_m2_18_16_r;
wire signed [`CalcTempBus]          temp_m2_18_16_i;
wire signed [`CalcTempBus]          temp_m2_18_17_r;
wire signed [`CalcTempBus]          temp_m2_18_17_i;
wire signed [`CalcTempBus]          temp_m2_18_18_r;
wire signed [`CalcTempBus]          temp_m2_18_18_i;
wire signed [`CalcTempBus]          temp_m2_18_19_r;
wire signed [`CalcTempBus]          temp_m2_18_19_i;
wire signed [`CalcTempBus]          temp_m2_18_20_r;
wire signed [`CalcTempBus]          temp_m2_18_20_i;
wire signed [`CalcTempBus]          temp_m2_18_21_r;
wire signed [`CalcTempBus]          temp_m2_18_21_i;
wire signed [`CalcTempBus]          temp_m2_18_22_r;
wire signed [`CalcTempBus]          temp_m2_18_22_i;
wire signed [`CalcTempBus]          temp_m2_18_23_r;
wire signed [`CalcTempBus]          temp_m2_18_23_i;
wire signed [`CalcTempBus]          temp_m2_18_24_r;
wire signed [`CalcTempBus]          temp_m2_18_24_i;
wire signed [`CalcTempBus]          temp_m2_18_25_r;
wire signed [`CalcTempBus]          temp_m2_18_25_i;
wire signed [`CalcTempBus]          temp_m2_18_26_r;
wire signed [`CalcTempBus]          temp_m2_18_26_i;
wire signed [`CalcTempBus]          temp_m2_18_27_r;
wire signed [`CalcTempBus]          temp_m2_18_27_i;
wire signed [`CalcTempBus]          temp_m2_18_28_r;
wire signed [`CalcTempBus]          temp_m2_18_28_i;
wire signed [`CalcTempBus]          temp_m2_18_29_r;
wire signed [`CalcTempBus]          temp_m2_18_29_i;
wire signed [`CalcTempBus]          temp_m2_18_30_r;
wire signed [`CalcTempBus]          temp_m2_18_30_i;
wire signed [`CalcTempBus]          temp_m2_18_31_r;
wire signed [`CalcTempBus]          temp_m2_18_31_i;
wire signed [`CalcTempBus]          temp_m2_18_32_r;
wire signed [`CalcTempBus]          temp_m2_18_32_i;
wire signed [`CalcTempBus]          temp_m2_19_1_r;
wire signed [`CalcTempBus]          temp_m2_19_1_i;
wire signed [`CalcTempBus]          temp_m2_19_2_r;
wire signed [`CalcTempBus]          temp_m2_19_2_i;
wire signed [`CalcTempBus]          temp_m2_19_3_r;
wire signed [`CalcTempBus]          temp_m2_19_3_i;
wire signed [`CalcTempBus]          temp_m2_19_4_r;
wire signed [`CalcTempBus]          temp_m2_19_4_i;
wire signed [`CalcTempBus]          temp_m2_19_5_r;
wire signed [`CalcTempBus]          temp_m2_19_5_i;
wire signed [`CalcTempBus]          temp_m2_19_6_r;
wire signed [`CalcTempBus]          temp_m2_19_6_i;
wire signed [`CalcTempBus]          temp_m2_19_7_r;
wire signed [`CalcTempBus]          temp_m2_19_7_i;
wire signed [`CalcTempBus]          temp_m2_19_8_r;
wire signed [`CalcTempBus]          temp_m2_19_8_i;
wire signed [`CalcTempBus]          temp_m2_19_9_r;
wire signed [`CalcTempBus]          temp_m2_19_9_i;
wire signed [`CalcTempBus]          temp_m2_19_10_r;
wire signed [`CalcTempBus]          temp_m2_19_10_i;
wire signed [`CalcTempBus]          temp_m2_19_11_r;
wire signed [`CalcTempBus]          temp_m2_19_11_i;
wire signed [`CalcTempBus]          temp_m2_19_12_r;
wire signed [`CalcTempBus]          temp_m2_19_12_i;
wire signed [`CalcTempBus]          temp_m2_19_13_r;
wire signed [`CalcTempBus]          temp_m2_19_13_i;
wire signed [`CalcTempBus]          temp_m2_19_14_r;
wire signed [`CalcTempBus]          temp_m2_19_14_i;
wire signed [`CalcTempBus]          temp_m2_19_15_r;
wire signed [`CalcTempBus]          temp_m2_19_15_i;
wire signed [`CalcTempBus]          temp_m2_19_16_r;
wire signed [`CalcTempBus]          temp_m2_19_16_i;
wire signed [`CalcTempBus]          temp_m2_19_17_r;
wire signed [`CalcTempBus]          temp_m2_19_17_i;
wire signed [`CalcTempBus]          temp_m2_19_18_r;
wire signed [`CalcTempBus]          temp_m2_19_18_i;
wire signed [`CalcTempBus]          temp_m2_19_19_r;
wire signed [`CalcTempBus]          temp_m2_19_19_i;
wire signed [`CalcTempBus]          temp_m2_19_20_r;
wire signed [`CalcTempBus]          temp_m2_19_20_i;
wire signed [`CalcTempBus]          temp_m2_19_21_r;
wire signed [`CalcTempBus]          temp_m2_19_21_i;
wire signed [`CalcTempBus]          temp_m2_19_22_r;
wire signed [`CalcTempBus]          temp_m2_19_22_i;
wire signed [`CalcTempBus]          temp_m2_19_23_r;
wire signed [`CalcTempBus]          temp_m2_19_23_i;
wire signed [`CalcTempBus]          temp_m2_19_24_r;
wire signed [`CalcTempBus]          temp_m2_19_24_i;
wire signed [`CalcTempBus]          temp_m2_19_25_r;
wire signed [`CalcTempBus]          temp_m2_19_25_i;
wire signed [`CalcTempBus]          temp_m2_19_26_r;
wire signed [`CalcTempBus]          temp_m2_19_26_i;
wire signed [`CalcTempBus]          temp_m2_19_27_r;
wire signed [`CalcTempBus]          temp_m2_19_27_i;
wire signed [`CalcTempBus]          temp_m2_19_28_r;
wire signed [`CalcTempBus]          temp_m2_19_28_i;
wire signed [`CalcTempBus]          temp_m2_19_29_r;
wire signed [`CalcTempBus]          temp_m2_19_29_i;
wire signed [`CalcTempBus]          temp_m2_19_30_r;
wire signed [`CalcTempBus]          temp_m2_19_30_i;
wire signed [`CalcTempBus]          temp_m2_19_31_r;
wire signed [`CalcTempBus]          temp_m2_19_31_i;
wire signed [`CalcTempBus]          temp_m2_19_32_r;
wire signed [`CalcTempBus]          temp_m2_19_32_i;
wire signed [`CalcTempBus]          temp_m2_20_1_r;
wire signed [`CalcTempBus]          temp_m2_20_1_i;
wire signed [`CalcTempBus]          temp_m2_20_2_r;
wire signed [`CalcTempBus]          temp_m2_20_2_i;
wire signed [`CalcTempBus]          temp_m2_20_3_r;
wire signed [`CalcTempBus]          temp_m2_20_3_i;
wire signed [`CalcTempBus]          temp_m2_20_4_r;
wire signed [`CalcTempBus]          temp_m2_20_4_i;
wire signed [`CalcTempBus]          temp_m2_20_5_r;
wire signed [`CalcTempBus]          temp_m2_20_5_i;
wire signed [`CalcTempBus]          temp_m2_20_6_r;
wire signed [`CalcTempBus]          temp_m2_20_6_i;
wire signed [`CalcTempBus]          temp_m2_20_7_r;
wire signed [`CalcTempBus]          temp_m2_20_7_i;
wire signed [`CalcTempBus]          temp_m2_20_8_r;
wire signed [`CalcTempBus]          temp_m2_20_8_i;
wire signed [`CalcTempBus]          temp_m2_20_9_r;
wire signed [`CalcTempBus]          temp_m2_20_9_i;
wire signed [`CalcTempBus]          temp_m2_20_10_r;
wire signed [`CalcTempBus]          temp_m2_20_10_i;
wire signed [`CalcTempBus]          temp_m2_20_11_r;
wire signed [`CalcTempBus]          temp_m2_20_11_i;
wire signed [`CalcTempBus]          temp_m2_20_12_r;
wire signed [`CalcTempBus]          temp_m2_20_12_i;
wire signed [`CalcTempBus]          temp_m2_20_13_r;
wire signed [`CalcTempBus]          temp_m2_20_13_i;
wire signed [`CalcTempBus]          temp_m2_20_14_r;
wire signed [`CalcTempBus]          temp_m2_20_14_i;
wire signed [`CalcTempBus]          temp_m2_20_15_r;
wire signed [`CalcTempBus]          temp_m2_20_15_i;
wire signed [`CalcTempBus]          temp_m2_20_16_r;
wire signed [`CalcTempBus]          temp_m2_20_16_i;
wire signed [`CalcTempBus]          temp_m2_20_17_r;
wire signed [`CalcTempBus]          temp_m2_20_17_i;
wire signed [`CalcTempBus]          temp_m2_20_18_r;
wire signed [`CalcTempBus]          temp_m2_20_18_i;
wire signed [`CalcTempBus]          temp_m2_20_19_r;
wire signed [`CalcTempBus]          temp_m2_20_19_i;
wire signed [`CalcTempBus]          temp_m2_20_20_r;
wire signed [`CalcTempBus]          temp_m2_20_20_i;
wire signed [`CalcTempBus]          temp_m2_20_21_r;
wire signed [`CalcTempBus]          temp_m2_20_21_i;
wire signed [`CalcTempBus]          temp_m2_20_22_r;
wire signed [`CalcTempBus]          temp_m2_20_22_i;
wire signed [`CalcTempBus]          temp_m2_20_23_r;
wire signed [`CalcTempBus]          temp_m2_20_23_i;
wire signed [`CalcTempBus]          temp_m2_20_24_r;
wire signed [`CalcTempBus]          temp_m2_20_24_i;
wire signed [`CalcTempBus]          temp_m2_20_25_r;
wire signed [`CalcTempBus]          temp_m2_20_25_i;
wire signed [`CalcTempBus]          temp_m2_20_26_r;
wire signed [`CalcTempBus]          temp_m2_20_26_i;
wire signed [`CalcTempBus]          temp_m2_20_27_r;
wire signed [`CalcTempBus]          temp_m2_20_27_i;
wire signed [`CalcTempBus]          temp_m2_20_28_r;
wire signed [`CalcTempBus]          temp_m2_20_28_i;
wire signed [`CalcTempBus]          temp_m2_20_29_r;
wire signed [`CalcTempBus]          temp_m2_20_29_i;
wire signed [`CalcTempBus]          temp_m2_20_30_r;
wire signed [`CalcTempBus]          temp_m2_20_30_i;
wire signed [`CalcTempBus]          temp_m2_20_31_r;
wire signed [`CalcTempBus]          temp_m2_20_31_i;
wire signed [`CalcTempBus]          temp_m2_20_32_r;
wire signed [`CalcTempBus]          temp_m2_20_32_i;
wire signed [`CalcTempBus]          temp_m2_21_1_r;
wire signed [`CalcTempBus]          temp_m2_21_1_i;
wire signed [`CalcTempBus]          temp_m2_21_2_r;
wire signed [`CalcTempBus]          temp_m2_21_2_i;
wire signed [`CalcTempBus]          temp_m2_21_3_r;
wire signed [`CalcTempBus]          temp_m2_21_3_i;
wire signed [`CalcTempBus]          temp_m2_21_4_r;
wire signed [`CalcTempBus]          temp_m2_21_4_i;
wire signed [`CalcTempBus]          temp_m2_21_5_r;
wire signed [`CalcTempBus]          temp_m2_21_5_i;
wire signed [`CalcTempBus]          temp_m2_21_6_r;
wire signed [`CalcTempBus]          temp_m2_21_6_i;
wire signed [`CalcTempBus]          temp_m2_21_7_r;
wire signed [`CalcTempBus]          temp_m2_21_7_i;
wire signed [`CalcTempBus]          temp_m2_21_8_r;
wire signed [`CalcTempBus]          temp_m2_21_8_i;
wire signed [`CalcTempBus]          temp_m2_21_9_r;
wire signed [`CalcTempBus]          temp_m2_21_9_i;
wire signed [`CalcTempBus]          temp_m2_21_10_r;
wire signed [`CalcTempBus]          temp_m2_21_10_i;
wire signed [`CalcTempBus]          temp_m2_21_11_r;
wire signed [`CalcTempBus]          temp_m2_21_11_i;
wire signed [`CalcTempBus]          temp_m2_21_12_r;
wire signed [`CalcTempBus]          temp_m2_21_12_i;
wire signed [`CalcTempBus]          temp_m2_21_13_r;
wire signed [`CalcTempBus]          temp_m2_21_13_i;
wire signed [`CalcTempBus]          temp_m2_21_14_r;
wire signed [`CalcTempBus]          temp_m2_21_14_i;
wire signed [`CalcTempBus]          temp_m2_21_15_r;
wire signed [`CalcTempBus]          temp_m2_21_15_i;
wire signed [`CalcTempBus]          temp_m2_21_16_r;
wire signed [`CalcTempBus]          temp_m2_21_16_i;
wire signed [`CalcTempBus]          temp_m2_21_17_r;
wire signed [`CalcTempBus]          temp_m2_21_17_i;
wire signed [`CalcTempBus]          temp_m2_21_18_r;
wire signed [`CalcTempBus]          temp_m2_21_18_i;
wire signed [`CalcTempBus]          temp_m2_21_19_r;
wire signed [`CalcTempBus]          temp_m2_21_19_i;
wire signed [`CalcTempBus]          temp_m2_21_20_r;
wire signed [`CalcTempBus]          temp_m2_21_20_i;
wire signed [`CalcTempBus]          temp_m2_21_21_r;
wire signed [`CalcTempBus]          temp_m2_21_21_i;
wire signed [`CalcTempBus]          temp_m2_21_22_r;
wire signed [`CalcTempBus]          temp_m2_21_22_i;
wire signed [`CalcTempBus]          temp_m2_21_23_r;
wire signed [`CalcTempBus]          temp_m2_21_23_i;
wire signed [`CalcTempBus]          temp_m2_21_24_r;
wire signed [`CalcTempBus]          temp_m2_21_24_i;
wire signed [`CalcTempBus]          temp_m2_21_25_r;
wire signed [`CalcTempBus]          temp_m2_21_25_i;
wire signed [`CalcTempBus]          temp_m2_21_26_r;
wire signed [`CalcTempBus]          temp_m2_21_26_i;
wire signed [`CalcTempBus]          temp_m2_21_27_r;
wire signed [`CalcTempBus]          temp_m2_21_27_i;
wire signed [`CalcTempBus]          temp_m2_21_28_r;
wire signed [`CalcTempBus]          temp_m2_21_28_i;
wire signed [`CalcTempBus]          temp_m2_21_29_r;
wire signed [`CalcTempBus]          temp_m2_21_29_i;
wire signed [`CalcTempBus]          temp_m2_21_30_r;
wire signed [`CalcTempBus]          temp_m2_21_30_i;
wire signed [`CalcTempBus]          temp_m2_21_31_r;
wire signed [`CalcTempBus]          temp_m2_21_31_i;
wire signed [`CalcTempBus]          temp_m2_21_32_r;
wire signed [`CalcTempBus]          temp_m2_21_32_i;
wire signed [`CalcTempBus]          temp_m2_22_1_r;
wire signed [`CalcTempBus]          temp_m2_22_1_i;
wire signed [`CalcTempBus]          temp_m2_22_2_r;
wire signed [`CalcTempBus]          temp_m2_22_2_i;
wire signed [`CalcTempBus]          temp_m2_22_3_r;
wire signed [`CalcTempBus]          temp_m2_22_3_i;
wire signed [`CalcTempBus]          temp_m2_22_4_r;
wire signed [`CalcTempBus]          temp_m2_22_4_i;
wire signed [`CalcTempBus]          temp_m2_22_5_r;
wire signed [`CalcTempBus]          temp_m2_22_5_i;
wire signed [`CalcTempBus]          temp_m2_22_6_r;
wire signed [`CalcTempBus]          temp_m2_22_6_i;
wire signed [`CalcTempBus]          temp_m2_22_7_r;
wire signed [`CalcTempBus]          temp_m2_22_7_i;
wire signed [`CalcTempBus]          temp_m2_22_8_r;
wire signed [`CalcTempBus]          temp_m2_22_8_i;
wire signed [`CalcTempBus]          temp_m2_22_9_r;
wire signed [`CalcTempBus]          temp_m2_22_9_i;
wire signed [`CalcTempBus]          temp_m2_22_10_r;
wire signed [`CalcTempBus]          temp_m2_22_10_i;
wire signed [`CalcTempBus]          temp_m2_22_11_r;
wire signed [`CalcTempBus]          temp_m2_22_11_i;
wire signed [`CalcTempBus]          temp_m2_22_12_r;
wire signed [`CalcTempBus]          temp_m2_22_12_i;
wire signed [`CalcTempBus]          temp_m2_22_13_r;
wire signed [`CalcTempBus]          temp_m2_22_13_i;
wire signed [`CalcTempBus]          temp_m2_22_14_r;
wire signed [`CalcTempBus]          temp_m2_22_14_i;
wire signed [`CalcTempBus]          temp_m2_22_15_r;
wire signed [`CalcTempBus]          temp_m2_22_15_i;
wire signed [`CalcTempBus]          temp_m2_22_16_r;
wire signed [`CalcTempBus]          temp_m2_22_16_i;
wire signed [`CalcTempBus]          temp_m2_22_17_r;
wire signed [`CalcTempBus]          temp_m2_22_17_i;
wire signed [`CalcTempBus]          temp_m2_22_18_r;
wire signed [`CalcTempBus]          temp_m2_22_18_i;
wire signed [`CalcTempBus]          temp_m2_22_19_r;
wire signed [`CalcTempBus]          temp_m2_22_19_i;
wire signed [`CalcTempBus]          temp_m2_22_20_r;
wire signed [`CalcTempBus]          temp_m2_22_20_i;
wire signed [`CalcTempBus]          temp_m2_22_21_r;
wire signed [`CalcTempBus]          temp_m2_22_21_i;
wire signed [`CalcTempBus]          temp_m2_22_22_r;
wire signed [`CalcTempBus]          temp_m2_22_22_i;
wire signed [`CalcTempBus]          temp_m2_22_23_r;
wire signed [`CalcTempBus]          temp_m2_22_23_i;
wire signed [`CalcTempBus]          temp_m2_22_24_r;
wire signed [`CalcTempBus]          temp_m2_22_24_i;
wire signed [`CalcTempBus]          temp_m2_22_25_r;
wire signed [`CalcTempBus]          temp_m2_22_25_i;
wire signed [`CalcTempBus]          temp_m2_22_26_r;
wire signed [`CalcTempBus]          temp_m2_22_26_i;
wire signed [`CalcTempBus]          temp_m2_22_27_r;
wire signed [`CalcTempBus]          temp_m2_22_27_i;
wire signed [`CalcTempBus]          temp_m2_22_28_r;
wire signed [`CalcTempBus]          temp_m2_22_28_i;
wire signed [`CalcTempBus]          temp_m2_22_29_r;
wire signed [`CalcTempBus]          temp_m2_22_29_i;
wire signed [`CalcTempBus]          temp_m2_22_30_r;
wire signed [`CalcTempBus]          temp_m2_22_30_i;
wire signed [`CalcTempBus]          temp_m2_22_31_r;
wire signed [`CalcTempBus]          temp_m2_22_31_i;
wire signed [`CalcTempBus]          temp_m2_22_32_r;
wire signed [`CalcTempBus]          temp_m2_22_32_i;
wire signed [`CalcTempBus]          temp_m2_23_1_r;
wire signed [`CalcTempBus]          temp_m2_23_1_i;
wire signed [`CalcTempBus]          temp_m2_23_2_r;
wire signed [`CalcTempBus]          temp_m2_23_2_i;
wire signed [`CalcTempBus]          temp_m2_23_3_r;
wire signed [`CalcTempBus]          temp_m2_23_3_i;
wire signed [`CalcTempBus]          temp_m2_23_4_r;
wire signed [`CalcTempBus]          temp_m2_23_4_i;
wire signed [`CalcTempBus]          temp_m2_23_5_r;
wire signed [`CalcTempBus]          temp_m2_23_5_i;
wire signed [`CalcTempBus]          temp_m2_23_6_r;
wire signed [`CalcTempBus]          temp_m2_23_6_i;
wire signed [`CalcTempBus]          temp_m2_23_7_r;
wire signed [`CalcTempBus]          temp_m2_23_7_i;
wire signed [`CalcTempBus]          temp_m2_23_8_r;
wire signed [`CalcTempBus]          temp_m2_23_8_i;
wire signed [`CalcTempBus]          temp_m2_23_9_r;
wire signed [`CalcTempBus]          temp_m2_23_9_i;
wire signed [`CalcTempBus]          temp_m2_23_10_r;
wire signed [`CalcTempBus]          temp_m2_23_10_i;
wire signed [`CalcTempBus]          temp_m2_23_11_r;
wire signed [`CalcTempBus]          temp_m2_23_11_i;
wire signed [`CalcTempBus]          temp_m2_23_12_r;
wire signed [`CalcTempBus]          temp_m2_23_12_i;
wire signed [`CalcTempBus]          temp_m2_23_13_r;
wire signed [`CalcTempBus]          temp_m2_23_13_i;
wire signed [`CalcTempBus]          temp_m2_23_14_r;
wire signed [`CalcTempBus]          temp_m2_23_14_i;
wire signed [`CalcTempBus]          temp_m2_23_15_r;
wire signed [`CalcTempBus]          temp_m2_23_15_i;
wire signed [`CalcTempBus]          temp_m2_23_16_r;
wire signed [`CalcTempBus]          temp_m2_23_16_i;
wire signed [`CalcTempBus]          temp_m2_23_17_r;
wire signed [`CalcTempBus]          temp_m2_23_17_i;
wire signed [`CalcTempBus]          temp_m2_23_18_r;
wire signed [`CalcTempBus]          temp_m2_23_18_i;
wire signed [`CalcTempBus]          temp_m2_23_19_r;
wire signed [`CalcTempBus]          temp_m2_23_19_i;
wire signed [`CalcTempBus]          temp_m2_23_20_r;
wire signed [`CalcTempBus]          temp_m2_23_20_i;
wire signed [`CalcTempBus]          temp_m2_23_21_r;
wire signed [`CalcTempBus]          temp_m2_23_21_i;
wire signed [`CalcTempBus]          temp_m2_23_22_r;
wire signed [`CalcTempBus]          temp_m2_23_22_i;
wire signed [`CalcTempBus]          temp_m2_23_23_r;
wire signed [`CalcTempBus]          temp_m2_23_23_i;
wire signed [`CalcTempBus]          temp_m2_23_24_r;
wire signed [`CalcTempBus]          temp_m2_23_24_i;
wire signed [`CalcTempBus]          temp_m2_23_25_r;
wire signed [`CalcTempBus]          temp_m2_23_25_i;
wire signed [`CalcTempBus]          temp_m2_23_26_r;
wire signed [`CalcTempBus]          temp_m2_23_26_i;
wire signed [`CalcTempBus]          temp_m2_23_27_r;
wire signed [`CalcTempBus]          temp_m2_23_27_i;
wire signed [`CalcTempBus]          temp_m2_23_28_r;
wire signed [`CalcTempBus]          temp_m2_23_28_i;
wire signed [`CalcTempBus]          temp_m2_23_29_r;
wire signed [`CalcTempBus]          temp_m2_23_29_i;
wire signed [`CalcTempBus]          temp_m2_23_30_r;
wire signed [`CalcTempBus]          temp_m2_23_30_i;
wire signed [`CalcTempBus]          temp_m2_23_31_r;
wire signed [`CalcTempBus]          temp_m2_23_31_i;
wire signed [`CalcTempBus]          temp_m2_23_32_r;
wire signed [`CalcTempBus]          temp_m2_23_32_i;
wire signed [`CalcTempBus]          temp_m2_24_1_r;
wire signed [`CalcTempBus]          temp_m2_24_1_i;
wire signed [`CalcTempBus]          temp_m2_24_2_r;
wire signed [`CalcTempBus]          temp_m2_24_2_i;
wire signed [`CalcTempBus]          temp_m2_24_3_r;
wire signed [`CalcTempBus]          temp_m2_24_3_i;
wire signed [`CalcTempBus]          temp_m2_24_4_r;
wire signed [`CalcTempBus]          temp_m2_24_4_i;
wire signed [`CalcTempBus]          temp_m2_24_5_r;
wire signed [`CalcTempBus]          temp_m2_24_5_i;
wire signed [`CalcTempBus]          temp_m2_24_6_r;
wire signed [`CalcTempBus]          temp_m2_24_6_i;
wire signed [`CalcTempBus]          temp_m2_24_7_r;
wire signed [`CalcTempBus]          temp_m2_24_7_i;
wire signed [`CalcTempBus]          temp_m2_24_8_r;
wire signed [`CalcTempBus]          temp_m2_24_8_i;
wire signed [`CalcTempBus]          temp_m2_24_9_r;
wire signed [`CalcTempBus]          temp_m2_24_9_i;
wire signed [`CalcTempBus]          temp_m2_24_10_r;
wire signed [`CalcTempBus]          temp_m2_24_10_i;
wire signed [`CalcTempBus]          temp_m2_24_11_r;
wire signed [`CalcTempBus]          temp_m2_24_11_i;
wire signed [`CalcTempBus]          temp_m2_24_12_r;
wire signed [`CalcTempBus]          temp_m2_24_12_i;
wire signed [`CalcTempBus]          temp_m2_24_13_r;
wire signed [`CalcTempBus]          temp_m2_24_13_i;
wire signed [`CalcTempBus]          temp_m2_24_14_r;
wire signed [`CalcTempBus]          temp_m2_24_14_i;
wire signed [`CalcTempBus]          temp_m2_24_15_r;
wire signed [`CalcTempBus]          temp_m2_24_15_i;
wire signed [`CalcTempBus]          temp_m2_24_16_r;
wire signed [`CalcTempBus]          temp_m2_24_16_i;
wire signed [`CalcTempBus]          temp_m2_24_17_r;
wire signed [`CalcTempBus]          temp_m2_24_17_i;
wire signed [`CalcTempBus]          temp_m2_24_18_r;
wire signed [`CalcTempBus]          temp_m2_24_18_i;
wire signed [`CalcTempBus]          temp_m2_24_19_r;
wire signed [`CalcTempBus]          temp_m2_24_19_i;
wire signed [`CalcTempBus]          temp_m2_24_20_r;
wire signed [`CalcTempBus]          temp_m2_24_20_i;
wire signed [`CalcTempBus]          temp_m2_24_21_r;
wire signed [`CalcTempBus]          temp_m2_24_21_i;
wire signed [`CalcTempBus]          temp_m2_24_22_r;
wire signed [`CalcTempBus]          temp_m2_24_22_i;
wire signed [`CalcTempBus]          temp_m2_24_23_r;
wire signed [`CalcTempBus]          temp_m2_24_23_i;
wire signed [`CalcTempBus]          temp_m2_24_24_r;
wire signed [`CalcTempBus]          temp_m2_24_24_i;
wire signed [`CalcTempBus]          temp_m2_24_25_r;
wire signed [`CalcTempBus]          temp_m2_24_25_i;
wire signed [`CalcTempBus]          temp_m2_24_26_r;
wire signed [`CalcTempBus]          temp_m2_24_26_i;
wire signed [`CalcTempBus]          temp_m2_24_27_r;
wire signed [`CalcTempBus]          temp_m2_24_27_i;
wire signed [`CalcTempBus]          temp_m2_24_28_r;
wire signed [`CalcTempBus]          temp_m2_24_28_i;
wire signed [`CalcTempBus]          temp_m2_24_29_r;
wire signed [`CalcTempBus]          temp_m2_24_29_i;
wire signed [`CalcTempBus]          temp_m2_24_30_r;
wire signed [`CalcTempBus]          temp_m2_24_30_i;
wire signed [`CalcTempBus]          temp_m2_24_31_r;
wire signed [`CalcTempBus]          temp_m2_24_31_i;
wire signed [`CalcTempBus]          temp_m2_24_32_r;
wire signed [`CalcTempBus]          temp_m2_24_32_i;
wire signed [`CalcTempBus]          temp_m2_25_1_r;
wire signed [`CalcTempBus]          temp_m2_25_1_i;
wire signed [`CalcTempBus]          temp_m2_25_2_r;
wire signed [`CalcTempBus]          temp_m2_25_2_i;
wire signed [`CalcTempBus]          temp_m2_25_3_r;
wire signed [`CalcTempBus]          temp_m2_25_3_i;
wire signed [`CalcTempBus]          temp_m2_25_4_r;
wire signed [`CalcTempBus]          temp_m2_25_4_i;
wire signed [`CalcTempBus]          temp_m2_25_5_r;
wire signed [`CalcTempBus]          temp_m2_25_5_i;
wire signed [`CalcTempBus]          temp_m2_25_6_r;
wire signed [`CalcTempBus]          temp_m2_25_6_i;
wire signed [`CalcTempBus]          temp_m2_25_7_r;
wire signed [`CalcTempBus]          temp_m2_25_7_i;
wire signed [`CalcTempBus]          temp_m2_25_8_r;
wire signed [`CalcTempBus]          temp_m2_25_8_i;
wire signed [`CalcTempBus]          temp_m2_25_9_r;
wire signed [`CalcTempBus]          temp_m2_25_9_i;
wire signed [`CalcTempBus]          temp_m2_25_10_r;
wire signed [`CalcTempBus]          temp_m2_25_10_i;
wire signed [`CalcTempBus]          temp_m2_25_11_r;
wire signed [`CalcTempBus]          temp_m2_25_11_i;
wire signed [`CalcTempBus]          temp_m2_25_12_r;
wire signed [`CalcTempBus]          temp_m2_25_12_i;
wire signed [`CalcTempBus]          temp_m2_25_13_r;
wire signed [`CalcTempBus]          temp_m2_25_13_i;
wire signed [`CalcTempBus]          temp_m2_25_14_r;
wire signed [`CalcTempBus]          temp_m2_25_14_i;
wire signed [`CalcTempBus]          temp_m2_25_15_r;
wire signed [`CalcTempBus]          temp_m2_25_15_i;
wire signed [`CalcTempBus]          temp_m2_25_16_r;
wire signed [`CalcTempBus]          temp_m2_25_16_i;
wire signed [`CalcTempBus]          temp_m2_25_17_r;
wire signed [`CalcTempBus]          temp_m2_25_17_i;
wire signed [`CalcTempBus]          temp_m2_25_18_r;
wire signed [`CalcTempBus]          temp_m2_25_18_i;
wire signed [`CalcTempBus]          temp_m2_25_19_r;
wire signed [`CalcTempBus]          temp_m2_25_19_i;
wire signed [`CalcTempBus]          temp_m2_25_20_r;
wire signed [`CalcTempBus]          temp_m2_25_20_i;
wire signed [`CalcTempBus]          temp_m2_25_21_r;
wire signed [`CalcTempBus]          temp_m2_25_21_i;
wire signed [`CalcTempBus]          temp_m2_25_22_r;
wire signed [`CalcTempBus]          temp_m2_25_22_i;
wire signed [`CalcTempBus]          temp_m2_25_23_r;
wire signed [`CalcTempBus]          temp_m2_25_23_i;
wire signed [`CalcTempBus]          temp_m2_25_24_r;
wire signed [`CalcTempBus]          temp_m2_25_24_i;
wire signed [`CalcTempBus]          temp_m2_25_25_r;
wire signed [`CalcTempBus]          temp_m2_25_25_i;
wire signed [`CalcTempBus]          temp_m2_25_26_r;
wire signed [`CalcTempBus]          temp_m2_25_26_i;
wire signed [`CalcTempBus]          temp_m2_25_27_r;
wire signed [`CalcTempBus]          temp_m2_25_27_i;
wire signed [`CalcTempBus]          temp_m2_25_28_r;
wire signed [`CalcTempBus]          temp_m2_25_28_i;
wire signed [`CalcTempBus]          temp_m2_25_29_r;
wire signed [`CalcTempBus]          temp_m2_25_29_i;
wire signed [`CalcTempBus]          temp_m2_25_30_r;
wire signed [`CalcTempBus]          temp_m2_25_30_i;
wire signed [`CalcTempBus]          temp_m2_25_31_r;
wire signed [`CalcTempBus]          temp_m2_25_31_i;
wire signed [`CalcTempBus]          temp_m2_25_32_r;
wire signed [`CalcTempBus]          temp_m2_25_32_i;
wire signed [`CalcTempBus]          temp_m2_26_1_r;
wire signed [`CalcTempBus]          temp_m2_26_1_i;
wire signed [`CalcTempBus]          temp_m2_26_2_r;
wire signed [`CalcTempBus]          temp_m2_26_2_i;
wire signed [`CalcTempBus]          temp_m2_26_3_r;
wire signed [`CalcTempBus]          temp_m2_26_3_i;
wire signed [`CalcTempBus]          temp_m2_26_4_r;
wire signed [`CalcTempBus]          temp_m2_26_4_i;
wire signed [`CalcTempBus]          temp_m2_26_5_r;
wire signed [`CalcTempBus]          temp_m2_26_5_i;
wire signed [`CalcTempBus]          temp_m2_26_6_r;
wire signed [`CalcTempBus]          temp_m2_26_6_i;
wire signed [`CalcTempBus]          temp_m2_26_7_r;
wire signed [`CalcTempBus]          temp_m2_26_7_i;
wire signed [`CalcTempBus]          temp_m2_26_8_r;
wire signed [`CalcTempBus]          temp_m2_26_8_i;
wire signed [`CalcTempBus]          temp_m2_26_9_r;
wire signed [`CalcTempBus]          temp_m2_26_9_i;
wire signed [`CalcTempBus]          temp_m2_26_10_r;
wire signed [`CalcTempBus]          temp_m2_26_10_i;
wire signed [`CalcTempBus]          temp_m2_26_11_r;
wire signed [`CalcTempBus]          temp_m2_26_11_i;
wire signed [`CalcTempBus]          temp_m2_26_12_r;
wire signed [`CalcTempBus]          temp_m2_26_12_i;
wire signed [`CalcTempBus]          temp_m2_26_13_r;
wire signed [`CalcTempBus]          temp_m2_26_13_i;
wire signed [`CalcTempBus]          temp_m2_26_14_r;
wire signed [`CalcTempBus]          temp_m2_26_14_i;
wire signed [`CalcTempBus]          temp_m2_26_15_r;
wire signed [`CalcTempBus]          temp_m2_26_15_i;
wire signed [`CalcTempBus]          temp_m2_26_16_r;
wire signed [`CalcTempBus]          temp_m2_26_16_i;
wire signed [`CalcTempBus]          temp_m2_26_17_r;
wire signed [`CalcTempBus]          temp_m2_26_17_i;
wire signed [`CalcTempBus]          temp_m2_26_18_r;
wire signed [`CalcTempBus]          temp_m2_26_18_i;
wire signed [`CalcTempBus]          temp_m2_26_19_r;
wire signed [`CalcTempBus]          temp_m2_26_19_i;
wire signed [`CalcTempBus]          temp_m2_26_20_r;
wire signed [`CalcTempBus]          temp_m2_26_20_i;
wire signed [`CalcTempBus]          temp_m2_26_21_r;
wire signed [`CalcTempBus]          temp_m2_26_21_i;
wire signed [`CalcTempBus]          temp_m2_26_22_r;
wire signed [`CalcTempBus]          temp_m2_26_22_i;
wire signed [`CalcTempBus]          temp_m2_26_23_r;
wire signed [`CalcTempBus]          temp_m2_26_23_i;
wire signed [`CalcTempBus]          temp_m2_26_24_r;
wire signed [`CalcTempBus]          temp_m2_26_24_i;
wire signed [`CalcTempBus]          temp_m2_26_25_r;
wire signed [`CalcTempBus]          temp_m2_26_25_i;
wire signed [`CalcTempBus]          temp_m2_26_26_r;
wire signed [`CalcTempBus]          temp_m2_26_26_i;
wire signed [`CalcTempBus]          temp_m2_26_27_r;
wire signed [`CalcTempBus]          temp_m2_26_27_i;
wire signed [`CalcTempBus]          temp_m2_26_28_r;
wire signed [`CalcTempBus]          temp_m2_26_28_i;
wire signed [`CalcTempBus]          temp_m2_26_29_r;
wire signed [`CalcTempBus]          temp_m2_26_29_i;
wire signed [`CalcTempBus]          temp_m2_26_30_r;
wire signed [`CalcTempBus]          temp_m2_26_30_i;
wire signed [`CalcTempBus]          temp_m2_26_31_r;
wire signed [`CalcTempBus]          temp_m2_26_31_i;
wire signed [`CalcTempBus]          temp_m2_26_32_r;
wire signed [`CalcTempBus]          temp_m2_26_32_i;
wire signed [`CalcTempBus]          temp_m2_27_1_r;
wire signed [`CalcTempBus]          temp_m2_27_1_i;
wire signed [`CalcTempBus]          temp_m2_27_2_r;
wire signed [`CalcTempBus]          temp_m2_27_2_i;
wire signed [`CalcTempBus]          temp_m2_27_3_r;
wire signed [`CalcTempBus]          temp_m2_27_3_i;
wire signed [`CalcTempBus]          temp_m2_27_4_r;
wire signed [`CalcTempBus]          temp_m2_27_4_i;
wire signed [`CalcTempBus]          temp_m2_27_5_r;
wire signed [`CalcTempBus]          temp_m2_27_5_i;
wire signed [`CalcTempBus]          temp_m2_27_6_r;
wire signed [`CalcTempBus]          temp_m2_27_6_i;
wire signed [`CalcTempBus]          temp_m2_27_7_r;
wire signed [`CalcTempBus]          temp_m2_27_7_i;
wire signed [`CalcTempBus]          temp_m2_27_8_r;
wire signed [`CalcTempBus]          temp_m2_27_8_i;
wire signed [`CalcTempBus]          temp_m2_27_9_r;
wire signed [`CalcTempBus]          temp_m2_27_9_i;
wire signed [`CalcTempBus]          temp_m2_27_10_r;
wire signed [`CalcTempBus]          temp_m2_27_10_i;
wire signed [`CalcTempBus]          temp_m2_27_11_r;
wire signed [`CalcTempBus]          temp_m2_27_11_i;
wire signed [`CalcTempBus]          temp_m2_27_12_r;
wire signed [`CalcTempBus]          temp_m2_27_12_i;
wire signed [`CalcTempBus]          temp_m2_27_13_r;
wire signed [`CalcTempBus]          temp_m2_27_13_i;
wire signed [`CalcTempBus]          temp_m2_27_14_r;
wire signed [`CalcTempBus]          temp_m2_27_14_i;
wire signed [`CalcTempBus]          temp_m2_27_15_r;
wire signed [`CalcTempBus]          temp_m2_27_15_i;
wire signed [`CalcTempBus]          temp_m2_27_16_r;
wire signed [`CalcTempBus]          temp_m2_27_16_i;
wire signed [`CalcTempBus]          temp_m2_27_17_r;
wire signed [`CalcTempBus]          temp_m2_27_17_i;
wire signed [`CalcTempBus]          temp_m2_27_18_r;
wire signed [`CalcTempBus]          temp_m2_27_18_i;
wire signed [`CalcTempBus]          temp_m2_27_19_r;
wire signed [`CalcTempBus]          temp_m2_27_19_i;
wire signed [`CalcTempBus]          temp_m2_27_20_r;
wire signed [`CalcTempBus]          temp_m2_27_20_i;
wire signed [`CalcTempBus]          temp_m2_27_21_r;
wire signed [`CalcTempBus]          temp_m2_27_21_i;
wire signed [`CalcTempBus]          temp_m2_27_22_r;
wire signed [`CalcTempBus]          temp_m2_27_22_i;
wire signed [`CalcTempBus]          temp_m2_27_23_r;
wire signed [`CalcTempBus]          temp_m2_27_23_i;
wire signed [`CalcTempBus]          temp_m2_27_24_r;
wire signed [`CalcTempBus]          temp_m2_27_24_i;
wire signed [`CalcTempBus]          temp_m2_27_25_r;
wire signed [`CalcTempBus]          temp_m2_27_25_i;
wire signed [`CalcTempBus]          temp_m2_27_26_r;
wire signed [`CalcTempBus]          temp_m2_27_26_i;
wire signed [`CalcTempBus]          temp_m2_27_27_r;
wire signed [`CalcTempBus]          temp_m2_27_27_i;
wire signed [`CalcTempBus]          temp_m2_27_28_r;
wire signed [`CalcTempBus]          temp_m2_27_28_i;
wire signed [`CalcTempBus]          temp_m2_27_29_r;
wire signed [`CalcTempBus]          temp_m2_27_29_i;
wire signed [`CalcTempBus]          temp_m2_27_30_r;
wire signed [`CalcTempBus]          temp_m2_27_30_i;
wire signed [`CalcTempBus]          temp_m2_27_31_r;
wire signed [`CalcTempBus]          temp_m2_27_31_i;
wire signed [`CalcTempBus]          temp_m2_27_32_r;
wire signed [`CalcTempBus]          temp_m2_27_32_i;
wire signed [`CalcTempBus]          temp_m2_28_1_r;
wire signed [`CalcTempBus]          temp_m2_28_1_i;
wire signed [`CalcTempBus]          temp_m2_28_2_r;
wire signed [`CalcTempBus]          temp_m2_28_2_i;
wire signed [`CalcTempBus]          temp_m2_28_3_r;
wire signed [`CalcTempBus]          temp_m2_28_3_i;
wire signed [`CalcTempBus]          temp_m2_28_4_r;
wire signed [`CalcTempBus]          temp_m2_28_4_i;
wire signed [`CalcTempBus]          temp_m2_28_5_r;
wire signed [`CalcTempBus]          temp_m2_28_5_i;
wire signed [`CalcTempBus]          temp_m2_28_6_r;
wire signed [`CalcTempBus]          temp_m2_28_6_i;
wire signed [`CalcTempBus]          temp_m2_28_7_r;
wire signed [`CalcTempBus]          temp_m2_28_7_i;
wire signed [`CalcTempBus]          temp_m2_28_8_r;
wire signed [`CalcTempBus]          temp_m2_28_8_i;
wire signed [`CalcTempBus]          temp_m2_28_9_r;
wire signed [`CalcTempBus]          temp_m2_28_9_i;
wire signed [`CalcTempBus]          temp_m2_28_10_r;
wire signed [`CalcTempBus]          temp_m2_28_10_i;
wire signed [`CalcTempBus]          temp_m2_28_11_r;
wire signed [`CalcTempBus]          temp_m2_28_11_i;
wire signed [`CalcTempBus]          temp_m2_28_12_r;
wire signed [`CalcTempBus]          temp_m2_28_12_i;
wire signed [`CalcTempBus]          temp_m2_28_13_r;
wire signed [`CalcTempBus]          temp_m2_28_13_i;
wire signed [`CalcTempBus]          temp_m2_28_14_r;
wire signed [`CalcTempBus]          temp_m2_28_14_i;
wire signed [`CalcTempBus]          temp_m2_28_15_r;
wire signed [`CalcTempBus]          temp_m2_28_15_i;
wire signed [`CalcTempBus]          temp_m2_28_16_r;
wire signed [`CalcTempBus]          temp_m2_28_16_i;
wire signed [`CalcTempBus]          temp_m2_28_17_r;
wire signed [`CalcTempBus]          temp_m2_28_17_i;
wire signed [`CalcTempBus]          temp_m2_28_18_r;
wire signed [`CalcTempBus]          temp_m2_28_18_i;
wire signed [`CalcTempBus]          temp_m2_28_19_r;
wire signed [`CalcTempBus]          temp_m2_28_19_i;
wire signed [`CalcTempBus]          temp_m2_28_20_r;
wire signed [`CalcTempBus]          temp_m2_28_20_i;
wire signed [`CalcTempBus]          temp_m2_28_21_r;
wire signed [`CalcTempBus]          temp_m2_28_21_i;
wire signed [`CalcTempBus]          temp_m2_28_22_r;
wire signed [`CalcTempBus]          temp_m2_28_22_i;
wire signed [`CalcTempBus]          temp_m2_28_23_r;
wire signed [`CalcTempBus]          temp_m2_28_23_i;
wire signed [`CalcTempBus]          temp_m2_28_24_r;
wire signed [`CalcTempBus]          temp_m2_28_24_i;
wire signed [`CalcTempBus]          temp_m2_28_25_r;
wire signed [`CalcTempBus]          temp_m2_28_25_i;
wire signed [`CalcTempBus]          temp_m2_28_26_r;
wire signed [`CalcTempBus]          temp_m2_28_26_i;
wire signed [`CalcTempBus]          temp_m2_28_27_r;
wire signed [`CalcTempBus]          temp_m2_28_27_i;
wire signed [`CalcTempBus]          temp_m2_28_28_r;
wire signed [`CalcTempBus]          temp_m2_28_28_i;
wire signed [`CalcTempBus]          temp_m2_28_29_r;
wire signed [`CalcTempBus]          temp_m2_28_29_i;
wire signed [`CalcTempBus]          temp_m2_28_30_r;
wire signed [`CalcTempBus]          temp_m2_28_30_i;
wire signed [`CalcTempBus]          temp_m2_28_31_r;
wire signed [`CalcTempBus]          temp_m2_28_31_i;
wire signed [`CalcTempBus]          temp_m2_28_32_r;
wire signed [`CalcTempBus]          temp_m2_28_32_i;
wire signed [`CalcTempBus]          temp_m2_29_1_r;
wire signed [`CalcTempBus]          temp_m2_29_1_i;
wire signed [`CalcTempBus]          temp_m2_29_2_r;
wire signed [`CalcTempBus]          temp_m2_29_2_i;
wire signed [`CalcTempBus]          temp_m2_29_3_r;
wire signed [`CalcTempBus]          temp_m2_29_3_i;
wire signed [`CalcTempBus]          temp_m2_29_4_r;
wire signed [`CalcTempBus]          temp_m2_29_4_i;
wire signed [`CalcTempBus]          temp_m2_29_5_r;
wire signed [`CalcTempBus]          temp_m2_29_5_i;
wire signed [`CalcTempBus]          temp_m2_29_6_r;
wire signed [`CalcTempBus]          temp_m2_29_6_i;
wire signed [`CalcTempBus]          temp_m2_29_7_r;
wire signed [`CalcTempBus]          temp_m2_29_7_i;
wire signed [`CalcTempBus]          temp_m2_29_8_r;
wire signed [`CalcTempBus]          temp_m2_29_8_i;
wire signed [`CalcTempBus]          temp_m2_29_9_r;
wire signed [`CalcTempBus]          temp_m2_29_9_i;
wire signed [`CalcTempBus]          temp_m2_29_10_r;
wire signed [`CalcTempBus]          temp_m2_29_10_i;
wire signed [`CalcTempBus]          temp_m2_29_11_r;
wire signed [`CalcTempBus]          temp_m2_29_11_i;
wire signed [`CalcTempBus]          temp_m2_29_12_r;
wire signed [`CalcTempBus]          temp_m2_29_12_i;
wire signed [`CalcTempBus]          temp_m2_29_13_r;
wire signed [`CalcTempBus]          temp_m2_29_13_i;
wire signed [`CalcTempBus]          temp_m2_29_14_r;
wire signed [`CalcTempBus]          temp_m2_29_14_i;
wire signed [`CalcTempBus]          temp_m2_29_15_r;
wire signed [`CalcTempBus]          temp_m2_29_15_i;
wire signed [`CalcTempBus]          temp_m2_29_16_r;
wire signed [`CalcTempBus]          temp_m2_29_16_i;
wire signed [`CalcTempBus]          temp_m2_29_17_r;
wire signed [`CalcTempBus]          temp_m2_29_17_i;
wire signed [`CalcTempBus]          temp_m2_29_18_r;
wire signed [`CalcTempBus]          temp_m2_29_18_i;
wire signed [`CalcTempBus]          temp_m2_29_19_r;
wire signed [`CalcTempBus]          temp_m2_29_19_i;
wire signed [`CalcTempBus]          temp_m2_29_20_r;
wire signed [`CalcTempBus]          temp_m2_29_20_i;
wire signed [`CalcTempBus]          temp_m2_29_21_r;
wire signed [`CalcTempBus]          temp_m2_29_21_i;
wire signed [`CalcTempBus]          temp_m2_29_22_r;
wire signed [`CalcTempBus]          temp_m2_29_22_i;
wire signed [`CalcTempBus]          temp_m2_29_23_r;
wire signed [`CalcTempBus]          temp_m2_29_23_i;
wire signed [`CalcTempBus]          temp_m2_29_24_r;
wire signed [`CalcTempBus]          temp_m2_29_24_i;
wire signed [`CalcTempBus]          temp_m2_29_25_r;
wire signed [`CalcTempBus]          temp_m2_29_25_i;
wire signed [`CalcTempBus]          temp_m2_29_26_r;
wire signed [`CalcTempBus]          temp_m2_29_26_i;
wire signed [`CalcTempBus]          temp_m2_29_27_r;
wire signed [`CalcTempBus]          temp_m2_29_27_i;
wire signed [`CalcTempBus]          temp_m2_29_28_r;
wire signed [`CalcTempBus]          temp_m2_29_28_i;
wire signed [`CalcTempBus]          temp_m2_29_29_r;
wire signed [`CalcTempBus]          temp_m2_29_29_i;
wire signed [`CalcTempBus]          temp_m2_29_30_r;
wire signed [`CalcTempBus]          temp_m2_29_30_i;
wire signed [`CalcTempBus]          temp_m2_29_31_r;
wire signed [`CalcTempBus]          temp_m2_29_31_i;
wire signed [`CalcTempBus]          temp_m2_29_32_r;
wire signed [`CalcTempBus]          temp_m2_29_32_i;
wire signed [`CalcTempBus]          temp_m2_30_1_r;
wire signed [`CalcTempBus]          temp_m2_30_1_i;
wire signed [`CalcTempBus]          temp_m2_30_2_r;
wire signed [`CalcTempBus]          temp_m2_30_2_i;
wire signed [`CalcTempBus]          temp_m2_30_3_r;
wire signed [`CalcTempBus]          temp_m2_30_3_i;
wire signed [`CalcTempBus]          temp_m2_30_4_r;
wire signed [`CalcTempBus]          temp_m2_30_4_i;
wire signed [`CalcTempBus]          temp_m2_30_5_r;
wire signed [`CalcTempBus]          temp_m2_30_5_i;
wire signed [`CalcTempBus]          temp_m2_30_6_r;
wire signed [`CalcTempBus]          temp_m2_30_6_i;
wire signed [`CalcTempBus]          temp_m2_30_7_r;
wire signed [`CalcTempBus]          temp_m2_30_7_i;
wire signed [`CalcTempBus]          temp_m2_30_8_r;
wire signed [`CalcTempBus]          temp_m2_30_8_i;
wire signed [`CalcTempBus]          temp_m2_30_9_r;
wire signed [`CalcTempBus]          temp_m2_30_9_i;
wire signed [`CalcTempBus]          temp_m2_30_10_r;
wire signed [`CalcTempBus]          temp_m2_30_10_i;
wire signed [`CalcTempBus]          temp_m2_30_11_r;
wire signed [`CalcTempBus]          temp_m2_30_11_i;
wire signed [`CalcTempBus]          temp_m2_30_12_r;
wire signed [`CalcTempBus]          temp_m2_30_12_i;
wire signed [`CalcTempBus]          temp_m2_30_13_r;
wire signed [`CalcTempBus]          temp_m2_30_13_i;
wire signed [`CalcTempBus]          temp_m2_30_14_r;
wire signed [`CalcTempBus]          temp_m2_30_14_i;
wire signed [`CalcTempBus]          temp_m2_30_15_r;
wire signed [`CalcTempBus]          temp_m2_30_15_i;
wire signed [`CalcTempBus]          temp_m2_30_16_r;
wire signed [`CalcTempBus]          temp_m2_30_16_i;
wire signed [`CalcTempBus]          temp_m2_30_17_r;
wire signed [`CalcTempBus]          temp_m2_30_17_i;
wire signed [`CalcTempBus]          temp_m2_30_18_r;
wire signed [`CalcTempBus]          temp_m2_30_18_i;
wire signed [`CalcTempBus]          temp_m2_30_19_r;
wire signed [`CalcTempBus]          temp_m2_30_19_i;
wire signed [`CalcTempBus]          temp_m2_30_20_r;
wire signed [`CalcTempBus]          temp_m2_30_20_i;
wire signed [`CalcTempBus]          temp_m2_30_21_r;
wire signed [`CalcTempBus]          temp_m2_30_21_i;
wire signed [`CalcTempBus]          temp_m2_30_22_r;
wire signed [`CalcTempBus]          temp_m2_30_22_i;
wire signed [`CalcTempBus]          temp_m2_30_23_r;
wire signed [`CalcTempBus]          temp_m2_30_23_i;
wire signed [`CalcTempBus]          temp_m2_30_24_r;
wire signed [`CalcTempBus]          temp_m2_30_24_i;
wire signed [`CalcTempBus]          temp_m2_30_25_r;
wire signed [`CalcTempBus]          temp_m2_30_25_i;
wire signed [`CalcTempBus]          temp_m2_30_26_r;
wire signed [`CalcTempBus]          temp_m2_30_26_i;
wire signed [`CalcTempBus]          temp_m2_30_27_r;
wire signed [`CalcTempBus]          temp_m2_30_27_i;
wire signed [`CalcTempBus]          temp_m2_30_28_r;
wire signed [`CalcTempBus]          temp_m2_30_28_i;
wire signed [`CalcTempBus]          temp_m2_30_29_r;
wire signed [`CalcTempBus]          temp_m2_30_29_i;
wire signed [`CalcTempBus]          temp_m2_30_30_r;
wire signed [`CalcTempBus]          temp_m2_30_30_i;
wire signed [`CalcTempBus]          temp_m2_30_31_r;
wire signed [`CalcTempBus]          temp_m2_30_31_i;
wire signed [`CalcTempBus]          temp_m2_30_32_r;
wire signed [`CalcTempBus]          temp_m2_30_32_i;
wire signed [`CalcTempBus]          temp_m2_31_1_r;
wire signed [`CalcTempBus]          temp_m2_31_1_i;
wire signed [`CalcTempBus]          temp_m2_31_2_r;
wire signed [`CalcTempBus]          temp_m2_31_2_i;
wire signed [`CalcTempBus]          temp_m2_31_3_r;
wire signed [`CalcTempBus]          temp_m2_31_3_i;
wire signed [`CalcTempBus]          temp_m2_31_4_r;
wire signed [`CalcTempBus]          temp_m2_31_4_i;
wire signed [`CalcTempBus]          temp_m2_31_5_r;
wire signed [`CalcTempBus]          temp_m2_31_5_i;
wire signed [`CalcTempBus]          temp_m2_31_6_r;
wire signed [`CalcTempBus]          temp_m2_31_6_i;
wire signed [`CalcTempBus]          temp_m2_31_7_r;
wire signed [`CalcTempBus]          temp_m2_31_7_i;
wire signed [`CalcTempBus]          temp_m2_31_8_r;
wire signed [`CalcTempBus]          temp_m2_31_8_i;
wire signed [`CalcTempBus]          temp_m2_31_9_r;
wire signed [`CalcTempBus]          temp_m2_31_9_i;
wire signed [`CalcTempBus]          temp_m2_31_10_r;
wire signed [`CalcTempBus]          temp_m2_31_10_i;
wire signed [`CalcTempBus]          temp_m2_31_11_r;
wire signed [`CalcTempBus]          temp_m2_31_11_i;
wire signed [`CalcTempBus]          temp_m2_31_12_r;
wire signed [`CalcTempBus]          temp_m2_31_12_i;
wire signed [`CalcTempBus]          temp_m2_31_13_r;
wire signed [`CalcTempBus]          temp_m2_31_13_i;
wire signed [`CalcTempBus]          temp_m2_31_14_r;
wire signed [`CalcTempBus]          temp_m2_31_14_i;
wire signed [`CalcTempBus]          temp_m2_31_15_r;
wire signed [`CalcTempBus]          temp_m2_31_15_i;
wire signed [`CalcTempBus]          temp_m2_31_16_r;
wire signed [`CalcTempBus]          temp_m2_31_16_i;
wire signed [`CalcTempBus]          temp_m2_31_17_r;
wire signed [`CalcTempBus]          temp_m2_31_17_i;
wire signed [`CalcTempBus]          temp_m2_31_18_r;
wire signed [`CalcTempBus]          temp_m2_31_18_i;
wire signed [`CalcTempBus]          temp_m2_31_19_r;
wire signed [`CalcTempBus]          temp_m2_31_19_i;
wire signed [`CalcTempBus]          temp_m2_31_20_r;
wire signed [`CalcTempBus]          temp_m2_31_20_i;
wire signed [`CalcTempBus]          temp_m2_31_21_r;
wire signed [`CalcTempBus]          temp_m2_31_21_i;
wire signed [`CalcTempBus]          temp_m2_31_22_r;
wire signed [`CalcTempBus]          temp_m2_31_22_i;
wire signed [`CalcTempBus]          temp_m2_31_23_r;
wire signed [`CalcTempBus]          temp_m2_31_23_i;
wire signed [`CalcTempBus]          temp_m2_31_24_r;
wire signed [`CalcTempBus]          temp_m2_31_24_i;
wire signed [`CalcTempBus]          temp_m2_31_25_r;
wire signed [`CalcTempBus]          temp_m2_31_25_i;
wire signed [`CalcTempBus]          temp_m2_31_26_r;
wire signed [`CalcTempBus]          temp_m2_31_26_i;
wire signed [`CalcTempBus]          temp_m2_31_27_r;
wire signed [`CalcTempBus]          temp_m2_31_27_i;
wire signed [`CalcTempBus]          temp_m2_31_28_r;
wire signed [`CalcTempBus]          temp_m2_31_28_i;
wire signed [`CalcTempBus]          temp_m2_31_29_r;
wire signed [`CalcTempBus]          temp_m2_31_29_i;
wire signed [`CalcTempBus]          temp_m2_31_30_r;
wire signed [`CalcTempBus]          temp_m2_31_30_i;
wire signed [`CalcTempBus]          temp_m2_31_31_r;
wire signed [`CalcTempBus]          temp_m2_31_31_i;
wire signed [`CalcTempBus]          temp_m2_31_32_r;
wire signed [`CalcTempBus]          temp_m2_31_32_i;
wire signed [`CalcTempBus]          temp_m2_32_1_r;
wire signed [`CalcTempBus]          temp_m2_32_1_i;
wire signed [`CalcTempBus]          temp_m2_32_2_r;
wire signed [`CalcTempBus]          temp_m2_32_2_i;
wire signed [`CalcTempBus]          temp_m2_32_3_r;
wire signed [`CalcTempBus]          temp_m2_32_3_i;
wire signed [`CalcTempBus]          temp_m2_32_4_r;
wire signed [`CalcTempBus]          temp_m2_32_4_i;
wire signed [`CalcTempBus]          temp_m2_32_5_r;
wire signed [`CalcTempBus]          temp_m2_32_5_i;
wire signed [`CalcTempBus]          temp_m2_32_6_r;
wire signed [`CalcTempBus]          temp_m2_32_6_i;
wire signed [`CalcTempBus]          temp_m2_32_7_r;
wire signed [`CalcTempBus]          temp_m2_32_7_i;
wire signed [`CalcTempBus]          temp_m2_32_8_r;
wire signed [`CalcTempBus]          temp_m2_32_8_i;
wire signed [`CalcTempBus]          temp_m2_32_9_r;
wire signed [`CalcTempBus]          temp_m2_32_9_i;
wire signed [`CalcTempBus]          temp_m2_32_10_r;
wire signed [`CalcTempBus]          temp_m2_32_10_i;
wire signed [`CalcTempBus]          temp_m2_32_11_r;
wire signed [`CalcTempBus]          temp_m2_32_11_i;
wire signed [`CalcTempBus]          temp_m2_32_12_r;
wire signed [`CalcTempBus]          temp_m2_32_12_i;
wire signed [`CalcTempBus]          temp_m2_32_13_r;
wire signed [`CalcTempBus]          temp_m2_32_13_i;
wire signed [`CalcTempBus]          temp_m2_32_14_r;
wire signed [`CalcTempBus]          temp_m2_32_14_i;
wire signed [`CalcTempBus]          temp_m2_32_15_r;
wire signed [`CalcTempBus]          temp_m2_32_15_i;
wire signed [`CalcTempBus]          temp_m2_32_16_r;
wire signed [`CalcTempBus]          temp_m2_32_16_i;
wire signed [`CalcTempBus]          temp_m2_32_17_r;
wire signed [`CalcTempBus]          temp_m2_32_17_i;
wire signed [`CalcTempBus]          temp_m2_32_18_r;
wire signed [`CalcTempBus]          temp_m2_32_18_i;
wire signed [`CalcTempBus]          temp_m2_32_19_r;
wire signed [`CalcTempBus]          temp_m2_32_19_i;
wire signed [`CalcTempBus]          temp_m2_32_20_r;
wire signed [`CalcTempBus]          temp_m2_32_20_i;
wire signed [`CalcTempBus]          temp_m2_32_21_r;
wire signed [`CalcTempBus]          temp_m2_32_21_i;
wire signed [`CalcTempBus]          temp_m2_32_22_r;
wire signed [`CalcTempBus]          temp_m2_32_22_i;
wire signed [`CalcTempBus]          temp_m2_32_23_r;
wire signed [`CalcTempBus]          temp_m2_32_23_i;
wire signed [`CalcTempBus]          temp_m2_32_24_r;
wire signed [`CalcTempBus]          temp_m2_32_24_i;
wire signed [`CalcTempBus]          temp_m2_32_25_r;
wire signed [`CalcTempBus]          temp_m2_32_25_i;
wire signed [`CalcTempBus]          temp_m2_32_26_r;
wire signed [`CalcTempBus]          temp_m2_32_26_i;
wire signed [`CalcTempBus]          temp_m2_32_27_r;
wire signed [`CalcTempBus]          temp_m2_32_27_i;
wire signed [`CalcTempBus]          temp_m2_32_28_r;
wire signed [`CalcTempBus]          temp_m2_32_28_i;
wire signed [`CalcTempBus]          temp_m2_32_29_r;
wire signed [`CalcTempBus]          temp_m2_32_29_i;
wire signed [`CalcTempBus]          temp_m2_32_30_r;
wire signed [`CalcTempBus]          temp_m2_32_30_i;
wire signed [`CalcTempBus]          temp_m2_32_31_r;
wire signed [`CalcTempBus]          temp_m2_32_31_i;
wire signed [`CalcTempBus]          temp_m2_32_32_r;
wire signed [`CalcTempBus]          temp_m2_32_32_i;
wire signed [`CalcTempBus]          temp_m3_1_1_r;
wire signed [`CalcTempBus]          temp_m3_1_1_i;
wire signed [`CalcTempBus]          temp_m3_1_2_r;
wire signed [`CalcTempBus]          temp_m3_1_2_i;
wire signed [`CalcTempBus]          temp_m3_1_3_r;
wire signed [`CalcTempBus]          temp_m3_1_3_i;
wire signed [`CalcTempBus]          temp_m3_1_4_r;
wire signed [`CalcTempBus]          temp_m3_1_4_i;
wire signed [`CalcTempBus]          temp_m3_1_5_r;
wire signed [`CalcTempBus]          temp_m3_1_5_i;
wire signed [`CalcTempBus]          temp_m3_1_6_r;
wire signed [`CalcTempBus]          temp_m3_1_6_i;
wire signed [`CalcTempBus]          temp_m3_1_7_r;
wire signed [`CalcTempBus]          temp_m3_1_7_i;
wire signed [`CalcTempBus]          temp_m3_1_8_r;
wire signed [`CalcTempBus]          temp_m3_1_8_i;
wire signed [`CalcTempBus]          temp_m3_1_9_r;
wire signed [`CalcTempBus]          temp_m3_1_9_i;
wire signed [`CalcTempBus]          temp_m3_1_10_r;
wire signed [`CalcTempBus]          temp_m3_1_10_i;
wire signed [`CalcTempBus]          temp_m3_1_11_r;
wire signed [`CalcTempBus]          temp_m3_1_11_i;
wire signed [`CalcTempBus]          temp_m3_1_12_r;
wire signed [`CalcTempBus]          temp_m3_1_12_i;
wire signed [`CalcTempBus]          temp_m3_1_13_r;
wire signed [`CalcTempBus]          temp_m3_1_13_i;
wire signed [`CalcTempBus]          temp_m3_1_14_r;
wire signed [`CalcTempBus]          temp_m3_1_14_i;
wire signed [`CalcTempBus]          temp_m3_1_15_r;
wire signed [`CalcTempBus]          temp_m3_1_15_i;
wire signed [`CalcTempBus]          temp_m3_1_16_r;
wire signed [`CalcTempBus]          temp_m3_1_16_i;
wire signed [`CalcTempBus]          temp_m3_1_17_r;
wire signed [`CalcTempBus]          temp_m3_1_17_i;
wire signed [`CalcTempBus]          temp_m3_1_18_r;
wire signed [`CalcTempBus]          temp_m3_1_18_i;
wire signed [`CalcTempBus]          temp_m3_1_19_r;
wire signed [`CalcTempBus]          temp_m3_1_19_i;
wire signed [`CalcTempBus]          temp_m3_1_20_r;
wire signed [`CalcTempBus]          temp_m3_1_20_i;
wire signed [`CalcTempBus]          temp_m3_1_21_r;
wire signed [`CalcTempBus]          temp_m3_1_21_i;
wire signed [`CalcTempBus]          temp_m3_1_22_r;
wire signed [`CalcTempBus]          temp_m3_1_22_i;
wire signed [`CalcTempBus]          temp_m3_1_23_r;
wire signed [`CalcTempBus]          temp_m3_1_23_i;
wire signed [`CalcTempBus]          temp_m3_1_24_r;
wire signed [`CalcTempBus]          temp_m3_1_24_i;
wire signed [`CalcTempBus]          temp_m3_1_25_r;
wire signed [`CalcTempBus]          temp_m3_1_25_i;
wire signed [`CalcTempBus]          temp_m3_1_26_r;
wire signed [`CalcTempBus]          temp_m3_1_26_i;
wire signed [`CalcTempBus]          temp_m3_1_27_r;
wire signed [`CalcTempBus]          temp_m3_1_27_i;
wire signed [`CalcTempBus]          temp_m3_1_28_r;
wire signed [`CalcTempBus]          temp_m3_1_28_i;
wire signed [`CalcTempBus]          temp_m3_1_29_r;
wire signed [`CalcTempBus]          temp_m3_1_29_i;
wire signed [`CalcTempBus]          temp_m3_1_30_r;
wire signed [`CalcTempBus]          temp_m3_1_30_i;
wire signed [`CalcTempBus]          temp_m3_1_31_r;
wire signed [`CalcTempBus]          temp_m3_1_31_i;
wire signed [`CalcTempBus]          temp_m3_1_32_r;
wire signed [`CalcTempBus]          temp_m3_1_32_i;
wire signed [`CalcTempBus]          temp_m3_2_1_r;
wire signed [`CalcTempBus]          temp_m3_2_1_i;
wire signed [`CalcTempBus]          temp_m3_2_2_r;
wire signed [`CalcTempBus]          temp_m3_2_2_i;
wire signed [`CalcTempBus]          temp_m3_2_3_r;
wire signed [`CalcTempBus]          temp_m3_2_3_i;
wire signed [`CalcTempBus]          temp_m3_2_4_r;
wire signed [`CalcTempBus]          temp_m3_2_4_i;
wire signed [`CalcTempBus]          temp_m3_2_5_r;
wire signed [`CalcTempBus]          temp_m3_2_5_i;
wire signed [`CalcTempBus]          temp_m3_2_6_r;
wire signed [`CalcTempBus]          temp_m3_2_6_i;
wire signed [`CalcTempBus]          temp_m3_2_7_r;
wire signed [`CalcTempBus]          temp_m3_2_7_i;
wire signed [`CalcTempBus]          temp_m3_2_8_r;
wire signed [`CalcTempBus]          temp_m3_2_8_i;
wire signed [`CalcTempBus]          temp_m3_2_9_r;
wire signed [`CalcTempBus]          temp_m3_2_9_i;
wire signed [`CalcTempBus]          temp_m3_2_10_r;
wire signed [`CalcTempBus]          temp_m3_2_10_i;
wire signed [`CalcTempBus]          temp_m3_2_11_r;
wire signed [`CalcTempBus]          temp_m3_2_11_i;
wire signed [`CalcTempBus]          temp_m3_2_12_r;
wire signed [`CalcTempBus]          temp_m3_2_12_i;
wire signed [`CalcTempBus]          temp_m3_2_13_r;
wire signed [`CalcTempBus]          temp_m3_2_13_i;
wire signed [`CalcTempBus]          temp_m3_2_14_r;
wire signed [`CalcTempBus]          temp_m3_2_14_i;
wire signed [`CalcTempBus]          temp_m3_2_15_r;
wire signed [`CalcTempBus]          temp_m3_2_15_i;
wire signed [`CalcTempBus]          temp_m3_2_16_r;
wire signed [`CalcTempBus]          temp_m3_2_16_i;
wire signed [`CalcTempBus]          temp_m3_2_17_r;
wire signed [`CalcTempBus]          temp_m3_2_17_i;
wire signed [`CalcTempBus]          temp_m3_2_18_r;
wire signed [`CalcTempBus]          temp_m3_2_18_i;
wire signed [`CalcTempBus]          temp_m3_2_19_r;
wire signed [`CalcTempBus]          temp_m3_2_19_i;
wire signed [`CalcTempBus]          temp_m3_2_20_r;
wire signed [`CalcTempBus]          temp_m3_2_20_i;
wire signed [`CalcTempBus]          temp_m3_2_21_r;
wire signed [`CalcTempBus]          temp_m3_2_21_i;
wire signed [`CalcTempBus]          temp_m3_2_22_r;
wire signed [`CalcTempBus]          temp_m3_2_22_i;
wire signed [`CalcTempBus]          temp_m3_2_23_r;
wire signed [`CalcTempBus]          temp_m3_2_23_i;
wire signed [`CalcTempBus]          temp_m3_2_24_r;
wire signed [`CalcTempBus]          temp_m3_2_24_i;
wire signed [`CalcTempBus]          temp_m3_2_25_r;
wire signed [`CalcTempBus]          temp_m3_2_25_i;
wire signed [`CalcTempBus]          temp_m3_2_26_r;
wire signed [`CalcTempBus]          temp_m3_2_26_i;
wire signed [`CalcTempBus]          temp_m3_2_27_r;
wire signed [`CalcTempBus]          temp_m3_2_27_i;
wire signed [`CalcTempBus]          temp_m3_2_28_r;
wire signed [`CalcTempBus]          temp_m3_2_28_i;
wire signed [`CalcTempBus]          temp_m3_2_29_r;
wire signed [`CalcTempBus]          temp_m3_2_29_i;
wire signed [`CalcTempBus]          temp_m3_2_30_r;
wire signed [`CalcTempBus]          temp_m3_2_30_i;
wire signed [`CalcTempBus]          temp_m3_2_31_r;
wire signed [`CalcTempBus]          temp_m3_2_31_i;
wire signed [`CalcTempBus]          temp_m3_2_32_r;
wire signed [`CalcTempBus]          temp_m3_2_32_i;
wire signed [`CalcTempBus]          temp_m3_3_1_r;
wire signed [`CalcTempBus]          temp_m3_3_1_i;
wire signed [`CalcTempBus]          temp_m3_3_2_r;
wire signed [`CalcTempBus]          temp_m3_3_2_i;
wire signed [`CalcTempBus]          temp_m3_3_3_r;
wire signed [`CalcTempBus]          temp_m3_3_3_i;
wire signed [`CalcTempBus]          temp_m3_3_4_r;
wire signed [`CalcTempBus]          temp_m3_3_4_i;
wire signed [`CalcTempBus]          temp_m3_3_5_r;
wire signed [`CalcTempBus]          temp_m3_3_5_i;
wire signed [`CalcTempBus]          temp_m3_3_6_r;
wire signed [`CalcTempBus]          temp_m3_3_6_i;
wire signed [`CalcTempBus]          temp_m3_3_7_r;
wire signed [`CalcTempBus]          temp_m3_3_7_i;
wire signed [`CalcTempBus]          temp_m3_3_8_r;
wire signed [`CalcTempBus]          temp_m3_3_8_i;
wire signed [`CalcTempBus]          temp_m3_3_9_r;
wire signed [`CalcTempBus]          temp_m3_3_9_i;
wire signed [`CalcTempBus]          temp_m3_3_10_r;
wire signed [`CalcTempBus]          temp_m3_3_10_i;
wire signed [`CalcTempBus]          temp_m3_3_11_r;
wire signed [`CalcTempBus]          temp_m3_3_11_i;
wire signed [`CalcTempBus]          temp_m3_3_12_r;
wire signed [`CalcTempBus]          temp_m3_3_12_i;
wire signed [`CalcTempBus]          temp_m3_3_13_r;
wire signed [`CalcTempBus]          temp_m3_3_13_i;
wire signed [`CalcTempBus]          temp_m3_3_14_r;
wire signed [`CalcTempBus]          temp_m3_3_14_i;
wire signed [`CalcTempBus]          temp_m3_3_15_r;
wire signed [`CalcTempBus]          temp_m3_3_15_i;
wire signed [`CalcTempBus]          temp_m3_3_16_r;
wire signed [`CalcTempBus]          temp_m3_3_16_i;
wire signed [`CalcTempBus]          temp_m3_3_17_r;
wire signed [`CalcTempBus]          temp_m3_3_17_i;
wire signed [`CalcTempBus]          temp_m3_3_18_r;
wire signed [`CalcTempBus]          temp_m3_3_18_i;
wire signed [`CalcTempBus]          temp_m3_3_19_r;
wire signed [`CalcTempBus]          temp_m3_3_19_i;
wire signed [`CalcTempBus]          temp_m3_3_20_r;
wire signed [`CalcTempBus]          temp_m3_3_20_i;
wire signed [`CalcTempBus]          temp_m3_3_21_r;
wire signed [`CalcTempBus]          temp_m3_3_21_i;
wire signed [`CalcTempBus]          temp_m3_3_22_r;
wire signed [`CalcTempBus]          temp_m3_3_22_i;
wire signed [`CalcTempBus]          temp_m3_3_23_r;
wire signed [`CalcTempBus]          temp_m3_3_23_i;
wire signed [`CalcTempBus]          temp_m3_3_24_r;
wire signed [`CalcTempBus]          temp_m3_3_24_i;
wire signed [`CalcTempBus]          temp_m3_3_25_r;
wire signed [`CalcTempBus]          temp_m3_3_25_i;
wire signed [`CalcTempBus]          temp_m3_3_26_r;
wire signed [`CalcTempBus]          temp_m3_3_26_i;
wire signed [`CalcTempBus]          temp_m3_3_27_r;
wire signed [`CalcTempBus]          temp_m3_3_27_i;
wire signed [`CalcTempBus]          temp_m3_3_28_r;
wire signed [`CalcTempBus]          temp_m3_3_28_i;
wire signed [`CalcTempBus]          temp_m3_3_29_r;
wire signed [`CalcTempBus]          temp_m3_3_29_i;
wire signed [`CalcTempBus]          temp_m3_3_30_r;
wire signed [`CalcTempBus]          temp_m3_3_30_i;
wire signed [`CalcTempBus]          temp_m3_3_31_r;
wire signed [`CalcTempBus]          temp_m3_3_31_i;
wire signed [`CalcTempBus]          temp_m3_3_32_r;
wire signed [`CalcTempBus]          temp_m3_3_32_i;
wire signed [`CalcTempBus]          temp_m3_4_1_r;
wire signed [`CalcTempBus]          temp_m3_4_1_i;
wire signed [`CalcTempBus]          temp_m3_4_2_r;
wire signed [`CalcTempBus]          temp_m3_4_2_i;
wire signed [`CalcTempBus]          temp_m3_4_3_r;
wire signed [`CalcTempBus]          temp_m3_4_3_i;
wire signed [`CalcTempBus]          temp_m3_4_4_r;
wire signed [`CalcTempBus]          temp_m3_4_4_i;
wire signed [`CalcTempBus]          temp_m3_4_5_r;
wire signed [`CalcTempBus]          temp_m3_4_5_i;
wire signed [`CalcTempBus]          temp_m3_4_6_r;
wire signed [`CalcTempBus]          temp_m3_4_6_i;
wire signed [`CalcTempBus]          temp_m3_4_7_r;
wire signed [`CalcTempBus]          temp_m3_4_7_i;
wire signed [`CalcTempBus]          temp_m3_4_8_r;
wire signed [`CalcTempBus]          temp_m3_4_8_i;
wire signed [`CalcTempBus]          temp_m3_4_9_r;
wire signed [`CalcTempBus]          temp_m3_4_9_i;
wire signed [`CalcTempBus]          temp_m3_4_10_r;
wire signed [`CalcTempBus]          temp_m3_4_10_i;
wire signed [`CalcTempBus]          temp_m3_4_11_r;
wire signed [`CalcTempBus]          temp_m3_4_11_i;
wire signed [`CalcTempBus]          temp_m3_4_12_r;
wire signed [`CalcTempBus]          temp_m3_4_12_i;
wire signed [`CalcTempBus]          temp_m3_4_13_r;
wire signed [`CalcTempBus]          temp_m3_4_13_i;
wire signed [`CalcTempBus]          temp_m3_4_14_r;
wire signed [`CalcTempBus]          temp_m3_4_14_i;
wire signed [`CalcTempBus]          temp_m3_4_15_r;
wire signed [`CalcTempBus]          temp_m3_4_15_i;
wire signed [`CalcTempBus]          temp_m3_4_16_r;
wire signed [`CalcTempBus]          temp_m3_4_16_i;
wire signed [`CalcTempBus]          temp_m3_4_17_r;
wire signed [`CalcTempBus]          temp_m3_4_17_i;
wire signed [`CalcTempBus]          temp_m3_4_18_r;
wire signed [`CalcTempBus]          temp_m3_4_18_i;
wire signed [`CalcTempBus]          temp_m3_4_19_r;
wire signed [`CalcTempBus]          temp_m3_4_19_i;
wire signed [`CalcTempBus]          temp_m3_4_20_r;
wire signed [`CalcTempBus]          temp_m3_4_20_i;
wire signed [`CalcTempBus]          temp_m3_4_21_r;
wire signed [`CalcTempBus]          temp_m3_4_21_i;
wire signed [`CalcTempBus]          temp_m3_4_22_r;
wire signed [`CalcTempBus]          temp_m3_4_22_i;
wire signed [`CalcTempBus]          temp_m3_4_23_r;
wire signed [`CalcTempBus]          temp_m3_4_23_i;
wire signed [`CalcTempBus]          temp_m3_4_24_r;
wire signed [`CalcTempBus]          temp_m3_4_24_i;
wire signed [`CalcTempBus]          temp_m3_4_25_r;
wire signed [`CalcTempBus]          temp_m3_4_25_i;
wire signed [`CalcTempBus]          temp_m3_4_26_r;
wire signed [`CalcTempBus]          temp_m3_4_26_i;
wire signed [`CalcTempBus]          temp_m3_4_27_r;
wire signed [`CalcTempBus]          temp_m3_4_27_i;
wire signed [`CalcTempBus]          temp_m3_4_28_r;
wire signed [`CalcTempBus]          temp_m3_4_28_i;
wire signed [`CalcTempBus]          temp_m3_4_29_r;
wire signed [`CalcTempBus]          temp_m3_4_29_i;
wire signed [`CalcTempBus]          temp_m3_4_30_r;
wire signed [`CalcTempBus]          temp_m3_4_30_i;
wire signed [`CalcTempBus]          temp_m3_4_31_r;
wire signed [`CalcTempBus]          temp_m3_4_31_i;
wire signed [`CalcTempBus]          temp_m3_4_32_r;
wire signed [`CalcTempBus]          temp_m3_4_32_i;
wire signed [`CalcTempBus]          temp_m3_5_1_r;
wire signed [`CalcTempBus]          temp_m3_5_1_i;
wire signed [`CalcTempBus]          temp_m3_5_2_r;
wire signed [`CalcTempBus]          temp_m3_5_2_i;
wire signed [`CalcTempBus]          temp_m3_5_3_r;
wire signed [`CalcTempBus]          temp_m3_5_3_i;
wire signed [`CalcTempBus]          temp_m3_5_4_r;
wire signed [`CalcTempBus]          temp_m3_5_4_i;
wire signed [`CalcTempBus]          temp_m3_5_5_r;
wire signed [`CalcTempBus]          temp_m3_5_5_i;
wire signed [`CalcTempBus]          temp_m3_5_6_r;
wire signed [`CalcTempBus]          temp_m3_5_6_i;
wire signed [`CalcTempBus]          temp_m3_5_7_r;
wire signed [`CalcTempBus]          temp_m3_5_7_i;
wire signed [`CalcTempBus]          temp_m3_5_8_r;
wire signed [`CalcTempBus]          temp_m3_5_8_i;
wire signed [`CalcTempBus]          temp_m3_5_9_r;
wire signed [`CalcTempBus]          temp_m3_5_9_i;
wire signed [`CalcTempBus]          temp_m3_5_10_r;
wire signed [`CalcTempBus]          temp_m3_5_10_i;
wire signed [`CalcTempBus]          temp_m3_5_11_r;
wire signed [`CalcTempBus]          temp_m3_5_11_i;
wire signed [`CalcTempBus]          temp_m3_5_12_r;
wire signed [`CalcTempBus]          temp_m3_5_12_i;
wire signed [`CalcTempBus]          temp_m3_5_13_r;
wire signed [`CalcTempBus]          temp_m3_5_13_i;
wire signed [`CalcTempBus]          temp_m3_5_14_r;
wire signed [`CalcTempBus]          temp_m3_5_14_i;
wire signed [`CalcTempBus]          temp_m3_5_15_r;
wire signed [`CalcTempBus]          temp_m3_5_15_i;
wire signed [`CalcTempBus]          temp_m3_5_16_r;
wire signed [`CalcTempBus]          temp_m3_5_16_i;
wire signed [`CalcTempBus]          temp_m3_5_17_r;
wire signed [`CalcTempBus]          temp_m3_5_17_i;
wire signed [`CalcTempBus]          temp_m3_5_18_r;
wire signed [`CalcTempBus]          temp_m3_5_18_i;
wire signed [`CalcTempBus]          temp_m3_5_19_r;
wire signed [`CalcTempBus]          temp_m3_5_19_i;
wire signed [`CalcTempBus]          temp_m3_5_20_r;
wire signed [`CalcTempBus]          temp_m3_5_20_i;
wire signed [`CalcTempBus]          temp_m3_5_21_r;
wire signed [`CalcTempBus]          temp_m3_5_21_i;
wire signed [`CalcTempBus]          temp_m3_5_22_r;
wire signed [`CalcTempBus]          temp_m3_5_22_i;
wire signed [`CalcTempBus]          temp_m3_5_23_r;
wire signed [`CalcTempBus]          temp_m3_5_23_i;
wire signed [`CalcTempBus]          temp_m3_5_24_r;
wire signed [`CalcTempBus]          temp_m3_5_24_i;
wire signed [`CalcTempBus]          temp_m3_5_25_r;
wire signed [`CalcTempBus]          temp_m3_5_25_i;
wire signed [`CalcTempBus]          temp_m3_5_26_r;
wire signed [`CalcTempBus]          temp_m3_5_26_i;
wire signed [`CalcTempBus]          temp_m3_5_27_r;
wire signed [`CalcTempBus]          temp_m3_5_27_i;
wire signed [`CalcTempBus]          temp_m3_5_28_r;
wire signed [`CalcTempBus]          temp_m3_5_28_i;
wire signed [`CalcTempBus]          temp_m3_5_29_r;
wire signed [`CalcTempBus]          temp_m3_5_29_i;
wire signed [`CalcTempBus]          temp_m3_5_30_r;
wire signed [`CalcTempBus]          temp_m3_5_30_i;
wire signed [`CalcTempBus]          temp_m3_5_31_r;
wire signed [`CalcTempBus]          temp_m3_5_31_i;
wire signed [`CalcTempBus]          temp_m3_5_32_r;
wire signed [`CalcTempBus]          temp_m3_5_32_i;
wire signed [`CalcTempBus]          temp_m3_6_1_r;
wire signed [`CalcTempBus]          temp_m3_6_1_i;
wire signed [`CalcTempBus]          temp_m3_6_2_r;
wire signed [`CalcTempBus]          temp_m3_6_2_i;
wire signed [`CalcTempBus]          temp_m3_6_3_r;
wire signed [`CalcTempBus]          temp_m3_6_3_i;
wire signed [`CalcTempBus]          temp_m3_6_4_r;
wire signed [`CalcTempBus]          temp_m3_6_4_i;
wire signed [`CalcTempBus]          temp_m3_6_5_r;
wire signed [`CalcTempBus]          temp_m3_6_5_i;
wire signed [`CalcTempBus]          temp_m3_6_6_r;
wire signed [`CalcTempBus]          temp_m3_6_6_i;
wire signed [`CalcTempBus]          temp_m3_6_7_r;
wire signed [`CalcTempBus]          temp_m3_6_7_i;
wire signed [`CalcTempBus]          temp_m3_6_8_r;
wire signed [`CalcTempBus]          temp_m3_6_8_i;
wire signed [`CalcTempBus]          temp_m3_6_9_r;
wire signed [`CalcTempBus]          temp_m3_6_9_i;
wire signed [`CalcTempBus]          temp_m3_6_10_r;
wire signed [`CalcTempBus]          temp_m3_6_10_i;
wire signed [`CalcTempBus]          temp_m3_6_11_r;
wire signed [`CalcTempBus]          temp_m3_6_11_i;
wire signed [`CalcTempBus]          temp_m3_6_12_r;
wire signed [`CalcTempBus]          temp_m3_6_12_i;
wire signed [`CalcTempBus]          temp_m3_6_13_r;
wire signed [`CalcTempBus]          temp_m3_6_13_i;
wire signed [`CalcTempBus]          temp_m3_6_14_r;
wire signed [`CalcTempBus]          temp_m3_6_14_i;
wire signed [`CalcTempBus]          temp_m3_6_15_r;
wire signed [`CalcTempBus]          temp_m3_6_15_i;
wire signed [`CalcTempBus]          temp_m3_6_16_r;
wire signed [`CalcTempBus]          temp_m3_6_16_i;
wire signed [`CalcTempBus]          temp_m3_6_17_r;
wire signed [`CalcTempBus]          temp_m3_6_17_i;
wire signed [`CalcTempBus]          temp_m3_6_18_r;
wire signed [`CalcTempBus]          temp_m3_6_18_i;
wire signed [`CalcTempBus]          temp_m3_6_19_r;
wire signed [`CalcTempBus]          temp_m3_6_19_i;
wire signed [`CalcTempBus]          temp_m3_6_20_r;
wire signed [`CalcTempBus]          temp_m3_6_20_i;
wire signed [`CalcTempBus]          temp_m3_6_21_r;
wire signed [`CalcTempBus]          temp_m3_6_21_i;
wire signed [`CalcTempBus]          temp_m3_6_22_r;
wire signed [`CalcTempBus]          temp_m3_6_22_i;
wire signed [`CalcTempBus]          temp_m3_6_23_r;
wire signed [`CalcTempBus]          temp_m3_6_23_i;
wire signed [`CalcTempBus]          temp_m3_6_24_r;
wire signed [`CalcTempBus]          temp_m3_6_24_i;
wire signed [`CalcTempBus]          temp_m3_6_25_r;
wire signed [`CalcTempBus]          temp_m3_6_25_i;
wire signed [`CalcTempBus]          temp_m3_6_26_r;
wire signed [`CalcTempBus]          temp_m3_6_26_i;
wire signed [`CalcTempBus]          temp_m3_6_27_r;
wire signed [`CalcTempBus]          temp_m3_6_27_i;
wire signed [`CalcTempBus]          temp_m3_6_28_r;
wire signed [`CalcTempBus]          temp_m3_6_28_i;
wire signed [`CalcTempBus]          temp_m3_6_29_r;
wire signed [`CalcTempBus]          temp_m3_6_29_i;
wire signed [`CalcTempBus]          temp_m3_6_30_r;
wire signed [`CalcTempBus]          temp_m3_6_30_i;
wire signed [`CalcTempBus]          temp_m3_6_31_r;
wire signed [`CalcTempBus]          temp_m3_6_31_i;
wire signed [`CalcTempBus]          temp_m3_6_32_r;
wire signed [`CalcTempBus]          temp_m3_6_32_i;
wire signed [`CalcTempBus]          temp_m3_7_1_r;
wire signed [`CalcTempBus]          temp_m3_7_1_i;
wire signed [`CalcTempBus]          temp_m3_7_2_r;
wire signed [`CalcTempBus]          temp_m3_7_2_i;
wire signed [`CalcTempBus]          temp_m3_7_3_r;
wire signed [`CalcTempBus]          temp_m3_7_3_i;
wire signed [`CalcTempBus]          temp_m3_7_4_r;
wire signed [`CalcTempBus]          temp_m3_7_4_i;
wire signed [`CalcTempBus]          temp_m3_7_5_r;
wire signed [`CalcTempBus]          temp_m3_7_5_i;
wire signed [`CalcTempBus]          temp_m3_7_6_r;
wire signed [`CalcTempBus]          temp_m3_7_6_i;
wire signed [`CalcTempBus]          temp_m3_7_7_r;
wire signed [`CalcTempBus]          temp_m3_7_7_i;
wire signed [`CalcTempBus]          temp_m3_7_8_r;
wire signed [`CalcTempBus]          temp_m3_7_8_i;
wire signed [`CalcTempBus]          temp_m3_7_9_r;
wire signed [`CalcTempBus]          temp_m3_7_9_i;
wire signed [`CalcTempBus]          temp_m3_7_10_r;
wire signed [`CalcTempBus]          temp_m3_7_10_i;
wire signed [`CalcTempBus]          temp_m3_7_11_r;
wire signed [`CalcTempBus]          temp_m3_7_11_i;
wire signed [`CalcTempBus]          temp_m3_7_12_r;
wire signed [`CalcTempBus]          temp_m3_7_12_i;
wire signed [`CalcTempBus]          temp_m3_7_13_r;
wire signed [`CalcTempBus]          temp_m3_7_13_i;
wire signed [`CalcTempBus]          temp_m3_7_14_r;
wire signed [`CalcTempBus]          temp_m3_7_14_i;
wire signed [`CalcTempBus]          temp_m3_7_15_r;
wire signed [`CalcTempBus]          temp_m3_7_15_i;
wire signed [`CalcTempBus]          temp_m3_7_16_r;
wire signed [`CalcTempBus]          temp_m3_7_16_i;
wire signed [`CalcTempBus]          temp_m3_7_17_r;
wire signed [`CalcTempBus]          temp_m3_7_17_i;
wire signed [`CalcTempBus]          temp_m3_7_18_r;
wire signed [`CalcTempBus]          temp_m3_7_18_i;
wire signed [`CalcTempBus]          temp_m3_7_19_r;
wire signed [`CalcTempBus]          temp_m3_7_19_i;
wire signed [`CalcTempBus]          temp_m3_7_20_r;
wire signed [`CalcTempBus]          temp_m3_7_20_i;
wire signed [`CalcTempBus]          temp_m3_7_21_r;
wire signed [`CalcTempBus]          temp_m3_7_21_i;
wire signed [`CalcTempBus]          temp_m3_7_22_r;
wire signed [`CalcTempBus]          temp_m3_7_22_i;
wire signed [`CalcTempBus]          temp_m3_7_23_r;
wire signed [`CalcTempBus]          temp_m3_7_23_i;
wire signed [`CalcTempBus]          temp_m3_7_24_r;
wire signed [`CalcTempBus]          temp_m3_7_24_i;
wire signed [`CalcTempBus]          temp_m3_7_25_r;
wire signed [`CalcTempBus]          temp_m3_7_25_i;
wire signed [`CalcTempBus]          temp_m3_7_26_r;
wire signed [`CalcTempBus]          temp_m3_7_26_i;
wire signed [`CalcTempBus]          temp_m3_7_27_r;
wire signed [`CalcTempBus]          temp_m3_7_27_i;
wire signed [`CalcTempBus]          temp_m3_7_28_r;
wire signed [`CalcTempBus]          temp_m3_7_28_i;
wire signed [`CalcTempBus]          temp_m3_7_29_r;
wire signed [`CalcTempBus]          temp_m3_7_29_i;
wire signed [`CalcTempBus]          temp_m3_7_30_r;
wire signed [`CalcTempBus]          temp_m3_7_30_i;
wire signed [`CalcTempBus]          temp_m3_7_31_r;
wire signed [`CalcTempBus]          temp_m3_7_31_i;
wire signed [`CalcTempBus]          temp_m3_7_32_r;
wire signed [`CalcTempBus]          temp_m3_7_32_i;
wire signed [`CalcTempBus]          temp_m3_8_1_r;
wire signed [`CalcTempBus]          temp_m3_8_1_i;
wire signed [`CalcTempBus]          temp_m3_8_2_r;
wire signed [`CalcTempBus]          temp_m3_8_2_i;
wire signed [`CalcTempBus]          temp_m3_8_3_r;
wire signed [`CalcTempBus]          temp_m3_8_3_i;
wire signed [`CalcTempBus]          temp_m3_8_4_r;
wire signed [`CalcTempBus]          temp_m3_8_4_i;
wire signed [`CalcTempBus]          temp_m3_8_5_r;
wire signed [`CalcTempBus]          temp_m3_8_5_i;
wire signed [`CalcTempBus]          temp_m3_8_6_r;
wire signed [`CalcTempBus]          temp_m3_8_6_i;
wire signed [`CalcTempBus]          temp_m3_8_7_r;
wire signed [`CalcTempBus]          temp_m3_8_7_i;
wire signed [`CalcTempBus]          temp_m3_8_8_r;
wire signed [`CalcTempBus]          temp_m3_8_8_i;
wire signed [`CalcTempBus]          temp_m3_8_9_r;
wire signed [`CalcTempBus]          temp_m3_8_9_i;
wire signed [`CalcTempBus]          temp_m3_8_10_r;
wire signed [`CalcTempBus]          temp_m3_8_10_i;
wire signed [`CalcTempBus]          temp_m3_8_11_r;
wire signed [`CalcTempBus]          temp_m3_8_11_i;
wire signed [`CalcTempBus]          temp_m3_8_12_r;
wire signed [`CalcTempBus]          temp_m3_8_12_i;
wire signed [`CalcTempBus]          temp_m3_8_13_r;
wire signed [`CalcTempBus]          temp_m3_8_13_i;
wire signed [`CalcTempBus]          temp_m3_8_14_r;
wire signed [`CalcTempBus]          temp_m3_8_14_i;
wire signed [`CalcTempBus]          temp_m3_8_15_r;
wire signed [`CalcTempBus]          temp_m3_8_15_i;
wire signed [`CalcTempBus]          temp_m3_8_16_r;
wire signed [`CalcTempBus]          temp_m3_8_16_i;
wire signed [`CalcTempBus]          temp_m3_8_17_r;
wire signed [`CalcTempBus]          temp_m3_8_17_i;
wire signed [`CalcTempBus]          temp_m3_8_18_r;
wire signed [`CalcTempBus]          temp_m3_8_18_i;
wire signed [`CalcTempBus]          temp_m3_8_19_r;
wire signed [`CalcTempBus]          temp_m3_8_19_i;
wire signed [`CalcTempBus]          temp_m3_8_20_r;
wire signed [`CalcTempBus]          temp_m3_8_20_i;
wire signed [`CalcTempBus]          temp_m3_8_21_r;
wire signed [`CalcTempBus]          temp_m3_8_21_i;
wire signed [`CalcTempBus]          temp_m3_8_22_r;
wire signed [`CalcTempBus]          temp_m3_8_22_i;
wire signed [`CalcTempBus]          temp_m3_8_23_r;
wire signed [`CalcTempBus]          temp_m3_8_23_i;
wire signed [`CalcTempBus]          temp_m3_8_24_r;
wire signed [`CalcTempBus]          temp_m3_8_24_i;
wire signed [`CalcTempBus]          temp_m3_8_25_r;
wire signed [`CalcTempBus]          temp_m3_8_25_i;
wire signed [`CalcTempBus]          temp_m3_8_26_r;
wire signed [`CalcTempBus]          temp_m3_8_26_i;
wire signed [`CalcTempBus]          temp_m3_8_27_r;
wire signed [`CalcTempBus]          temp_m3_8_27_i;
wire signed [`CalcTempBus]          temp_m3_8_28_r;
wire signed [`CalcTempBus]          temp_m3_8_28_i;
wire signed [`CalcTempBus]          temp_m3_8_29_r;
wire signed [`CalcTempBus]          temp_m3_8_29_i;
wire signed [`CalcTempBus]          temp_m3_8_30_r;
wire signed [`CalcTempBus]          temp_m3_8_30_i;
wire signed [`CalcTempBus]          temp_m3_8_31_r;
wire signed [`CalcTempBus]          temp_m3_8_31_i;
wire signed [`CalcTempBus]          temp_m3_8_32_r;
wire signed [`CalcTempBus]          temp_m3_8_32_i;
wire signed [`CalcTempBus]          temp_m3_9_1_r;
wire signed [`CalcTempBus]          temp_m3_9_1_i;
wire signed [`CalcTempBus]          temp_m3_9_2_r;
wire signed [`CalcTempBus]          temp_m3_9_2_i;
wire signed [`CalcTempBus]          temp_m3_9_3_r;
wire signed [`CalcTempBus]          temp_m3_9_3_i;
wire signed [`CalcTempBus]          temp_m3_9_4_r;
wire signed [`CalcTempBus]          temp_m3_9_4_i;
wire signed [`CalcTempBus]          temp_m3_9_5_r;
wire signed [`CalcTempBus]          temp_m3_9_5_i;
wire signed [`CalcTempBus]          temp_m3_9_6_r;
wire signed [`CalcTempBus]          temp_m3_9_6_i;
wire signed [`CalcTempBus]          temp_m3_9_7_r;
wire signed [`CalcTempBus]          temp_m3_9_7_i;
wire signed [`CalcTempBus]          temp_m3_9_8_r;
wire signed [`CalcTempBus]          temp_m3_9_8_i;
wire signed [`CalcTempBus]          temp_m3_9_9_r;
wire signed [`CalcTempBus]          temp_m3_9_9_i;
wire signed [`CalcTempBus]          temp_m3_9_10_r;
wire signed [`CalcTempBus]          temp_m3_9_10_i;
wire signed [`CalcTempBus]          temp_m3_9_11_r;
wire signed [`CalcTempBus]          temp_m3_9_11_i;
wire signed [`CalcTempBus]          temp_m3_9_12_r;
wire signed [`CalcTempBus]          temp_m3_9_12_i;
wire signed [`CalcTempBus]          temp_m3_9_13_r;
wire signed [`CalcTempBus]          temp_m3_9_13_i;
wire signed [`CalcTempBus]          temp_m3_9_14_r;
wire signed [`CalcTempBus]          temp_m3_9_14_i;
wire signed [`CalcTempBus]          temp_m3_9_15_r;
wire signed [`CalcTempBus]          temp_m3_9_15_i;
wire signed [`CalcTempBus]          temp_m3_9_16_r;
wire signed [`CalcTempBus]          temp_m3_9_16_i;
wire signed [`CalcTempBus]          temp_m3_9_17_r;
wire signed [`CalcTempBus]          temp_m3_9_17_i;
wire signed [`CalcTempBus]          temp_m3_9_18_r;
wire signed [`CalcTempBus]          temp_m3_9_18_i;
wire signed [`CalcTempBus]          temp_m3_9_19_r;
wire signed [`CalcTempBus]          temp_m3_9_19_i;
wire signed [`CalcTempBus]          temp_m3_9_20_r;
wire signed [`CalcTempBus]          temp_m3_9_20_i;
wire signed [`CalcTempBus]          temp_m3_9_21_r;
wire signed [`CalcTempBus]          temp_m3_9_21_i;
wire signed [`CalcTempBus]          temp_m3_9_22_r;
wire signed [`CalcTempBus]          temp_m3_9_22_i;
wire signed [`CalcTempBus]          temp_m3_9_23_r;
wire signed [`CalcTempBus]          temp_m3_9_23_i;
wire signed [`CalcTempBus]          temp_m3_9_24_r;
wire signed [`CalcTempBus]          temp_m3_9_24_i;
wire signed [`CalcTempBus]          temp_m3_9_25_r;
wire signed [`CalcTempBus]          temp_m3_9_25_i;
wire signed [`CalcTempBus]          temp_m3_9_26_r;
wire signed [`CalcTempBus]          temp_m3_9_26_i;
wire signed [`CalcTempBus]          temp_m3_9_27_r;
wire signed [`CalcTempBus]          temp_m3_9_27_i;
wire signed [`CalcTempBus]          temp_m3_9_28_r;
wire signed [`CalcTempBus]          temp_m3_9_28_i;
wire signed [`CalcTempBus]          temp_m3_9_29_r;
wire signed [`CalcTempBus]          temp_m3_9_29_i;
wire signed [`CalcTempBus]          temp_m3_9_30_r;
wire signed [`CalcTempBus]          temp_m3_9_30_i;
wire signed [`CalcTempBus]          temp_m3_9_31_r;
wire signed [`CalcTempBus]          temp_m3_9_31_i;
wire signed [`CalcTempBus]          temp_m3_9_32_r;
wire signed [`CalcTempBus]          temp_m3_9_32_i;
wire signed [`CalcTempBus]          temp_m3_10_1_r;
wire signed [`CalcTempBus]          temp_m3_10_1_i;
wire signed [`CalcTempBus]          temp_m3_10_2_r;
wire signed [`CalcTempBus]          temp_m3_10_2_i;
wire signed [`CalcTempBus]          temp_m3_10_3_r;
wire signed [`CalcTempBus]          temp_m3_10_3_i;
wire signed [`CalcTempBus]          temp_m3_10_4_r;
wire signed [`CalcTempBus]          temp_m3_10_4_i;
wire signed [`CalcTempBus]          temp_m3_10_5_r;
wire signed [`CalcTempBus]          temp_m3_10_5_i;
wire signed [`CalcTempBus]          temp_m3_10_6_r;
wire signed [`CalcTempBus]          temp_m3_10_6_i;
wire signed [`CalcTempBus]          temp_m3_10_7_r;
wire signed [`CalcTempBus]          temp_m3_10_7_i;
wire signed [`CalcTempBus]          temp_m3_10_8_r;
wire signed [`CalcTempBus]          temp_m3_10_8_i;
wire signed [`CalcTempBus]          temp_m3_10_9_r;
wire signed [`CalcTempBus]          temp_m3_10_9_i;
wire signed [`CalcTempBus]          temp_m3_10_10_r;
wire signed [`CalcTempBus]          temp_m3_10_10_i;
wire signed [`CalcTempBus]          temp_m3_10_11_r;
wire signed [`CalcTempBus]          temp_m3_10_11_i;
wire signed [`CalcTempBus]          temp_m3_10_12_r;
wire signed [`CalcTempBus]          temp_m3_10_12_i;
wire signed [`CalcTempBus]          temp_m3_10_13_r;
wire signed [`CalcTempBus]          temp_m3_10_13_i;
wire signed [`CalcTempBus]          temp_m3_10_14_r;
wire signed [`CalcTempBus]          temp_m3_10_14_i;
wire signed [`CalcTempBus]          temp_m3_10_15_r;
wire signed [`CalcTempBus]          temp_m3_10_15_i;
wire signed [`CalcTempBus]          temp_m3_10_16_r;
wire signed [`CalcTempBus]          temp_m3_10_16_i;
wire signed [`CalcTempBus]          temp_m3_10_17_r;
wire signed [`CalcTempBus]          temp_m3_10_17_i;
wire signed [`CalcTempBus]          temp_m3_10_18_r;
wire signed [`CalcTempBus]          temp_m3_10_18_i;
wire signed [`CalcTempBus]          temp_m3_10_19_r;
wire signed [`CalcTempBus]          temp_m3_10_19_i;
wire signed [`CalcTempBus]          temp_m3_10_20_r;
wire signed [`CalcTempBus]          temp_m3_10_20_i;
wire signed [`CalcTempBus]          temp_m3_10_21_r;
wire signed [`CalcTempBus]          temp_m3_10_21_i;
wire signed [`CalcTempBus]          temp_m3_10_22_r;
wire signed [`CalcTempBus]          temp_m3_10_22_i;
wire signed [`CalcTempBus]          temp_m3_10_23_r;
wire signed [`CalcTempBus]          temp_m3_10_23_i;
wire signed [`CalcTempBus]          temp_m3_10_24_r;
wire signed [`CalcTempBus]          temp_m3_10_24_i;
wire signed [`CalcTempBus]          temp_m3_10_25_r;
wire signed [`CalcTempBus]          temp_m3_10_25_i;
wire signed [`CalcTempBus]          temp_m3_10_26_r;
wire signed [`CalcTempBus]          temp_m3_10_26_i;
wire signed [`CalcTempBus]          temp_m3_10_27_r;
wire signed [`CalcTempBus]          temp_m3_10_27_i;
wire signed [`CalcTempBus]          temp_m3_10_28_r;
wire signed [`CalcTempBus]          temp_m3_10_28_i;
wire signed [`CalcTempBus]          temp_m3_10_29_r;
wire signed [`CalcTempBus]          temp_m3_10_29_i;
wire signed [`CalcTempBus]          temp_m3_10_30_r;
wire signed [`CalcTempBus]          temp_m3_10_30_i;
wire signed [`CalcTempBus]          temp_m3_10_31_r;
wire signed [`CalcTempBus]          temp_m3_10_31_i;
wire signed [`CalcTempBus]          temp_m3_10_32_r;
wire signed [`CalcTempBus]          temp_m3_10_32_i;
wire signed [`CalcTempBus]          temp_m3_11_1_r;
wire signed [`CalcTempBus]          temp_m3_11_1_i;
wire signed [`CalcTempBus]          temp_m3_11_2_r;
wire signed [`CalcTempBus]          temp_m3_11_2_i;
wire signed [`CalcTempBus]          temp_m3_11_3_r;
wire signed [`CalcTempBus]          temp_m3_11_3_i;
wire signed [`CalcTempBus]          temp_m3_11_4_r;
wire signed [`CalcTempBus]          temp_m3_11_4_i;
wire signed [`CalcTempBus]          temp_m3_11_5_r;
wire signed [`CalcTempBus]          temp_m3_11_5_i;
wire signed [`CalcTempBus]          temp_m3_11_6_r;
wire signed [`CalcTempBus]          temp_m3_11_6_i;
wire signed [`CalcTempBus]          temp_m3_11_7_r;
wire signed [`CalcTempBus]          temp_m3_11_7_i;
wire signed [`CalcTempBus]          temp_m3_11_8_r;
wire signed [`CalcTempBus]          temp_m3_11_8_i;
wire signed [`CalcTempBus]          temp_m3_11_9_r;
wire signed [`CalcTempBus]          temp_m3_11_9_i;
wire signed [`CalcTempBus]          temp_m3_11_10_r;
wire signed [`CalcTempBus]          temp_m3_11_10_i;
wire signed [`CalcTempBus]          temp_m3_11_11_r;
wire signed [`CalcTempBus]          temp_m3_11_11_i;
wire signed [`CalcTempBus]          temp_m3_11_12_r;
wire signed [`CalcTempBus]          temp_m3_11_12_i;
wire signed [`CalcTempBus]          temp_m3_11_13_r;
wire signed [`CalcTempBus]          temp_m3_11_13_i;
wire signed [`CalcTempBus]          temp_m3_11_14_r;
wire signed [`CalcTempBus]          temp_m3_11_14_i;
wire signed [`CalcTempBus]          temp_m3_11_15_r;
wire signed [`CalcTempBus]          temp_m3_11_15_i;
wire signed [`CalcTempBus]          temp_m3_11_16_r;
wire signed [`CalcTempBus]          temp_m3_11_16_i;
wire signed [`CalcTempBus]          temp_m3_11_17_r;
wire signed [`CalcTempBus]          temp_m3_11_17_i;
wire signed [`CalcTempBus]          temp_m3_11_18_r;
wire signed [`CalcTempBus]          temp_m3_11_18_i;
wire signed [`CalcTempBus]          temp_m3_11_19_r;
wire signed [`CalcTempBus]          temp_m3_11_19_i;
wire signed [`CalcTempBus]          temp_m3_11_20_r;
wire signed [`CalcTempBus]          temp_m3_11_20_i;
wire signed [`CalcTempBus]          temp_m3_11_21_r;
wire signed [`CalcTempBus]          temp_m3_11_21_i;
wire signed [`CalcTempBus]          temp_m3_11_22_r;
wire signed [`CalcTempBus]          temp_m3_11_22_i;
wire signed [`CalcTempBus]          temp_m3_11_23_r;
wire signed [`CalcTempBus]          temp_m3_11_23_i;
wire signed [`CalcTempBus]          temp_m3_11_24_r;
wire signed [`CalcTempBus]          temp_m3_11_24_i;
wire signed [`CalcTempBus]          temp_m3_11_25_r;
wire signed [`CalcTempBus]          temp_m3_11_25_i;
wire signed [`CalcTempBus]          temp_m3_11_26_r;
wire signed [`CalcTempBus]          temp_m3_11_26_i;
wire signed [`CalcTempBus]          temp_m3_11_27_r;
wire signed [`CalcTempBus]          temp_m3_11_27_i;
wire signed [`CalcTempBus]          temp_m3_11_28_r;
wire signed [`CalcTempBus]          temp_m3_11_28_i;
wire signed [`CalcTempBus]          temp_m3_11_29_r;
wire signed [`CalcTempBus]          temp_m3_11_29_i;
wire signed [`CalcTempBus]          temp_m3_11_30_r;
wire signed [`CalcTempBus]          temp_m3_11_30_i;
wire signed [`CalcTempBus]          temp_m3_11_31_r;
wire signed [`CalcTempBus]          temp_m3_11_31_i;
wire signed [`CalcTempBus]          temp_m3_11_32_r;
wire signed [`CalcTempBus]          temp_m3_11_32_i;
wire signed [`CalcTempBus]          temp_m3_12_1_r;
wire signed [`CalcTempBus]          temp_m3_12_1_i;
wire signed [`CalcTempBus]          temp_m3_12_2_r;
wire signed [`CalcTempBus]          temp_m3_12_2_i;
wire signed [`CalcTempBus]          temp_m3_12_3_r;
wire signed [`CalcTempBus]          temp_m3_12_3_i;
wire signed [`CalcTempBus]          temp_m3_12_4_r;
wire signed [`CalcTempBus]          temp_m3_12_4_i;
wire signed [`CalcTempBus]          temp_m3_12_5_r;
wire signed [`CalcTempBus]          temp_m3_12_5_i;
wire signed [`CalcTempBus]          temp_m3_12_6_r;
wire signed [`CalcTempBus]          temp_m3_12_6_i;
wire signed [`CalcTempBus]          temp_m3_12_7_r;
wire signed [`CalcTempBus]          temp_m3_12_7_i;
wire signed [`CalcTempBus]          temp_m3_12_8_r;
wire signed [`CalcTempBus]          temp_m3_12_8_i;
wire signed [`CalcTempBus]          temp_m3_12_9_r;
wire signed [`CalcTempBus]          temp_m3_12_9_i;
wire signed [`CalcTempBus]          temp_m3_12_10_r;
wire signed [`CalcTempBus]          temp_m3_12_10_i;
wire signed [`CalcTempBus]          temp_m3_12_11_r;
wire signed [`CalcTempBus]          temp_m3_12_11_i;
wire signed [`CalcTempBus]          temp_m3_12_12_r;
wire signed [`CalcTempBus]          temp_m3_12_12_i;
wire signed [`CalcTempBus]          temp_m3_12_13_r;
wire signed [`CalcTempBus]          temp_m3_12_13_i;
wire signed [`CalcTempBus]          temp_m3_12_14_r;
wire signed [`CalcTempBus]          temp_m3_12_14_i;
wire signed [`CalcTempBus]          temp_m3_12_15_r;
wire signed [`CalcTempBus]          temp_m3_12_15_i;
wire signed [`CalcTempBus]          temp_m3_12_16_r;
wire signed [`CalcTempBus]          temp_m3_12_16_i;
wire signed [`CalcTempBus]          temp_m3_12_17_r;
wire signed [`CalcTempBus]          temp_m3_12_17_i;
wire signed [`CalcTempBus]          temp_m3_12_18_r;
wire signed [`CalcTempBus]          temp_m3_12_18_i;
wire signed [`CalcTempBus]          temp_m3_12_19_r;
wire signed [`CalcTempBus]          temp_m3_12_19_i;
wire signed [`CalcTempBus]          temp_m3_12_20_r;
wire signed [`CalcTempBus]          temp_m3_12_20_i;
wire signed [`CalcTempBus]          temp_m3_12_21_r;
wire signed [`CalcTempBus]          temp_m3_12_21_i;
wire signed [`CalcTempBus]          temp_m3_12_22_r;
wire signed [`CalcTempBus]          temp_m3_12_22_i;
wire signed [`CalcTempBus]          temp_m3_12_23_r;
wire signed [`CalcTempBus]          temp_m3_12_23_i;
wire signed [`CalcTempBus]          temp_m3_12_24_r;
wire signed [`CalcTempBus]          temp_m3_12_24_i;
wire signed [`CalcTempBus]          temp_m3_12_25_r;
wire signed [`CalcTempBus]          temp_m3_12_25_i;
wire signed [`CalcTempBus]          temp_m3_12_26_r;
wire signed [`CalcTempBus]          temp_m3_12_26_i;
wire signed [`CalcTempBus]          temp_m3_12_27_r;
wire signed [`CalcTempBus]          temp_m3_12_27_i;
wire signed [`CalcTempBus]          temp_m3_12_28_r;
wire signed [`CalcTempBus]          temp_m3_12_28_i;
wire signed [`CalcTempBus]          temp_m3_12_29_r;
wire signed [`CalcTempBus]          temp_m3_12_29_i;
wire signed [`CalcTempBus]          temp_m3_12_30_r;
wire signed [`CalcTempBus]          temp_m3_12_30_i;
wire signed [`CalcTempBus]          temp_m3_12_31_r;
wire signed [`CalcTempBus]          temp_m3_12_31_i;
wire signed [`CalcTempBus]          temp_m3_12_32_r;
wire signed [`CalcTempBus]          temp_m3_12_32_i;
wire signed [`CalcTempBus]          temp_m3_13_1_r;
wire signed [`CalcTempBus]          temp_m3_13_1_i;
wire signed [`CalcTempBus]          temp_m3_13_2_r;
wire signed [`CalcTempBus]          temp_m3_13_2_i;
wire signed [`CalcTempBus]          temp_m3_13_3_r;
wire signed [`CalcTempBus]          temp_m3_13_3_i;
wire signed [`CalcTempBus]          temp_m3_13_4_r;
wire signed [`CalcTempBus]          temp_m3_13_4_i;
wire signed [`CalcTempBus]          temp_m3_13_5_r;
wire signed [`CalcTempBus]          temp_m3_13_5_i;
wire signed [`CalcTempBus]          temp_m3_13_6_r;
wire signed [`CalcTempBus]          temp_m3_13_6_i;
wire signed [`CalcTempBus]          temp_m3_13_7_r;
wire signed [`CalcTempBus]          temp_m3_13_7_i;
wire signed [`CalcTempBus]          temp_m3_13_8_r;
wire signed [`CalcTempBus]          temp_m3_13_8_i;
wire signed [`CalcTempBus]          temp_m3_13_9_r;
wire signed [`CalcTempBus]          temp_m3_13_9_i;
wire signed [`CalcTempBus]          temp_m3_13_10_r;
wire signed [`CalcTempBus]          temp_m3_13_10_i;
wire signed [`CalcTempBus]          temp_m3_13_11_r;
wire signed [`CalcTempBus]          temp_m3_13_11_i;
wire signed [`CalcTempBus]          temp_m3_13_12_r;
wire signed [`CalcTempBus]          temp_m3_13_12_i;
wire signed [`CalcTempBus]          temp_m3_13_13_r;
wire signed [`CalcTempBus]          temp_m3_13_13_i;
wire signed [`CalcTempBus]          temp_m3_13_14_r;
wire signed [`CalcTempBus]          temp_m3_13_14_i;
wire signed [`CalcTempBus]          temp_m3_13_15_r;
wire signed [`CalcTempBus]          temp_m3_13_15_i;
wire signed [`CalcTempBus]          temp_m3_13_16_r;
wire signed [`CalcTempBus]          temp_m3_13_16_i;
wire signed [`CalcTempBus]          temp_m3_13_17_r;
wire signed [`CalcTempBus]          temp_m3_13_17_i;
wire signed [`CalcTempBus]          temp_m3_13_18_r;
wire signed [`CalcTempBus]          temp_m3_13_18_i;
wire signed [`CalcTempBus]          temp_m3_13_19_r;
wire signed [`CalcTempBus]          temp_m3_13_19_i;
wire signed [`CalcTempBus]          temp_m3_13_20_r;
wire signed [`CalcTempBus]          temp_m3_13_20_i;
wire signed [`CalcTempBus]          temp_m3_13_21_r;
wire signed [`CalcTempBus]          temp_m3_13_21_i;
wire signed [`CalcTempBus]          temp_m3_13_22_r;
wire signed [`CalcTempBus]          temp_m3_13_22_i;
wire signed [`CalcTempBus]          temp_m3_13_23_r;
wire signed [`CalcTempBus]          temp_m3_13_23_i;
wire signed [`CalcTempBus]          temp_m3_13_24_r;
wire signed [`CalcTempBus]          temp_m3_13_24_i;
wire signed [`CalcTempBus]          temp_m3_13_25_r;
wire signed [`CalcTempBus]          temp_m3_13_25_i;
wire signed [`CalcTempBus]          temp_m3_13_26_r;
wire signed [`CalcTempBus]          temp_m3_13_26_i;
wire signed [`CalcTempBus]          temp_m3_13_27_r;
wire signed [`CalcTempBus]          temp_m3_13_27_i;
wire signed [`CalcTempBus]          temp_m3_13_28_r;
wire signed [`CalcTempBus]          temp_m3_13_28_i;
wire signed [`CalcTempBus]          temp_m3_13_29_r;
wire signed [`CalcTempBus]          temp_m3_13_29_i;
wire signed [`CalcTempBus]          temp_m3_13_30_r;
wire signed [`CalcTempBus]          temp_m3_13_30_i;
wire signed [`CalcTempBus]          temp_m3_13_31_r;
wire signed [`CalcTempBus]          temp_m3_13_31_i;
wire signed [`CalcTempBus]          temp_m3_13_32_r;
wire signed [`CalcTempBus]          temp_m3_13_32_i;
wire signed [`CalcTempBus]          temp_m3_14_1_r;
wire signed [`CalcTempBus]          temp_m3_14_1_i;
wire signed [`CalcTempBus]          temp_m3_14_2_r;
wire signed [`CalcTempBus]          temp_m3_14_2_i;
wire signed [`CalcTempBus]          temp_m3_14_3_r;
wire signed [`CalcTempBus]          temp_m3_14_3_i;
wire signed [`CalcTempBus]          temp_m3_14_4_r;
wire signed [`CalcTempBus]          temp_m3_14_4_i;
wire signed [`CalcTempBus]          temp_m3_14_5_r;
wire signed [`CalcTempBus]          temp_m3_14_5_i;
wire signed [`CalcTempBus]          temp_m3_14_6_r;
wire signed [`CalcTempBus]          temp_m3_14_6_i;
wire signed [`CalcTempBus]          temp_m3_14_7_r;
wire signed [`CalcTempBus]          temp_m3_14_7_i;
wire signed [`CalcTempBus]          temp_m3_14_8_r;
wire signed [`CalcTempBus]          temp_m3_14_8_i;
wire signed [`CalcTempBus]          temp_m3_14_9_r;
wire signed [`CalcTempBus]          temp_m3_14_9_i;
wire signed [`CalcTempBus]          temp_m3_14_10_r;
wire signed [`CalcTempBus]          temp_m3_14_10_i;
wire signed [`CalcTempBus]          temp_m3_14_11_r;
wire signed [`CalcTempBus]          temp_m3_14_11_i;
wire signed [`CalcTempBus]          temp_m3_14_12_r;
wire signed [`CalcTempBus]          temp_m3_14_12_i;
wire signed [`CalcTempBus]          temp_m3_14_13_r;
wire signed [`CalcTempBus]          temp_m3_14_13_i;
wire signed [`CalcTempBus]          temp_m3_14_14_r;
wire signed [`CalcTempBus]          temp_m3_14_14_i;
wire signed [`CalcTempBus]          temp_m3_14_15_r;
wire signed [`CalcTempBus]          temp_m3_14_15_i;
wire signed [`CalcTempBus]          temp_m3_14_16_r;
wire signed [`CalcTempBus]          temp_m3_14_16_i;
wire signed [`CalcTempBus]          temp_m3_14_17_r;
wire signed [`CalcTempBus]          temp_m3_14_17_i;
wire signed [`CalcTempBus]          temp_m3_14_18_r;
wire signed [`CalcTempBus]          temp_m3_14_18_i;
wire signed [`CalcTempBus]          temp_m3_14_19_r;
wire signed [`CalcTempBus]          temp_m3_14_19_i;
wire signed [`CalcTempBus]          temp_m3_14_20_r;
wire signed [`CalcTempBus]          temp_m3_14_20_i;
wire signed [`CalcTempBus]          temp_m3_14_21_r;
wire signed [`CalcTempBus]          temp_m3_14_21_i;
wire signed [`CalcTempBus]          temp_m3_14_22_r;
wire signed [`CalcTempBus]          temp_m3_14_22_i;
wire signed [`CalcTempBus]          temp_m3_14_23_r;
wire signed [`CalcTempBus]          temp_m3_14_23_i;
wire signed [`CalcTempBus]          temp_m3_14_24_r;
wire signed [`CalcTempBus]          temp_m3_14_24_i;
wire signed [`CalcTempBus]          temp_m3_14_25_r;
wire signed [`CalcTempBus]          temp_m3_14_25_i;
wire signed [`CalcTempBus]          temp_m3_14_26_r;
wire signed [`CalcTempBus]          temp_m3_14_26_i;
wire signed [`CalcTempBus]          temp_m3_14_27_r;
wire signed [`CalcTempBus]          temp_m3_14_27_i;
wire signed [`CalcTempBus]          temp_m3_14_28_r;
wire signed [`CalcTempBus]          temp_m3_14_28_i;
wire signed [`CalcTempBus]          temp_m3_14_29_r;
wire signed [`CalcTempBus]          temp_m3_14_29_i;
wire signed [`CalcTempBus]          temp_m3_14_30_r;
wire signed [`CalcTempBus]          temp_m3_14_30_i;
wire signed [`CalcTempBus]          temp_m3_14_31_r;
wire signed [`CalcTempBus]          temp_m3_14_31_i;
wire signed [`CalcTempBus]          temp_m3_14_32_r;
wire signed [`CalcTempBus]          temp_m3_14_32_i;
wire signed [`CalcTempBus]          temp_m3_15_1_r;
wire signed [`CalcTempBus]          temp_m3_15_1_i;
wire signed [`CalcTempBus]          temp_m3_15_2_r;
wire signed [`CalcTempBus]          temp_m3_15_2_i;
wire signed [`CalcTempBus]          temp_m3_15_3_r;
wire signed [`CalcTempBus]          temp_m3_15_3_i;
wire signed [`CalcTempBus]          temp_m3_15_4_r;
wire signed [`CalcTempBus]          temp_m3_15_4_i;
wire signed [`CalcTempBus]          temp_m3_15_5_r;
wire signed [`CalcTempBus]          temp_m3_15_5_i;
wire signed [`CalcTempBus]          temp_m3_15_6_r;
wire signed [`CalcTempBus]          temp_m3_15_6_i;
wire signed [`CalcTempBus]          temp_m3_15_7_r;
wire signed [`CalcTempBus]          temp_m3_15_7_i;
wire signed [`CalcTempBus]          temp_m3_15_8_r;
wire signed [`CalcTempBus]          temp_m3_15_8_i;
wire signed [`CalcTempBus]          temp_m3_15_9_r;
wire signed [`CalcTempBus]          temp_m3_15_9_i;
wire signed [`CalcTempBus]          temp_m3_15_10_r;
wire signed [`CalcTempBus]          temp_m3_15_10_i;
wire signed [`CalcTempBus]          temp_m3_15_11_r;
wire signed [`CalcTempBus]          temp_m3_15_11_i;
wire signed [`CalcTempBus]          temp_m3_15_12_r;
wire signed [`CalcTempBus]          temp_m3_15_12_i;
wire signed [`CalcTempBus]          temp_m3_15_13_r;
wire signed [`CalcTempBus]          temp_m3_15_13_i;
wire signed [`CalcTempBus]          temp_m3_15_14_r;
wire signed [`CalcTempBus]          temp_m3_15_14_i;
wire signed [`CalcTempBus]          temp_m3_15_15_r;
wire signed [`CalcTempBus]          temp_m3_15_15_i;
wire signed [`CalcTempBus]          temp_m3_15_16_r;
wire signed [`CalcTempBus]          temp_m3_15_16_i;
wire signed [`CalcTempBus]          temp_m3_15_17_r;
wire signed [`CalcTempBus]          temp_m3_15_17_i;
wire signed [`CalcTempBus]          temp_m3_15_18_r;
wire signed [`CalcTempBus]          temp_m3_15_18_i;
wire signed [`CalcTempBus]          temp_m3_15_19_r;
wire signed [`CalcTempBus]          temp_m3_15_19_i;
wire signed [`CalcTempBus]          temp_m3_15_20_r;
wire signed [`CalcTempBus]          temp_m3_15_20_i;
wire signed [`CalcTempBus]          temp_m3_15_21_r;
wire signed [`CalcTempBus]          temp_m3_15_21_i;
wire signed [`CalcTempBus]          temp_m3_15_22_r;
wire signed [`CalcTempBus]          temp_m3_15_22_i;
wire signed [`CalcTempBus]          temp_m3_15_23_r;
wire signed [`CalcTempBus]          temp_m3_15_23_i;
wire signed [`CalcTempBus]          temp_m3_15_24_r;
wire signed [`CalcTempBus]          temp_m3_15_24_i;
wire signed [`CalcTempBus]          temp_m3_15_25_r;
wire signed [`CalcTempBus]          temp_m3_15_25_i;
wire signed [`CalcTempBus]          temp_m3_15_26_r;
wire signed [`CalcTempBus]          temp_m3_15_26_i;
wire signed [`CalcTempBus]          temp_m3_15_27_r;
wire signed [`CalcTempBus]          temp_m3_15_27_i;
wire signed [`CalcTempBus]          temp_m3_15_28_r;
wire signed [`CalcTempBus]          temp_m3_15_28_i;
wire signed [`CalcTempBus]          temp_m3_15_29_r;
wire signed [`CalcTempBus]          temp_m3_15_29_i;
wire signed [`CalcTempBus]          temp_m3_15_30_r;
wire signed [`CalcTempBus]          temp_m3_15_30_i;
wire signed [`CalcTempBus]          temp_m3_15_31_r;
wire signed [`CalcTempBus]          temp_m3_15_31_i;
wire signed [`CalcTempBus]          temp_m3_15_32_r;
wire signed [`CalcTempBus]          temp_m3_15_32_i;
wire signed [`CalcTempBus]          temp_m3_16_1_r;
wire signed [`CalcTempBus]          temp_m3_16_1_i;
wire signed [`CalcTempBus]          temp_m3_16_2_r;
wire signed [`CalcTempBus]          temp_m3_16_2_i;
wire signed [`CalcTempBus]          temp_m3_16_3_r;
wire signed [`CalcTempBus]          temp_m3_16_3_i;
wire signed [`CalcTempBus]          temp_m3_16_4_r;
wire signed [`CalcTempBus]          temp_m3_16_4_i;
wire signed [`CalcTempBus]          temp_m3_16_5_r;
wire signed [`CalcTempBus]          temp_m3_16_5_i;
wire signed [`CalcTempBus]          temp_m3_16_6_r;
wire signed [`CalcTempBus]          temp_m3_16_6_i;
wire signed [`CalcTempBus]          temp_m3_16_7_r;
wire signed [`CalcTempBus]          temp_m3_16_7_i;
wire signed [`CalcTempBus]          temp_m3_16_8_r;
wire signed [`CalcTempBus]          temp_m3_16_8_i;
wire signed [`CalcTempBus]          temp_m3_16_9_r;
wire signed [`CalcTempBus]          temp_m3_16_9_i;
wire signed [`CalcTempBus]          temp_m3_16_10_r;
wire signed [`CalcTempBus]          temp_m3_16_10_i;
wire signed [`CalcTempBus]          temp_m3_16_11_r;
wire signed [`CalcTempBus]          temp_m3_16_11_i;
wire signed [`CalcTempBus]          temp_m3_16_12_r;
wire signed [`CalcTempBus]          temp_m3_16_12_i;
wire signed [`CalcTempBus]          temp_m3_16_13_r;
wire signed [`CalcTempBus]          temp_m3_16_13_i;
wire signed [`CalcTempBus]          temp_m3_16_14_r;
wire signed [`CalcTempBus]          temp_m3_16_14_i;
wire signed [`CalcTempBus]          temp_m3_16_15_r;
wire signed [`CalcTempBus]          temp_m3_16_15_i;
wire signed [`CalcTempBus]          temp_m3_16_16_r;
wire signed [`CalcTempBus]          temp_m3_16_16_i;
wire signed [`CalcTempBus]          temp_m3_16_17_r;
wire signed [`CalcTempBus]          temp_m3_16_17_i;
wire signed [`CalcTempBus]          temp_m3_16_18_r;
wire signed [`CalcTempBus]          temp_m3_16_18_i;
wire signed [`CalcTempBus]          temp_m3_16_19_r;
wire signed [`CalcTempBus]          temp_m3_16_19_i;
wire signed [`CalcTempBus]          temp_m3_16_20_r;
wire signed [`CalcTempBus]          temp_m3_16_20_i;
wire signed [`CalcTempBus]          temp_m3_16_21_r;
wire signed [`CalcTempBus]          temp_m3_16_21_i;
wire signed [`CalcTempBus]          temp_m3_16_22_r;
wire signed [`CalcTempBus]          temp_m3_16_22_i;
wire signed [`CalcTempBus]          temp_m3_16_23_r;
wire signed [`CalcTempBus]          temp_m3_16_23_i;
wire signed [`CalcTempBus]          temp_m3_16_24_r;
wire signed [`CalcTempBus]          temp_m3_16_24_i;
wire signed [`CalcTempBus]          temp_m3_16_25_r;
wire signed [`CalcTempBus]          temp_m3_16_25_i;
wire signed [`CalcTempBus]          temp_m3_16_26_r;
wire signed [`CalcTempBus]          temp_m3_16_26_i;
wire signed [`CalcTempBus]          temp_m3_16_27_r;
wire signed [`CalcTempBus]          temp_m3_16_27_i;
wire signed [`CalcTempBus]          temp_m3_16_28_r;
wire signed [`CalcTempBus]          temp_m3_16_28_i;
wire signed [`CalcTempBus]          temp_m3_16_29_r;
wire signed [`CalcTempBus]          temp_m3_16_29_i;
wire signed [`CalcTempBus]          temp_m3_16_30_r;
wire signed [`CalcTempBus]          temp_m3_16_30_i;
wire signed [`CalcTempBus]          temp_m3_16_31_r;
wire signed [`CalcTempBus]          temp_m3_16_31_i;
wire signed [`CalcTempBus]          temp_m3_16_32_r;
wire signed [`CalcTempBus]          temp_m3_16_32_i;
wire signed [`CalcTempBus]          temp_m3_17_1_r;
wire signed [`CalcTempBus]          temp_m3_17_1_i;
wire signed [`CalcTempBus]          temp_m3_17_2_r;
wire signed [`CalcTempBus]          temp_m3_17_2_i;
wire signed [`CalcTempBus]          temp_m3_17_3_r;
wire signed [`CalcTempBus]          temp_m3_17_3_i;
wire signed [`CalcTempBus]          temp_m3_17_4_r;
wire signed [`CalcTempBus]          temp_m3_17_4_i;
wire signed [`CalcTempBus]          temp_m3_17_5_r;
wire signed [`CalcTempBus]          temp_m3_17_5_i;
wire signed [`CalcTempBus]          temp_m3_17_6_r;
wire signed [`CalcTempBus]          temp_m3_17_6_i;
wire signed [`CalcTempBus]          temp_m3_17_7_r;
wire signed [`CalcTempBus]          temp_m3_17_7_i;
wire signed [`CalcTempBus]          temp_m3_17_8_r;
wire signed [`CalcTempBus]          temp_m3_17_8_i;
wire signed [`CalcTempBus]          temp_m3_17_9_r;
wire signed [`CalcTempBus]          temp_m3_17_9_i;
wire signed [`CalcTempBus]          temp_m3_17_10_r;
wire signed [`CalcTempBus]          temp_m3_17_10_i;
wire signed [`CalcTempBus]          temp_m3_17_11_r;
wire signed [`CalcTempBus]          temp_m3_17_11_i;
wire signed [`CalcTempBus]          temp_m3_17_12_r;
wire signed [`CalcTempBus]          temp_m3_17_12_i;
wire signed [`CalcTempBus]          temp_m3_17_13_r;
wire signed [`CalcTempBus]          temp_m3_17_13_i;
wire signed [`CalcTempBus]          temp_m3_17_14_r;
wire signed [`CalcTempBus]          temp_m3_17_14_i;
wire signed [`CalcTempBus]          temp_m3_17_15_r;
wire signed [`CalcTempBus]          temp_m3_17_15_i;
wire signed [`CalcTempBus]          temp_m3_17_16_r;
wire signed [`CalcTempBus]          temp_m3_17_16_i;
wire signed [`CalcTempBus]          temp_m3_17_17_r;
wire signed [`CalcTempBus]          temp_m3_17_17_i;
wire signed [`CalcTempBus]          temp_m3_17_18_r;
wire signed [`CalcTempBus]          temp_m3_17_18_i;
wire signed [`CalcTempBus]          temp_m3_17_19_r;
wire signed [`CalcTempBus]          temp_m3_17_19_i;
wire signed [`CalcTempBus]          temp_m3_17_20_r;
wire signed [`CalcTempBus]          temp_m3_17_20_i;
wire signed [`CalcTempBus]          temp_m3_17_21_r;
wire signed [`CalcTempBus]          temp_m3_17_21_i;
wire signed [`CalcTempBus]          temp_m3_17_22_r;
wire signed [`CalcTempBus]          temp_m3_17_22_i;
wire signed [`CalcTempBus]          temp_m3_17_23_r;
wire signed [`CalcTempBus]          temp_m3_17_23_i;
wire signed [`CalcTempBus]          temp_m3_17_24_r;
wire signed [`CalcTempBus]          temp_m3_17_24_i;
wire signed [`CalcTempBus]          temp_m3_17_25_r;
wire signed [`CalcTempBus]          temp_m3_17_25_i;
wire signed [`CalcTempBus]          temp_m3_17_26_r;
wire signed [`CalcTempBus]          temp_m3_17_26_i;
wire signed [`CalcTempBus]          temp_m3_17_27_r;
wire signed [`CalcTempBus]          temp_m3_17_27_i;
wire signed [`CalcTempBus]          temp_m3_17_28_r;
wire signed [`CalcTempBus]          temp_m3_17_28_i;
wire signed [`CalcTempBus]          temp_m3_17_29_r;
wire signed [`CalcTempBus]          temp_m3_17_29_i;
wire signed [`CalcTempBus]          temp_m3_17_30_r;
wire signed [`CalcTempBus]          temp_m3_17_30_i;
wire signed [`CalcTempBus]          temp_m3_17_31_r;
wire signed [`CalcTempBus]          temp_m3_17_31_i;
wire signed [`CalcTempBus]          temp_m3_17_32_r;
wire signed [`CalcTempBus]          temp_m3_17_32_i;
wire signed [`CalcTempBus]          temp_m3_18_1_r;
wire signed [`CalcTempBus]          temp_m3_18_1_i;
wire signed [`CalcTempBus]          temp_m3_18_2_r;
wire signed [`CalcTempBus]          temp_m3_18_2_i;
wire signed [`CalcTempBus]          temp_m3_18_3_r;
wire signed [`CalcTempBus]          temp_m3_18_3_i;
wire signed [`CalcTempBus]          temp_m3_18_4_r;
wire signed [`CalcTempBus]          temp_m3_18_4_i;
wire signed [`CalcTempBus]          temp_m3_18_5_r;
wire signed [`CalcTempBus]          temp_m3_18_5_i;
wire signed [`CalcTempBus]          temp_m3_18_6_r;
wire signed [`CalcTempBus]          temp_m3_18_6_i;
wire signed [`CalcTempBus]          temp_m3_18_7_r;
wire signed [`CalcTempBus]          temp_m3_18_7_i;
wire signed [`CalcTempBus]          temp_m3_18_8_r;
wire signed [`CalcTempBus]          temp_m3_18_8_i;
wire signed [`CalcTempBus]          temp_m3_18_9_r;
wire signed [`CalcTempBus]          temp_m3_18_9_i;
wire signed [`CalcTempBus]          temp_m3_18_10_r;
wire signed [`CalcTempBus]          temp_m3_18_10_i;
wire signed [`CalcTempBus]          temp_m3_18_11_r;
wire signed [`CalcTempBus]          temp_m3_18_11_i;
wire signed [`CalcTempBus]          temp_m3_18_12_r;
wire signed [`CalcTempBus]          temp_m3_18_12_i;
wire signed [`CalcTempBus]          temp_m3_18_13_r;
wire signed [`CalcTempBus]          temp_m3_18_13_i;
wire signed [`CalcTempBus]          temp_m3_18_14_r;
wire signed [`CalcTempBus]          temp_m3_18_14_i;
wire signed [`CalcTempBus]          temp_m3_18_15_r;
wire signed [`CalcTempBus]          temp_m3_18_15_i;
wire signed [`CalcTempBus]          temp_m3_18_16_r;
wire signed [`CalcTempBus]          temp_m3_18_16_i;
wire signed [`CalcTempBus]          temp_m3_18_17_r;
wire signed [`CalcTempBus]          temp_m3_18_17_i;
wire signed [`CalcTempBus]          temp_m3_18_18_r;
wire signed [`CalcTempBus]          temp_m3_18_18_i;
wire signed [`CalcTempBus]          temp_m3_18_19_r;
wire signed [`CalcTempBus]          temp_m3_18_19_i;
wire signed [`CalcTempBus]          temp_m3_18_20_r;
wire signed [`CalcTempBus]          temp_m3_18_20_i;
wire signed [`CalcTempBus]          temp_m3_18_21_r;
wire signed [`CalcTempBus]          temp_m3_18_21_i;
wire signed [`CalcTempBus]          temp_m3_18_22_r;
wire signed [`CalcTempBus]          temp_m3_18_22_i;
wire signed [`CalcTempBus]          temp_m3_18_23_r;
wire signed [`CalcTempBus]          temp_m3_18_23_i;
wire signed [`CalcTempBus]          temp_m3_18_24_r;
wire signed [`CalcTempBus]          temp_m3_18_24_i;
wire signed [`CalcTempBus]          temp_m3_18_25_r;
wire signed [`CalcTempBus]          temp_m3_18_25_i;
wire signed [`CalcTempBus]          temp_m3_18_26_r;
wire signed [`CalcTempBus]          temp_m3_18_26_i;
wire signed [`CalcTempBus]          temp_m3_18_27_r;
wire signed [`CalcTempBus]          temp_m3_18_27_i;
wire signed [`CalcTempBus]          temp_m3_18_28_r;
wire signed [`CalcTempBus]          temp_m3_18_28_i;
wire signed [`CalcTempBus]          temp_m3_18_29_r;
wire signed [`CalcTempBus]          temp_m3_18_29_i;
wire signed [`CalcTempBus]          temp_m3_18_30_r;
wire signed [`CalcTempBus]          temp_m3_18_30_i;
wire signed [`CalcTempBus]          temp_m3_18_31_r;
wire signed [`CalcTempBus]          temp_m3_18_31_i;
wire signed [`CalcTempBus]          temp_m3_18_32_r;
wire signed [`CalcTempBus]          temp_m3_18_32_i;
wire signed [`CalcTempBus]          temp_m3_19_1_r;
wire signed [`CalcTempBus]          temp_m3_19_1_i;
wire signed [`CalcTempBus]          temp_m3_19_2_r;
wire signed [`CalcTempBus]          temp_m3_19_2_i;
wire signed [`CalcTempBus]          temp_m3_19_3_r;
wire signed [`CalcTempBus]          temp_m3_19_3_i;
wire signed [`CalcTempBus]          temp_m3_19_4_r;
wire signed [`CalcTempBus]          temp_m3_19_4_i;
wire signed [`CalcTempBus]          temp_m3_19_5_r;
wire signed [`CalcTempBus]          temp_m3_19_5_i;
wire signed [`CalcTempBus]          temp_m3_19_6_r;
wire signed [`CalcTempBus]          temp_m3_19_6_i;
wire signed [`CalcTempBus]          temp_m3_19_7_r;
wire signed [`CalcTempBus]          temp_m3_19_7_i;
wire signed [`CalcTempBus]          temp_m3_19_8_r;
wire signed [`CalcTempBus]          temp_m3_19_8_i;
wire signed [`CalcTempBus]          temp_m3_19_9_r;
wire signed [`CalcTempBus]          temp_m3_19_9_i;
wire signed [`CalcTempBus]          temp_m3_19_10_r;
wire signed [`CalcTempBus]          temp_m3_19_10_i;
wire signed [`CalcTempBus]          temp_m3_19_11_r;
wire signed [`CalcTempBus]          temp_m3_19_11_i;
wire signed [`CalcTempBus]          temp_m3_19_12_r;
wire signed [`CalcTempBus]          temp_m3_19_12_i;
wire signed [`CalcTempBus]          temp_m3_19_13_r;
wire signed [`CalcTempBus]          temp_m3_19_13_i;
wire signed [`CalcTempBus]          temp_m3_19_14_r;
wire signed [`CalcTempBus]          temp_m3_19_14_i;
wire signed [`CalcTempBus]          temp_m3_19_15_r;
wire signed [`CalcTempBus]          temp_m3_19_15_i;
wire signed [`CalcTempBus]          temp_m3_19_16_r;
wire signed [`CalcTempBus]          temp_m3_19_16_i;
wire signed [`CalcTempBus]          temp_m3_19_17_r;
wire signed [`CalcTempBus]          temp_m3_19_17_i;
wire signed [`CalcTempBus]          temp_m3_19_18_r;
wire signed [`CalcTempBus]          temp_m3_19_18_i;
wire signed [`CalcTempBus]          temp_m3_19_19_r;
wire signed [`CalcTempBus]          temp_m3_19_19_i;
wire signed [`CalcTempBus]          temp_m3_19_20_r;
wire signed [`CalcTempBus]          temp_m3_19_20_i;
wire signed [`CalcTempBus]          temp_m3_19_21_r;
wire signed [`CalcTempBus]          temp_m3_19_21_i;
wire signed [`CalcTempBus]          temp_m3_19_22_r;
wire signed [`CalcTempBus]          temp_m3_19_22_i;
wire signed [`CalcTempBus]          temp_m3_19_23_r;
wire signed [`CalcTempBus]          temp_m3_19_23_i;
wire signed [`CalcTempBus]          temp_m3_19_24_r;
wire signed [`CalcTempBus]          temp_m3_19_24_i;
wire signed [`CalcTempBus]          temp_m3_19_25_r;
wire signed [`CalcTempBus]          temp_m3_19_25_i;
wire signed [`CalcTempBus]          temp_m3_19_26_r;
wire signed [`CalcTempBus]          temp_m3_19_26_i;
wire signed [`CalcTempBus]          temp_m3_19_27_r;
wire signed [`CalcTempBus]          temp_m3_19_27_i;
wire signed [`CalcTempBus]          temp_m3_19_28_r;
wire signed [`CalcTempBus]          temp_m3_19_28_i;
wire signed [`CalcTempBus]          temp_m3_19_29_r;
wire signed [`CalcTempBus]          temp_m3_19_29_i;
wire signed [`CalcTempBus]          temp_m3_19_30_r;
wire signed [`CalcTempBus]          temp_m3_19_30_i;
wire signed [`CalcTempBus]          temp_m3_19_31_r;
wire signed [`CalcTempBus]          temp_m3_19_31_i;
wire signed [`CalcTempBus]          temp_m3_19_32_r;
wire signed [`CalcTempBus]          temp_m3_19_32_i;
wire signed [`CalcTempBus]          temp_m3_20_1_r;
wire signed [`CalcTempBus]          temp_m3_20_1_i;
wire signed [`CalcTempBus]          temp_m3_20_2_r;
wire signed [`CalcTempBus]          temp_m3_20_2_i;
wire signed [`CalcTempBus]          temp_m3_20_3_r;
wire signed [`CalcTempBus]          temp_m3_20_3_i;
wire signed [`CalcTempBus]          temp_m3_20_4_r;
wire signed [`CalcTempBus]          temp_m3_20_4_i;
wire signed [`CalcTempBus]          temp_m3_20_5_r;
wire signed [`CalcTempBus]          temp_m3_20_5_i;
wire signed [`CalcTempBus]          temp_m3_20_6_r;
wire signed [`CalcTempBus]          temp_m3_20_6_i;
wire signed [`CalcTempBus]          temp_m3_20_7_r;
wire signed [`CalcTempBus]          temp_m3_20_7_i;
wire signed [`CalcTempBus]          temp_m3_20_8_r;
wire signed [`CalcTempBus]          temp_m3_20_8_i;
wire signed [`CalcTempBus]          temp_m3_20_9_r;
wire signed [`CalcTempBus]          temp_m3_20_9_i;
wire signed [`CalcTempBus]          temp_m3_20_10_r;
wire signed [`CalcTempBus]          temp_m3_20_10_i;
wire signed [`CalcTempBus]          temp_m3_20_11_r;
wire signed [`CalcTempBus]          temp_m3_20_11_i;
wire signed [`CalcTempBus]          temp_m3_20_12_r;
wire signed [`CalcTempBus]          temp_m3_20_12_i;
wire signed [`CalcTempBus]          temp_m3_20_13_r;
wire signed [`CalcTempBus]          temp_m3_20_13_i;
wire signed [`CalcTempBus]          temp_m3_20_14_r;
wire signed [`CalcTempBus]          temp_m3_20_14_i;
wire signed [`CalcTempBus]          temp_m3_20_15_r;
wire signed [`CalcTempBus]          temp_m3_20_15_i;
wire signed [`CalcTempBus]          temp_m3_20_16_r;
wire signed [`CalcTempBus]          temp_m3_20_16_i;
wire signed [`CalcTempBus]          temp_m3_20_17_r;
wire signed [`CalcTempBus]          temp_m3_20_17_i;
wire signed [`CalcTempBus]          temp_m3_20_18_r;
wire signed [`CalcTempBus]          temp_m3_20_18_i;
wire signed [`CalcTempBus]          temp_m3_20_19_r;
wire signed [`CalcTempBus]          temp_m3_20_19_i;
wire signed [`CalcTempBus]          temp_m3_20_20_r;
wire signed [`CalcTempBus]          temp_m3_20_20_i;
wire signed [`CalcTempBus]          temp_m3_20_21_r;
wire signed [`CalcTempBus]          temp_m3_20_21_i;
wire signed [`CalcTempBus]          temp_m3_20_22_r;
wire signed [`CalcTempBus]          temp_m3_20_22_i;
wire signed [`CalcTempBus]          temp_m3_20_23_r;
wire signed [`CalcTempBus]          temp_m3_20_23_i;
wire signed [`CalcTempBus]          temp_m3_20_24_r;
wire signed [`CalcTempBus]          temp_m3_20_24_i;
wire signed [`CalcTempBus]          temp_m3_20_25_r;
wire signed [`CalcTempBus]          temp_m3_20_25_i;
wire signed [`CalcTempBus]          temp_m3_20_26_r;
wire signed [`CalcTempBus]          temp_m3_20_26_i;
wire signed [`CalcTempBus]          temp_m3_20_27_r;
wire signed [`CalcTempBus]          temp_m3_20_27_i;
wire signed [`CalcTempBus]          temp_m3_20_28_r;
wire signed [`CalcTempBus]          temp_m3_20_28_i;
wire signed [`CalcTempBus]          temp_m3_20_29_r;
wire signed [`CalcTempBus]          temp_m3_20_29_i;
wire signed [`CalcTempBus]          temp_m3_20_30_r;
wire signed [`CalcTempBus]          temp_m3_20_30_i;
wire signed [`CalcTempBus]          temp_m3_20_31_r;
wire signed [`CalcTempBus]          temp_m3_20_31_i;
wire signed [`CalcTempBus]          temp_m3_20_32_r;
wire signed [`CalcTempBus]          temp_m3_20_32_i;
wire signed [`CalcTempBus]          temp_m3_21_1_r;
wire signed [`CalcTempBus]          temp_m3_21_1_i;
wire signed [`CalcTempBus]          temp_m3_21_2_r;
wire signed [`CalcTempBus]          temp_m3_21_2_i;
wire signed [`CalcTempBus]          temp_m3_21_3_r;
wire signed [`CalcTempBus]          temp_m3_21_3_i;
wire signed [`CalcTempBus]          temp_m3_21_4_r;
wire signed [`CalcTempBus]          temp_m3_21_4_i;
wire signed [`CalcTempBus]          temp_m3_21_5_r;
wire signed [`CalcTempBus]          temp_m3_21_5_i;
wire signed [`CalcTempBus]          temp_m3_21_6_r;
wire signed [`CalcTempBus]          temp_m3_21_6_i;
wire signed [`CalcTempBus]          temp_m3_21_7_r;
wire signed [`CalcTempBus]          temp_m3_21_7_i;
wire signed [`CalcTempBus]          temp_m3_21_8_r;
wire signed [`CalcTempBus]          temp_m3_21_8_i;
wire signed [`CalcTempBus]          temp_m3_21_9_r;
wire signed [`CalcTempBus]          temp_m3_21_9_i;
wire signed [`CalcTempBus]          temp_m3_21_10_r;
wire signed [`CalcTempBus]          temp_m3_21_10_i;
wire signed [`CalcTempBus]          temp_m3_21_11_r;
wire signed [`CalcTempBus]          temp_m3_21_11_i;
wire signed [`CalcTempBus]          temp_m3_21_12_r;
wire signed [`CalcTempBus]          temp_m3_21_12_i;
wire signed [`CalcTempBus]          temp_m3_21_13_r;
wire signed [`CalcTempBus]          temp_m3_21_13_i;
wire signed [`CalcTempBus]          temp_m3_21_14_r;
wire signed [`CalcTempBus]          temp_m3_21_14_i;
wire signed [`CalcTempBus]          temp_m3_21_15_r;
wire signed [`CalcTempBus]          temp_m3_21_15_i;
wire signed [`CalcTempBus]          temp_m3_21_16_r;
wire signed [`CalcTempBus]          temp_m3_21_16_i;
wire signed [`CalcTempBus]          temp_m3_21_17_r;
wire signed [`CalcTempBus]          temp_m3_21_17_i;
wire signed [`CalcTempBus]          temp_m3_21_18_r;
wire signed [`CalcTempBus]          temp_m3_21_18_i;
wire signed [`CalcTempBus]          temp_m3_21_19_r;
wire signed [`CalcTempBus]          temp_m3_21_19_i;
wire signed [`CalcTempBus]          temp_m3_21_20_r;
wire signed [`CalcTempBus]          temp_m3_21_20_i;
wire signed [`CalcTempBus]          temp_m3_21_21_r;
wire signed [`CalcTempBus]          temp_m3_21_21_i;
wire signed [`CalcTempBus]          temp_m3_21_22_r;
wire signed [`CalcTempBus]          temp_m3_21_22_i;
wire signed [`CalcTempBus]          temp_m3_21_23_r;
wire signed [`CalcTempBus]          temp_m3_21_23_i;
wire signed [`CalcTempBus]          temp_m3_21_24_r;
wire signed [`CalcTempBus]          temp_m3_21_24_i;
wire signed [`CalcTempBus]          temp_m3_21_25_r;
wire signed [`CalcTempBus]          temp_m3_21_25_i;
wire signed [`CalcTempBus]          temp_m3_21_26_r;
wire signed [`CalcTempBus]          temp_m3_21_26_i;
wire signed [`CalcTempBus]          temp_m3_21_27_r;
wire signed [`CalcTempBus]          temp_m3_21_27_i;
wire signed [`CalcTempBus]          temp_m3_21_28_r;
wire signed [`CalcTempBus]          temp_m3_21_28_i;
wire signed [`CalcTempBus]          temp_m3_21_29_r;
wire signed [`CalcTempBus]          temp_m3_21_29_i;
wire signed [`CalcTempBus]          temp_m3_21_30_r;
wire signed [`CalcTempBus]          temp_m3_21_30_i;
wire signed [`CalcTempBus]          temp_m3_21_31_r;
wire signed [`CalcTempBus]          temp_m3_21_31_i;
wire signed [`CalcTempBus]          temp_m3_21_32_r;
wire signed [`CalcTempBus]          temp_m3_21_32_i;
wire signed [`CalcTempBus]          temp_m3_22_1_r;
wire signed [`CalcTempBus]          temp_m3_22_1_i;
wire signed [`CalcTempBus]          temp_m3_22_2_r;
wire signed [`CalcTempBus]          temp_m3_22_2_i;
wire signed [`CalcTempBus]          temp_m3_22_3_r;
wire signed [`CalcTempBus]          temp_m3_22_3_i;
wire signed [`CalcTempBus]          temp_m3_22_4_r;
wire signed [`CalcTempBus]          temp_m3_22_4_i;
wire signed [`CalcTempBus]          temp_m3_22_5_r;
wire signed [`CalcTempBus]          temp_m3_22_5_i;
wire signed [`CalcTempBus]          temp_m3_22_6_r;
wire signed [`CalcTempBus]          temp_m3_22_6_i;
wire signed [`CalcTempBus]          temp_m3_22_7_r;
wire signed [`CalcTempBus]          temp_m3_22_7_i;
wire signed [`CalcTempBus]          temp_m3_22_8_r;
wire signed [`CalcTempBus]          temp_m3_22_8_i;
wire signed [`CalcTempBus]          temp_m3_22_9_r;
wire signed [`CalcTempBus]          temp_m3_22_9_i;
wire signed [`CalcTempBus]          temp_m3_22_10_r;
wire signed [`CalcTempBus]          temp_m3_22_10_i;
wire signed [`CalcTempBus]          temp_m3_22_11_r;
wire signed [`CalcTempBus]          temp_m3_22_11_i;
wire signed [`CalcTempBus]          temp_m3_22_12_r;
wire signed [`CalcTempBus]          temp_m3_22_12_i;
wire signed [`CalcTempBus]          temp_m3_22_13_r;
wire signed [`CalcTempBus]          temp_m3_22_13_i;
wire signed [`CalcTempBus]          temp_m3_22_14_r;
wire signed [`CalcTempBus]          temp_m3_22_14_i;
wire signed [`CalcTempBus]          temp_m3_22_15_r;
wire signed [`CalcTempBus]          temp_m3_22_15_i;
wire signed [`CalcTempBus]          temp_m3_22_16_r;
wire signed [`CalcTempBus]          temp_m3_22_16_i;
wire signed [`CalcTempBus]          temp_m3_22_17_r;
wire signed [`CalcTempBus]          temp_m3_22_17_i;
wire signed [`CalcTempBus]          temp_m3_22_18_r;
wire signed [`CalcTempBus]          temp_m3_22_18_i;
wire signed [`CalcTempBus]          temp_m3_22_19_r;
wire signed [`CalcTempBus]          temp_m3_22_19_i;
wire signed [`CalcTempBus]          temp_m3_22_20_r;
wire signed [`CalcTempBus]          temp_m3_22_20_i;
wire signed [`CalcTempBus]          temp_m3_22_21_r;
wire signed [`CalcTempBus]          temp_m3_22_21_i;
wire signed [`CalcTempBus]          temp_m3_22_22_r;
wire signed [`CalcTempBus]          temp_m3_22_22_i;
wire signed [`CalcTempBus]          temp_m3_22_23_r;
wire signed [`CalcTempBus]          temp_m3_22_23_i;
wire signed [`CalcTempBus]          temp_m3_22_24_r;
wire signed [`CalcTempBus]          temp_m3_22_24_i;
wire signed [`CalcTempBus]          temp_m3_22_25_r;
wire signed [`CalcTempBus]          temp_m3_22_25_i;
wire signed [`CalcTempBus]          temp_m3_22_26_r;
wire signed [`CalcTempBus]          temp_m3_22_26_i;
wire signed [`CalcTempBus]          temp_m3_22_27_r;
wire signed [`CalcTempBus]          temp_m3_22_27_i;
wire signed [`CalcTempBus]          temp_m3_22_28_r;
wire signed [`CalcTempBus]          temp_m3_22_28_i;
wire signed [`CalcTempBus]          temp_m3_22_29_r;
wire signed [`CalcTempBus]          temp_m3_22_29_i;
wire signed [`CalcTempBus]          temp_m3_22_30_r;
wire signed [`CalcTempBus]          temp_m3_22_30_i;
wire signed [`CalcTempBus]          temp_m3_22_31_r;
wire signed [`CalcTempBus]          temp_m3_22_31_i;
wire signed [`CalcTempBus]          temp_m3_22_32_r;
wire signed [`CalcTempBus]          temp_m3_22_32_i;
wire signed [`CalcTempBus]          temp_m3_23_1_r;
wire signed [`CalcTempBus]          temp_m3_23_1_i;
wire signed [`CalcTempBus]          temp_m3_23_2_r;
wire signed [`CalcTempBus]          temp_m3_23_2_i;
wire signed [`CalcTempBus]          temp_m3_23_3_r;
wire signed [`CalcTempBus]          temp_m3_23_3_i;
wire signed [`CalcTempBus]          temp_m3_23_4_r;
wire signed [`CalcTempBus]          temp_m3_23_4_i;
wire signed [`CalcTempBus]          temp_m3_23_5_r;
wire signed [`CalcTempBus]          temp_m3_23_5_i;
wire signed [`CalcTempBus]          temp_m3_23_6_r;
wire signed [`CalcTempBus]          temp_m3_23_6_i;
wire signed [`CalcTempBus]          temp_m3_23_7_r;
wire signed [`CalcTempBus]          temp_m3_23_7_i;
wire signed [`CalcTempBus]          temp_m3_23_8_r;
wire signed [`CalcTempBus]          temp_m3_23_8_i;
wire signed [`CalcTempBus]          temp_m3_23_9_r;
wire signed [`CalcTempBus]          temp_m3_23_9_i;
wire signed [`CalcTempBus]          temp_m3_23_10_r;
wire signed [`CalcTempBus]          temp_m3_23_10_i;
wire signed [`CalcTempBus]          temp_m3_23_11_r;
wire signed [`CalcTempBus]          temp_m3_23_11_i;
wire signed [`CalcTempBus]          temp_m3_23_12_r;
wire signed [`CalcTempBus]          temp_m3_23_12_i;
wire signed [`CalcTempBus]          temp_m3_23_13_r;
wire signed [`CalcTempBus]          temp_m3_23_13_i;
wire signed [`CalcTempBus]          temp_m3_23_14_r;
wire signed [`CalcTempBus]          temp_m3_23_14_i;
wire signed [`CalcTempBus]          temp_m3_23_15_r;
wire signed [`CalcTempBus]          temp_m3_23_15_i;
wire signed [`CalcTempBus]          temp_m3_23_16_r;
wire signed [`CalcTempBus]          temp_m3_23_16_i;
wire signed [`CalcTempBus]          temp_m3_23_17_r;
wire signed [`CalcTempBus]          temp_m3_23_17_i;
wire signed [`CalcTempBus]          temp_m3_23_18_r;
wire signed [`CalcTempBus]          temp_m3_23_18_i;
wire signed [`CalcTempBus]          temp_m3_23_19_r;
wire signed [`CalcTempBus]          temp_m3_23_19_i;
wire signed [`CalcTempBus]          temp_m3_23_20_r;
wire signed [`CalcTempBus]          temp_m3_23_20_i;
wire signed [`CalcTempBus]          temp_m3_23_21_r;
wire signed [`CalcTempBus]          temp_m3_23_21_i;
wire signed [`CalcTempBus]          temp_m3_23_22_r;
wire signed [`CalcTempBus]          temp_m3_23_22_i;
wire signed [`CalcTempBus]          temp_m3_23_23_r;
wire signed [`CalcTempBus]          temp_m3_23_23_i;
wire signed [`CalcTempBus]          temp_m3_23_24_r;
wire signed [`CalcTempBus]          temp_m3_23_24_i;
wire signed [`CalcTempBus]          temp_m3_23_25_r;
wire signed [`CalcTempBus]          temp_m3_23_25_i;
wire signed [`CalcTempBus]          temp_m3_23_26_r;
wire signed [`CalcTempBus]          temp_m3_23_26_i;
wire signed [`CalcTempBus]          temp_m3_23_27_r;
wire signed [`CalcTempBus]          temp_m3_23_27_i;
wire signed [`CalcTempBus]          temp_m3_23_28_r;
wire signed [`CalcTempBus]          temp_m3_23_28_i;
wire signed [`CalcTempBus]          temp_m3_23_29_r;
wire signed [`CalcTempBus]          temp_m3_23_29_i;
wire signed [`CalcTempBus]          temp_m3_23_30_r;
wire signed [`CalcTempBus]          temp_m3_23_30_i;
wire signed [`CalcTempBus]          temp_m3_23_31_r;
wire signed [`CalcTempBus]          temp_m3_23_31_i;
wire signed [`CalcTempBus]          temp_m3_23_32_r;
wire signed [`CalcTempBus]          temp_m3_23_32_i;
wire signed [`CalcTempBus]          temp_m3_24_1_r;
wire signed [`CalcTempBus]          temp_m3_24_1_i;
wire signed [`CalcTempBus]          temp_m3_24_2_r;
wire signed [`CalcTempBus]          temp_m3_24_2_i;
wire signed [`CalcTempBus]          temp_m3_24_3_r;
wire signed [`CalcTempBus]          temp_m3_24_3_i;
wire signed [`CalcTempBus]          temp_m3_24_4_r;
wire signed [`CalcTempBus]          temp_m3_24_4_i;
wire signed [`CalcTempBus]          temp_m3_24_5_r;
wire signed [`CalcTempBus]          temp_m3_24_5_i;
wire signed [`CalcTempBus]          temp_m3_24_6_r;
wire signed [`CalcTempBus]          temp_m3_24_6_i;
wire signed [`CalcTempBus]          temp_m3_24_7_r;
wire signed [`CalcTempBus]          temp_m3_24_7_i;
wire signed [`CalcTempBus]          temp_m3_24_8_r;
wire signed [`CalcTempBus]          temp_m3_24_8_i;
wire signed [`CalcTempBus]          temp_m3_24_9_r;
wire signed [`CalcTempBus]          temp_m3_24_9_i;
wire signed [`CalcTempBus]          temp_m3_24_10_r;
wire signed [`CalcTempBus]          temp_m3_24_10_i;
wire signed [`CalcTempBus]          temp_m3_24_11_r;
wire signed [`CalcTempBus]          temp_m3_24_11_i;
wire signed [`CalcTempBus]          temp_m3_24_12_r;
wire signed [`CalcTempBus]          temp_m3_24_12_i;
wire signed [`CalcTempBus]          temp_m3_24_13_r;
wire signed [`CalcTempBus]          temp_m3_24_13_i;
wire signed [`CalcTempBus]          temp_m3_24_14_r;
wire signed [`CalcTempBus]          temp_m3_24_14_i;
wire signed [`CalcTempBus]          temp_m3_24_15_r;
wire signed [`CalcTempBus]          temp_m3_24_15_i;
wire signed [`CalcTempBus]          temp_m3_24_16_r;
wire signed [`CalcTempBus]          temp_m3_24_16_i;
wire signed [`CalcTempBus]          temp_m3_24_17_r;
wire signed [`CalcTempBus]          temp_m3_24_17_i;
wire signed [`CalcTempBus]          temp_m3_24_18_r;
wire signed [`CalcTempBus]          temp_m3_24_18_i;
wire signed [`CalcTempBus]          temp_m3_24_19_r;
wire signed [`CalcTempBus]          temp_m3_24_19_i;
wire signed [`CalcTempBus]          temp_m3_24_20_r;
wire signed [`CalcTempBus]          temp_m3_24_20_i;
wire signed [`CalcTempBus]          temp_m3_24_21_r;
wire signed [`CalcTempBus]          temp_m3_24_21_i;
wire signed [`CalcTempBus]          temp_m3_24_22_r;
wire signed [`CalcTempBus]          temp_m3_24_22_i;
wire signed [`CalcTempBus]          temp_m3_24_23_r;
wire signed [`CalcTempBus]          temp_m3_24_23_i;
wire signed [`CalcTempBus]          temp_m3_24_24_r;
wire signed [`CalcTempBus]          temp_m3_24_24_i;
wire signed [`CalcTempBus]          temp_m3_24_25_r;
wire signed [`CalcTempBus]          temp_m3_24_25_i;
wire signed [`CalcTempBus]          temp_m3_24_26_r;
wire signed [`CalcTempBus]          temp_m3_24_26_i;
wire signed [`CalcTempBus]          temp_m3_24_27_r;
wire signed [`CalcTempBus]          temp_m3_24_27_i;
wire signed [`CalcTempBus]          temp_m3_24_28_r;
wire signed [`CalcTempBus]          temp_m3_24_28_i;
wire signed [`CalcTempBus]          temp_m3_24_29_r;
wire signed [`CalcTempBus]          temp_m3_24_29_i;
wire signed [`CalcTempBus]          temp_m3_24_30_r;
wire signed [`CalcTempBus]          temp_m3_24_30_i;
wire signed [`CalcTempBus]          temp_m3_24_31_r;
wire signed [`CalcTempBus]          temp_m3_24_31_i;
wire signed [`CalcTempBus]          temp_m3_24_32_r;
wire signed [`CalcTempBus]          temp_m3_24_32_i;
wire signed [`CalcTempBus]          temp_m3_25_1_r;
wire signed [`CalcTempBus]          temp_m3_25_1_i;
wire signed [`CalcTempBus]          temp_m3_25_2_r;
wire signed [`CalcTempBus]          temp_m3_25_2_i;
wire signed [`CalcTempBus]          temp_m3_25_3_r;
wire signed [`CalcTempBus]          temp_m3_25_3_i;
wire signed [`CalcTempBus]          temp_m3_25_4_r;
wire signed [`CalcTempBus]          temp_m3_25_4_i;
wire signed [`CalcTempBus]          temp_m3_25_5_r;
wire signed [`CalcTempBus]          temp_m3_25_5_i;
wire signed [`CalcTempBus]          temp_m3_25_6_r;
wire signed [`CalcTempBus]          temp_m3_25_6_i;
wire signed [`CalcTempBus]          temp_m3_25_7_r;
wire signed [`CalcTempBus]          temp_m3_25_7_i;
wire signed [`CalcTempBus]          temp_m3_25_8_r;
wire signed [`CalcTempBus]          temp_m3_25_8_i;
wire signed [`CalcTempBus]          temp_m3_25_9_r;
wire signed [`CalcTempBus]          temp_m3_25_9_i;
wire signed [`CalcTempBus]          temp_m3_25_10_r;
wire signed [`CalcTempBus]          temp_m3_25_10_i;
wire signed [`CalcTempBus]          temp_m3_25_11_r;
wire signed [`CalcTempBus]          temp_m3_25_11_i;
wire signed [`CalcTempBus]          temp_m3_25_12_r;
wire signed [`CalcTempBus]          temp_m3_25_12_i;
wire signed [`CalcTempBus]          temp_m3_25_13_r;
wire signed [`CalcTempBus]          temp_m3_25_13_i;
wire signed [`CalcTempBus]          temp_m3_25_14_r;
wire signed [`CalcTempBus]          temp_m3_25_14_i;
wire signed [`CalcTempBus]          temp_m3_25_15_r;
wire signed [`CalcTempBus]          temp_m3_25_15_i;
wire signed [`CalcTempBus]          temp_m3_25_16_r;
wire signed [`CalcTempBus]          temp_m3_25_16_i;
wire signed [`CalcTempBus]          temp_m3_25_17_r;
wire signed [`CalcTempBus]          temp_m3_25_17_i;
wire signed [`CalcTempBus]          temp_m3_25_18_r;
wire signed [`CalcTempBus]          temp_m3_25_18_i;
wire signed [`CalcTempBus]          temp_m3_25_19_r;
wire signed [`CalcTempBus]          temp_m3_25_19_i;
wire signed [`CalcTempBus]          temp_m3_25_20_r;
wire signed [`CalcTempBus]          temp_m3_25_20_i;
wire signed [`CalcTempBus]          temp_m3_25_21_r;
wire signed [`CalcTempBus]          temp_m3_25_21_i;
wire signed [`CalcTempBus]          temp_m3_25_22_r;
wire signed [`CalcTempBus]          temp_m3_25_22_i;
wire signed [`CalcTempBus]          temp_m3_25_23_r;
wire signed [`CalcTempBus]          temp_m3_25_23_i;
wire signed [`CalcTempBus]          temp_m3_25_24_r;
wire signed [`CalcTempBus]          temp_m3_25_24_i;
wire signed [`CalcTempBus]          temp_m3_25_25_r;
wire signed [`CalcTempBus]          temp_m3_25_25_i;
wire signed [`CalcTempBus]          temp_m3_25_26_r;
wire signed [`CalcTempBus]          temp_m3_25_26_i;
wire signed [`CalcTempBus]          temp_m3_25_27_r;
wire signed [`CalcTempBus]          temp_m3_25_27_i;
wire signed [`CalcTempBus]          temp_m3_25_28_r;
wire signed [`CalcTempBus]          temp_m3_25_28_i;
wire signed [`CalcTempBus]          temp_m3_25_29_r;
wire signed [`CalcTempBus]          temp_m3_25_29_i;
wire signed [`CalcTempBus]          temp_m3_25_30_r;
wire signed [`CalcTempBus]          temp_m3_25_30_i;
wire signed [`CalcTempBus]          temp_m3_25_31_r;
wire signed [`CalcTempBus]          temp_m3_25_31_i;
wire signed [`CalcTempBus]          temp_m3_25_32_r;
wire signed [`CalcTempBus]          temp_m3_25_32_i;
wire signed [`CalcTempBus]          temp_m3_26_1_r;
wire signed [`CalcTempBus]          temp_m3_26_1_i;
wire signed [`CalcTempBus]          temp_m3_26_2_r;
wire signed [`CalcTempBus]          temp_m3_26_2_i;
wire signed [`CalcTempBus]          temp_m3_26_3_r;
wire signed [`CalcTempBus]          temp_m3_26_3_i;
wire signed [`CalcTempBus]          temp_m3_26_4_r;
wire signed [`CalcTempBus]          temp_m3_26_4_i;
wire signed [`CalcTempBus]          temp_m3_26_5_r;
wire signed [`CalcTempBus]          temp_m3_26_5_i;
wire signed [`CalcTempBus]          temp_m3_26_6_r;
wire signed [`CalcTempBus]          temp_m3_26_6_i;
wire signed [`CalcTempBus]          temp_m3_26_7_r;
wire signed [`CalcTempBus]          temp_m3_26_7_i;
wire signed [`CalcTempBus]          temp_m3_26_8_r;
wire signed [`CalcTempBus]          temp_m3_26_8_i;
wire signed [`CalcTempBus]          temp_m3_26_9_r;
wire signed [`CalcTempBus]          temp_m3_26_9_i;
wire signed [`CalcTempBus]          temp_m3_26_10_r;
wire signed [`CalcTempBus]          temp_m3_26_10_i;
wire signed [`CalcTempBus]          temp_m3_26_11_r;
wire signed [`CalcTempBus]          temp_m3_26_11_i;
wire signed [`CalcTempBus]          temp_m3_26_12_r;
wire signed [`CalcTempBus]          temp_m3_26_12_i;
wire signed [`CalcTempBus]          temp_m3_26_13_r;
wire signed [`CalcTempBus]          temp_m3_26_13_i;
wire signed [`CalcTempBus]          temp_m3_26_14_r;
wire signed [`CalcTempBus]          temp_m3_26_14_i;
wire signed [`CalcTempBus]          temp_m3_26_15_r;
wire signed [`CalcTempBus]          temp_m3_26_15_i;
wire signed [`CalcTempBus]          temp_m3_26_16_r;
wire signed [`CalcTempBus]          temp_m3_26_16_i;
wire signed [`CalcTempBus]          temp_m3_26_17_r;
wire signed [`CalcTempBus]          temp_m3_26_17_i;
wire signed [`CalcTempBus]          temp_m3_26_18_r;
wire signed [`CalcTempBus]          temp_m3_26_18_i;
wire signed [`CalcTempBus]          temp_m3_26_19_r;
wire signed [`CalcTempBus]          temp_m3_26_19_i;
wire signed [`CalcTempBus]          temp_m3_26_20_r;
wire signed [`CalcTempBus]          temp_m3_26_20_i;
wire signed [`CalcTempBus]          temp_m3_26_21_r;
wire signed [`CalcTempBus]          temp_m3_26_21_i;
wire signed [`CalcTempBus]          temp_m3_26_22_r;
wire signed [`CalcTempBus]          temp_m3_26_22_i;
wire signed [`CalcTempBus]          temp_m3_26_23_r;
wire signed [`CalcTempBus]          temp_m3_26_23_i;
wire signed [`CalcTempBus]          temp_m3_26_24_r;
wire signed [`CalcTempBus]          temp_m3_26_24_i;
wire signed [`CalcTempBus]          temp_m3_26_25_r;
wire signed [`CalcTempBus]          temp_m3_26_25_i;
wire signed [`CalcTempBus]          temp_m3_26_26_r;
wire signed [`CalcTempBus]          temp_m3_26_26_i;
wire signed [`CalcTempBus]          temp_m3_26_27_r;
wire signed [`CalcTempBus]          temp_m3_26_27_i;
wire signed [`CalcTempBus]          temp_m3_26_28_r;
wire signed [`CalcTempBus]          temp_m3_26_28_i;
wire signed [`CalcTempBus]          temp_m3_26_29_r;
wire signed [`CalcTempBus]          temp_m3_26_29_i;
wire signed [`CalcTempBus]          temp_m3_26_30_r;
wire signed [`CalcTempBus]          temp_m3_26_30_i;
wire signed [`CalcTempBus]          temp_m3_26_31_r;
wire signed [`CalcTempBus]          temp_m3_26_31_i;
wire signed [`CalcTempBus]          temp_m3_26_32_r;
wire signed [`CalcTempBus]          temp_m3_26_32_i;
wire signed [`CalcTempBus]          temp_m3_27_1_r;
wire signed [`CalcTempBus]          temp_m3_27_1_i;
wire signed [`CalcTempBus]          temp_m3_27_2_r;
wire signed [`CalcTempBus]          temp_m3_27_2_i;
wire signed [`CalcTempBus]          temp_m3_27_3_r;
wire signed [`CalcTempBus]          temp_m3_27_3_i;
wire signed [`CalcTempBus]          temp_m3_27_4_r;
wire signed [`CalcTempBus]          temp_m3_27_4_i;
wire signed [`CalcTempBus]          temp_m3_27_5_r;
wire signed [`CalcTempBus]          temp_m3_27_5_i;
wire signed [`CalcTempBus]          temp_m3_27_6_r;
wire signed [`CalcTempBus]          temp_m3_27_6_i;
wire signed [`CalcTempBus]          temp_m3_27_7_r;
wire signed [`CalcTempBus]          temp_m3_27_7_i;
wire signed [`CalcTempBus]          temp_m3_27_8_r;
wire signed [`CalcTempBus]          temp_m3_27_8_i;
wire signed [`CalcTempBus]          temp_m3_27_9_r;
wire signed [`CalcTempBus]          temp_m3_27_9_i;
wire signed [`CalcTempBus]          temp_m3_27_10_r;
wire signed [`CalcTempBus]          temp_m3_27_10_i;
wire signed [`CalcTempBus]          temp_m3_27_11_r;
wire signed [`CalcTempBus]          temp_m3_27_11_i;
wire signed [`CalcTempBus]          temp_m3_27_12_r;
wire signed [`CalcTempBus]          temp_m3_27_12_i;
wire signed [`CalcTempBus]          temp_m3_27_13_r;
wire signed [`CalcTempBus]          temp_m3_27_13_i;
wire signed [`CalcTempBus]          temp_m3_27_14_r;
wire signed [`CalcTempBus]          temp_m3_27_14_i;
wire signed [`CalcTempBus]          temp_m3_27_15_r;
wire signed [`CalcTempBus]          temp_m3_27_15_i;
wire signed [`CalcTempBus]          temp_m3_27_16_r;
wire signed [`CalcTempBus]          temp_m3_27_16_i;
wire signed [`CalcTempBus]          temp_m3_27_17_r;
wire signed [`CalcTempBus]          temp_m3_27_17_i;
wire signed [`CalcTempBus]          temp_m3_27_18_r;
wire signed [`CalcTempBus]          temp_m3_27_18_i;
wire signed [`CalcTempBus]          temp_m3_27_19_r;
wire signed [`CalcTempBus]          temp_m3_27_19_i;
wire signed [`CalcTempBus]          temp_m3_27_20_r;
wire signed [`CalcTempBus]          temp_m3_27_20_i;
wire signed [`CalcTempBus]          temp_m3_27_21_r;
wire signed [`CalcTempBus]          temp_m3_27_21_i;
wire signed [`CalcTempBus]          temp_m3_27_22_r;
wire signed [`CalcTempBus]          temp_m3_27_22_i;
wire signed [`CalcTempBus]          temp_m3_27_23_r;
wire signed [`CalcTempBus]          temp_m3_27_23_i;
wire signed [`CalcTempBus]          temp_m3_27_24_r;
wire signed [`CalcTempBus]          temp_m3_27_24_i;
wire signed [`CalcTempBus]          temp_m3_27_25_r;
wire signed [`CalcTempBus]          temp_m3_27_25_i;
wire signed [`CalcTempBus]          temp_m3_27_26_r;
wire signed [`CalcTempBus]          temp_m3_27_26_i;
wire signed [`CalcTempBus]          temp_m3_27_27_r;
wire signed [`CalcTempBus]          temp_m3_27_27_i;
wire signed [`CalcTempBus]          temp_m3_27_28_r;
wire signed [`CalcTempBus]          temp_m3_27_28_i;
wire signed [`CalcTempBus]          temp_m3_27_29_r;
wire signed [`CalcTempBus]          temp_m3_27_29_i;
wire signed [`CalcTempBus]          temp_m3_27_30_r;
wire signed [`CalcTempBus]          temp_m3_27_30_i;
wire signed [`CalcTempBus]          temp_m3_27_31_r;
wire signed [`CalcTempBus]          temp_m3_27_31_i;
wire signed [`CalcTempBus]          temp_m3_27_32_r;
wire signed [`CalcTempBus]          temp_m3_27_32_i;
wire signed [`CalcTempBus]          temp_m3_28_1_r;
wire signed [`CalcTempBus]          temp_m3_28_1_i;
wire signed [`CalcTempBus]          temp_m3_28_2_r;
wire signed [`CalcTempBus]          temp_m3_28_2_i;
wire signed [`CalcTempBus]          temp_m3_28_3_r;
wire signed [`CalcTempBus]          temp_m3_28_3_i;
wire signed [`CalcTempBus]          temp_m3_28_4_r;
wire signed [`CalcTempBus]          temp_m3_28_4_i;
wire signed [`CalcTempBus]          temp_m3_28_5_r;
wire signed [`CalcTempBus]          temp_m3_28_5_i;
wire signed [`CalcTempBus]          temp_m3_28_6_r;
wire signed [`CalcTempBus]          temp_m3_28_6_i;
wire signed [`CalcTempBus]          temp_m3_28_7_r;
wire signed [`CalcTempBus]          temp_m3_28_7_i;
wire signed [`CalcTempBus]          temp_m3_28_8_r;
wire signed [`CalcTempBus]          temp_m3_28_8_i;
wire signed [`CalcTempBus]          temp_m3_28_9_r;
wire signed [`CalcTempBus]          temp_m3_28_9_i;
wire signed [`CalcTempBus]          temp_m3_28_10_r;
wire signed [`CalcTempBus]          temp_m3_28_10_i;
wire signed [`CalcTempBus]          temp_m3_28_11_r;
wire signed [`CalcTempBus]          temp_m3_28_11_i;
wire signed [`CalcTempBus]          temp_m3_28_12_r;
wire signed [`CalcTempBus]          temp_m3_28_12_i;
wire signed [`CalcTempBus]          temp_m3_28_13_r;
wire signed [`CalcTempBus]          temp_m3_28_13_i;
wire signed [`CalcTempBus]          temp_m3_28_14_r;
wire signed [`CalcTempBus]          temp_m3_28_14_i;
wire signed [`CalcTempBus]          temp_m3_28_15_r;
wire signed [`CalcTempBus]          temp_m3_28_15_i;
wire signed [`CalcTempBus]          temp_m3_28_16_r;
wire signed [`CalcTempBus]          temp_m3_28_16_i;
wire signed [`CalcTempBus]          temp_m3_28_17_r;
wire signed [`CalcTempBus]          temp_m3_28_17_i;
wire signed [`CalcTempBus]          temp_m3_28_18_r;
wire signed [`CalcTempBus]          temp_m3_28_18_i;
wire signed [`CalcTempBus]          temp_m3_28_19_r;
wire signed [`CalcTempBus]          temp_m3_28_19_i;
wire signed [`CalcTempBus]          temp_m3_28_20_r;
wire signed [`CalcTempBus]          temp_m3_28_20_i;
wire signed [`CalcTempBus]          temp_m3_28_21_r;
wire signed [`CalcTempBus]          temp_m3_28_21_i;
wire signed [`CalcTempBus]          temp_m3_28_22_r;
wire signed [`CalcTempBus]          temp_m3_28_22_i;
wire signed [`CalcTempBus]          temp_m3_28_23_r;
wire signed [`CalcTempBus]          temp_m3_28_23_i;
wire signed [`CalcTempBus]          temp_m3_28_24_r;
wire signed [`CalcTempBus]          temp_m3_28_24_i;
wire signed [`CalcTempBus]          temp_m3_28_25_r;
wire signed [`CalcTempBus]          temp_m3_28_25_i;
wire signed [`CalcTempBus]          temp_m3_28_26_r;
wire signed [`CalcTempBus]          temp_m3_28_26_i;
wire signed [`CalcTempBus]          temp_m3_28_27_r;
wire signed [`CalcTempBus]          temp_m3_28_27_i;
wire signed [`CalcTempBus]          temp_m3_28_28_r;
wire signed [`CalcTempBus]          temp_m3_28_28_i;
wire signed [`CalcTempBus]          temp_m3_28_29_r;
wire signed [`CalcTempBus]          temp_m3_28_29_i;
wire signed [`CalcTempBus]          temp_m3_28_30_r;
wire signed [`CalcTempBus]          temp_m3_28_30_i;
wire signed [`CalcTempBus]          temp_m3_28_31_r;
wire signed [`CalcTempBus]          temp_m3_28_31_i;
wire signed [`CalcTempBus]          temp_m3_28_32_r;
wire signed [`CalcTempBus]          temp_m3_28_32_i;
wire signed [`CalcTempBus]          temp_m3_29_1_r;
wire signed [`CalcTempBus]          temp_m3_29_1_i;
wire signed [`CalcTempBus]          temp_m3_29_2_r;
wire signed [`CalcTempBus]          temp_m3_29_2_i;
wire signed [`CalcTempBus]          temp_m3_29_3_r;
wire signed [`CalcTempBus]          temp_m3_29_3_i;
wire signed [`CalcTempBus]          temp_m3_29_4_r;
wire signed [`CalcTempBus]          temp_m3_29_4_i;
wire signed [`CalcTempBus]          temp_m3_29_5_r;
wire signed [`CalcTempBus]          temp_m3_29_5_i;
wire signed [`CalcTempBus]          temp_m3_29_6_r;
wire signed [`CalcTempBus]          temp_m3_29_6_i;
wire signed [`CalcTempBus]          temp_m3_29_7_r;
wire signed [`CalcTempBus]          temp_m3_29_7_i;
wire signed [`CalcTempBus]          temp_m3_29_8_r;
wire signed [`CalcTempBus]          temp_m3_29_8_i;
wire signed [`CalcTempBus]          temp_m3_29_9_r;
wire signed [`CalcTempBus]          temp_m3_29_9_i;
wire signed [`CalcTempBus]          temp_m3_29_10_r;
wire signed [`CalcTempBus]          temp_m3_29_10_i;
wire signed [`CalcTempBus]          temp_m3_29_11_r;
wire signed [`CalcTempBus]          temp_m3_29_11_i;
wire signed [`CalcTempBus]          temp_m3_29_12_r;
wire signed [`CalcTempBus]          temp_m3_29_12_i;
wire signed [`CalcTempBus]          temp_m3_29_13_r;
wire signed [`CalcTempBus]          temp_m3_29_13_i;
wire signed [`CalcTempBus]          temp_m3_29_14_r;
wire signed [`CalcTempBus]          temp_m3_29_14_i;
wire signed [`CalcTempBus]          temp_m3_29_15_r;
wire signed [`CalcTempBus]          temp_m3_29_15_i;
wire signed [`CalcTempBus]          temp_m3_29_16_r;
wire signed [`CalcTempBus]          temp_m3_29_16_i;
wire signed [`CalcTempBus]          temp_m3_29_17_r;
wire signed [`CalcTempBus]          temp_m3_29_17_i;
wire signed [`CalcTempBus]          temp_m3_29_18_r;
wire signed [`CalcTempBus]          temp_m3_29_18_i;
wire signed [`CalcTempBus]          temp_m3_29_19_r;
wire signed [`CalcTempBus]          temp_m3_29_19_i;
wire signed [`CalcTempBus]          temp_m3_29_20_r;
wire signed [`CalcTempBus]          temp_m3_29_20_i;
wire signed [`CalcTempBus]          temp_m3_29_21_r;
wire signed [`CalcTempBus]          temp_m3_29_21_i;
wire signed [`CalcTempBus]          temp_m3_29_22_r;
wire signed [`CalcTempBus]          temp_m3_29_22_i;
wire signed [`CalcTempBus]          temp_m3_29_23_r;
wire signed [`CalcTempBus]          temp_m3_29_23_i;
wire signed [`CalcTempBus]          temp_m3_29_24_r;
wire signed [`CalcTempBus]          temp_m3_29_24_i;
wire signed [`CalcTempBus]          temp_m3_29_25_r;
wire signed [`CalcTempBus]          temp_m3_29_25_i;
wire signed [`CalcTempBus]          temp_m3_29_26_r;
wire signed [`CalcTempBus]          temp_m3_29_26_i;
wire signed [`CalcTempBus]          temp_m3_29_27_r;
wire signed [`CalcTempBus]          temp_m3_29_27_i;
wire signed [`CalcTempBus]          temp_m3_29_28_r;
wire signed [`CalcTempBus]          temp_m3_29_28_i;
wire signed [`CalcTempBus]          temp_m3_29_29_r;
wire signed [`CalcTempBus]          temp_m3_29_29_i;
wire signed [`CalcTempBus]          temp_m3_29_30_r;
wire signed [`CalcTempBus]          temp_m3_29_30_i;
wire signed [`CalcTempBus]          temp_m3_29_31_r;
wire signed [`CalcTempBus]          temp_m3_29_31_i;
wire signed [`CalcTempBus]          temp_m3_29_32_r;
wire signed [`CalcTempBus]          temp_m3_29_32_i;
wire signed [`CalcTempBus]          temp_m3_30_1_r;
wire signed [`CalcTempBus]          temp_m3_30_1_i;
wire signed [`CalcTempBus]          temp_m3_30_2_r;
wire signed [`CalcTempBus]          temp_m3_30_2_i;
wire signed [`CalcTempBus]          temp_m3_30_3_r;
wire signed [`CalcTempBus]          temp_m3_30_3_i;
wire signed [`CalcTempBus]          temp_m3_30_4_r;
wire signed [`CalcTempBus]          temp_m3_30_4_i;
wire signed [`CalcTempBus]          temp_m3_30_5_r;
wire signed [`CalcTempBus]          temp_m3_30_5_i;
wire signed [`CalcTempBus]          temp_m3_30_6_r;
wire signed [`CalcTempBus]          temp_m3_30_6_i;
wire signed [`CalcTempBus]          temp_m3_30_7_r;
wire signed [`CalcTempBus]          temp_m3_30_7_i;
wire signed [`CalcTempBus]          temp_m3_30_8_r;
wire signed [`CalcTempBus]          temp_m3_30_8_i;
wire signed [`CalcTempBus]          temp_m3_30_9_r;
wire signed [`CalcTempBus]          temp_m3_30_9_i;
wire signed [`CalcTempBus]          temp_m3_30_10_r;
wire signed [`CalcTempBus]          temp_m3_30_10_i;
wire signed [`CalcTempBus]          temp_m3_30_11_r;
wire signed [`CalcTempBus]          temp_m3_30_11_i;
wire signed [`CalcTempBus]          temp_m3_30_12_r;
wire signed [`CalcTempBus]          temp_m3_30_12_i;
wire signed [`CalcTempBus]          temp_m3_30_13_r;
wire signed [`CalcTempBus]          temp_m3_30_13_i;
wire signed [`CalcTempBus]          temp_m3_30_14_r;
wire signed [`CalcTempBus]          temp_m3_30_14_i;
wire signed [`CalcTempBus]          temp_m3_30_15_r;
wire signed [`CalcTempBus]          temp_m3_30_15_i;
wire signed [`CalcTempBus]          temp_m3_30_16_r;
wire signed [`CalcTempBus]          temp_m3_30_16_i;
wire signed [`CalcTempBus]          temp_m3_30_17_r;
wire signed [`CalcTempBus]          temp_m3_30_17_i;
wire signed [`CalcTempBus]          temp_m3_30_18_r;
wire signed [`CalcTempBus]          temp_m3_30_18_i;
wire signed [`CalcTempBus]          temp_m3_30_19_r;
wire signed [`CalcTempBus]          temp_m3_30_19_i;
wire signed [`CalcTempBus]          temp_m3_30_20_r;
wire signed [`CalcTempBus]          temp_m3_30_20_i;
wire signed [`CalcTempBus]          temp_m3_30_21_r;
wire signed [`CalcTempBus]          temp_m3_30_21_i;
wire signed [`CalcTempBus]          temp_m3_30_22_r;
wire signed [`CalcTempBus]          temp_m3_30_22_i;
wire signed [`CalcTempBus]          temp_m3_30_23_r;
wire signed [`CalcTempBus]          temp_m3_30_23_i;
wire signed [`CalcTempBus]          temp_m3_30_24_r;
wire signed [`CalcTempBus]          temp_m3_30_24_i;
wire signed [`CalcTempBus]          temp_m3_30_25_r;
wire signed [`CalcTempBus]          temp_m3_30_25_i;
wire signed [`CalcTempBus]          temp_m3_30_26_r;
wire signed [`CalcTempBus]          temp_m3_30_26_i;
wire signed [`CalcTempBus]          temp_m3_30_27_r;
wire signed [`CalcTempBus]          temp_m3_30_27_i;
wire signed [`CalcTempBus]          temp_m3_30_28_r;
wire signed [`CalcTempBus]          temp_m3_30_28_i;
wire signed [`CalcTempBus]          temp_m3_30_29_r;
wire signed [`CalcTempBus]          temp_m3_30_29_i;
wire signed [`CalcTempBus]          temp_m3_30_30_r;
wire signed [`CalcTempBus]          temp_m3_30_30_i;
wire signed [`CalcTempBus]          temp_m3_30_31_r;
wire signed [`CalcTempBus]          temp_m3_30_31_i;
wire signed [`CalcTempBus]          temp_m3_30_32_r;
wire signed [`CalcTempBus]          temp_m3_30_32_i;
wire signed [`CalcTempBus]          temp_m3_31_1_r;
wire signed [`CalcTempBus]          temp_m3_31_1_i;
wire signed [`CalcTempBus]          temp_m3_31_2_r;
wire signed [`CalcTempBus]          temp_m3_31_2_i;
wire signed [`CalcTempBus]          temp_m3_31_3_r;
wire signed [`CalcTempBus]          temp_m3_31_3_i;
wire signed [`CalcTempBus]          temp_m3_31_4_r;
wire signed [`CalcTempBus]          temp_m3_31_4_i;
wire signed [`CalcTempBus]          temp_m3_31_5_r;
wire signed [`CalcTempBus]          temp_m3_31_5_i;
wire signed [`CalcTempBus]          temp_m3_31_6_r;
wire signed [`CalcTempBus]          temp_m3_31_6_i;
wire signed [`CalcTempBus]          temp_m3_31_7_r;
wire signed [`CalcTempBus]          temp_m3_31_7_i;
wire signed [`CalcTempBus]          temp_m3_31_8_r;
wire signed [`CalcTempBus]          temp_m3_31_8_i;
wire signed [`CalcTempBus]          temp_m3_31_9_r;
wire signed [`CalcTempBus]          temp_m3_31_9_i;
wire signed [`CalcTempBus]          temp_m3_31_10_r;
wire signed [`CalcTempBus]          temp_m3_31_10_i;
wire signed [`CalcTempBus]          temp_m3_31_11_r;
wire signed [`CalcTempBus]          temp_m3_31_11_i;
wire signed [`CalcTempBus]          temp_m3_31_12_r;
wire signed [`CalcTempBus]          temp_m3_31_12_i;
wire signed [`CalcTempBus]          temp_m3_31_13_r;
wire signed [`CalcTempBus]          temp_m3_31_13_i;
wire signed [`CalcTempBus]          temp_m3_31_14_r;
wire signed [`CalcTempBus]          temp_m3_31_14_i;
wire signed [`CalcTempBus]          temp_m3_31_15_r;
wire signed [`CalcTempBus]          temp_m3_31_15_i;
wire signed [`CalcTempBus]          temp_m3_31_16_r;
wire signed [`CalcTempBus]          temp_m3_31_16_i;
wire signed [`CalcTempBus]          temp_m3_31_17_r;
wire signed [`CalcTempBus]          temp_m3_31_17_i;
wire signed [`CalcTempBus]          temp_m3_31_18_r;
wire signed [`CalcTempBus]          temp_m3_31_18_i;
wire signed [`CalcTempBus]          temp_m3_31_19_r;
wire signed [`CalcTempBus]          temp_m3_31_19_i;
wire signed [`CalcTempBus]          temp_m3_31_20_r;
wire signed [`CalcTempBus]          temp_m3_31_20_i;
wire signed [`CalcTempBus]          temp_m3_31_21_r;
wire signed [`CalcTempBus]          temp_m3_31_21_i;
wire signed [`CalcTempBus]          temp_m3_31_22_r;
wire signed [`CalcTempBus]          temp_m3_31_22_i;
wire signed [`CalcTempBus]          temp_m3_31_23_r;
wire signed [`CalcTempBus]          temp_m3_31_23_i;
wire signed [`CalcTempBus]          temp_m3_31_24_r;
wire signed [`CalcTempBus]          temp_m3_31_24_i;
wire signed [`CalcTempBus]          temp_m3_31_25_r;
wire signed [`CalcTempBus]          temp_m3_31_25_i;
wire signed [`CalcTempBus]          temp_m3_31_26_r;
wire signed [`CalcTempBus]          temp_m3_31_26_i;
wire signed [`CalcTempBus]          temp_m3_31_27_r;
wire signed [`CalcTempBus]          temp_m3_31_27_i;
wire signed [`CalcTempBus]          temp_m3_31_28_r;
wire signed [`CalcTempBus]          temp_m3_31_28_i;
wire signed [`CalcTempBus]          temp_m3_31_29_r;
wire signed [`CalcTempBus]          temp_m3_31_29_i;
wire signed [`CalcTempBus]          temp_m3_31_30_r;
wire signed [`CalcTempBus]          temp_m3_31_30_i;
wire signed [`CalcTempBus]          temp_m3_31_31_r;
wire signed [`CalcTempBus]          temp_m3_31_31_i;
wire signed [`CalcTempBus]          temp_m3_31_32_r;
wire signed [`CalcTempBus]          temp_m3_31_32_i;
wire signed [`CalcTempBus]          temp_m3_32_1_r;
wire signed [`CalcTempBus]          temp_m3_32_1_i;
wire signed [`CalcTempBus]          temp_m3_32_2_r;
wire signed [`CalcTempBus]          temp_m3_32_2_i;
wire signed [`CalcTempBus]          temp_m3_32_3_r;
wire signed [`CalcTempBus]          temp_m3_32_3_i;
wire signed [`CalcTempBus]          temp_m3_32_4_r;
wire signed [`CalcTempBus]          temp_m3_32_4_i;
wire signed [`CalcTempBus]          temp_m3_32_5_r;
wire signed [`CalcTempBus]          temp_m3_32_5_i;
wire signed [`CalcTempBus]          temp_m3_32_6_r;
wire signed [`CalcTempBus]          temp_m3_32_6_i;
wire signed [`CalcTempBus]          temp_m3_32_7_r;
wire signed [`CalcTempBus]          temp_m3_32_7_i;
wire signed [`CalcTempBus]          temp_m3_32_8_r;
wire signed [`CalcTempBus]          temp_m3_32_8_i;
wire signed [`CalcTempBus]          temp_m3_32_9_r;
wire signed [`CalcTempBus]          temp_m3_32_9_i;
wire signed [`CalcTempBus]          temp_m3_32_10_r;
wire signed [`CalcTempBus]          temp_m3_32_10_i;
wire signed [`CalcTempBus]          temp_m3_32_11_r;
wire signed [`CalcTempBus]          temp_m3_32_11_i;
wire signed [`CalcTempBus]          temp_m3_32_12_r;
wire signed [`CalcTempBus]          temp_m3_32_12_i;
wire signed [`CalcTempBus]          temp_m3_32_13_r;
wire signed [`CalcTempBus]          temp_m3_32_13_i;
wire signed [`CalcTempBus]          temp_m3_32_14_r;
wire signed [`CalcTempBus]          temp_m3_32_14_i;
wire signed [`CalcTempBus]          temp_m3_32_15_r;
wire signed [`CalcTempBus]          temp_m3_32_15_i;
wire signed [`CalcTempBus]          temp_m3_32_16_r;
wire signed [`CalcTempBus]          temp_m3_32_16_i;
wire signed [`CalcTempBus]          temp_m3_32_17_r;
wire signed [`CalcTempBus]          temp_m3_32_17_i;
wire signed [`CalcTempBus]          temp_m3_32_18_r;
wire signed [`CalcTempBus]          temp_m3_32_18_i;
wire signed [`CalcTempBus]          temp_m3_32_19_r;
wire signed [`CalcTempBus]          temp_m3_32_19_i;
wire signed [`CalcTempBus]          temp_m3_32_20_r;
wire signed [`CalcTempBus]          temp_m3_32_20_i;
wire signed [`CalcTempBus]          temp_m3_32_21_r;
wire signed [`CalcTempBus]          temp_m3_32_21_i;
wire signed [`CalcTempBus]          temp_m3_32_22_r;
wire signed [`CalcTempBus]          temp_m3_32_22_i;
wire signed [`CalcTempBus]          temp_m3_32_23_r;
wire signed [`CalcTempBus]          temp_m3_32_23_i;
wire signed [`CalcTempBus]          temp_m3_32_24_r;
wire signed [`CalcTempBus]          temp_m3_32_24_i;
wire signed [`CalcTempBus]          temp_m3_32_25_r;
wire signed [`CalcTempBus]          temp_m3_32_25_i;
wire signed [`CalcTempBus]          temp_m3_32_26_r;
wire signed [`CalcTempBus]          temp_m3_32_26_i;
wire signed [`CalcTempBus]          temp_m3_32_27_r;
wire signed [`CalcTempBus]          temp_m3_32_27_i;
wire signed [`CalcTempBus]          temp_m3_32_28_r;
wire signed [`CalcTempBus]          temp_m3_32_28_i;
wire signed [`CalcTempBus]          temp_m3_32_29_r;
wire signed [`CalcTempBus]          temp_m3_32_29_i;
wire signed [`CalcTempBus]          temp_m3_32_30_r;
wire signed [`CalcTempBus]          temp_m3_32_30_i;
wire signed [`CalcTempBus]          temp_m3_32_31_r;
wire signed [`CalcTempBus]          temp_m3_32_31_i;
wire signed [`CalcTempBus]          temp_m3_32_32_r;
wire signed [`CalcTempBus]          temp_m3_32_32_i;
wire signed [`CalcTempBus]          temp_m4_1_1_r;
wire signed [`CalcTempBus]          temp_m4_1_1_i;
wire signed [`CalcTempBus]          temp_m4_1_2_r;
wire signed [`CalcTempBus]          temp_m4_1_2_i;
wire signed [`CalcTempBus]          temp_m4_1_3_r;
wire signed [`CalcTempBus]          temp_m4_1_3_i;
wire signed [`CalcTempBus]          temp_m4_1_4_r;
wire signed [`CalcTempBus]          temp_m4_1_4_i;
wire signed [`CalcTempBus]          temp_m4_1_5_r;
wire signed [`CalcTempBus]          temp_m4_1_5_i;
wire signed [`CalcTempBus]          temp_m4_1_6_r;
wire signed [`CalcTempBus]          temp_m4_1_6_i;
wire signed [`CalcTempBus]          temp_m4_1_7_r;
wire signed [`CalcTempBus]          temp_m4_1_7_i;
wire signed [`CalcTempBus]          temp_m4_1_8_r;
wire signed [`CalcTempBus]          temp_m4_1_8_i;
wire signed [`CalcTempBus]          temp_m4_1_9_r;
wire signed [`CalcTempBus]          temp_m4_1_9_i;
wire signed [`CalcTempBus]          temp_m4_1_10_r;
wire signed [`CalcTempBus]          temp_m4_1_10_i;
wire signed [`CalcTempBus]          temp_m4_1_11_r;
wire signed [`CalcTempBus]          temp_m4_1_11_i;
wire signed [`CalcTempBus]          temp_m4_1_12_r;
wire signed [`CalcTempBus]          temp_m4_1_12_i;
wire signed [`CalcTempBus]          temp_m4_1_13_r;
wire signed [`CalcTempBus]          temp_m4_1_13_i;
wire signed [`CalcTempBus]          temp_m4_1_14_r;
wire signed [`CalcTempBus]          temp_m4_1_14_i;
wire signed [`CalcTempBus]          temp_m4_1_15_r;
wire signed [`CalcTempBus]          temp_m4_1_15_i;
wire signed [`CalcTempBus]          temp_m4_1_16_r;
wire signed [`CalcTempBus]          temp_m4_1_16_i;
wire signed [`CalcTempBus]          temp_m4_1_17_r;
wire signed [`CalcTempBus]          temp_m4_1_17_i;
wire signed [`CalcTempBus]          temp_m4_1_18_r;
wire signed [`CalcTempBus]          temp_m4_1_18_i;
wire signed [`CalcTempBus]          temp_m4_1_19_r;
wire signed [`CalcTempBus]          temp_m4_1_19_i;
wire signed [`CalcTempBus]          temp_m4_1_20_r;
wire signed [`CalcTempBus]          temp_m4_1_20_i;
wire signed [`CalcTempBus]          temp_m4_1_21_r;
wire signed [`CalcTempBus]          temp_m4_1_21_i;
wire signed [`CalcTempBus]          temp_m4_1_22_r;
wire signed [`CalcTempBus]          temp_m4_1_22_i;
wire signed [`CalcTempBus]          temp_m4_1_23_r;
wire signed [`CalcTempBus]          temp_m4_1_23_i;
wire signed [`CalcTempBus]          temp_m4_1_24_r;
wire signed [`CalcTempBus]          temp_m4_1_24_i;
wire signed [`CalcTempBus]          temp_m4_1_25_r;
wire signed [`CalcTempBus]          temp_m4_1_25_i;
wire signed [`CalcTempBus]          temp_m4_1_26_r;
wire signed [`CalcTempBus]          temp_m4_1_26_i;
wire signed [`CalcTempBus]          temp_m4_1_27_r;
wire signed [`CalcTempBus]          temp_m4_1_27_i;
wire signed [`CalcTempBus]          temp_m4_1_28_r;
wire signed [`CalcTempBus]          temp_m4_1_28_i;
wire signed [`CalcTempBus]          temp_m4_1_29_r;
wire signed [`CalcTempBus]          temp_m4_1_29_i;
wire signed [`CalcTempBus]          temp_m4_1_30_r;
wire signed [`CalcTempBus]          temp_m4_1_30_i;
wire signed [`CalcTempBus]          temp_m4_1_31_r;
wire signed [`CalcTempBus]          temp_m4_1_31_i;
wire signed [`CalcTempBus]          temp_m4_1_32_r;
wire signed [`CalcTempBus]          temp_m4_1_32_i;
wire signed [`CalcTempBus]          temp_m4_2_1_r;
wire signed [`CalcTempBus]          temp_m4_2_1_i;
wire signed [`CalcTempBus]          temp_m4_2_2_r;
wire signed [`CalcTempBus]          temp_m4_2_2_i;
wire signed [`CalcTempBus]          temp_m4_2_3_r;
wire signed [`CalcTempBus]          temp_m4_2_3_i;
wire signed [`CalcTempBus]          temp_m4_2_4_r;
wire signed [`CalcTempBus]          temp_m4_2_4_i;
wire signed [`CalcTempBus]          temp_m4_2_5_r;
wire signed [`CalcTempBus]          temp_m4_2_5_i;
wire signed [`CalcTempBus]          temp_m4_2_6_r;
wire signed [`CalcTempBus]          temp_m4_2_6_i;
wire signed [`CalcTempBus]          temp_m4_2_7_r;
wire signed [`CalcTempBus]          temp_m4_2_7_i;
wire signed [`CalcTempBus]          temp_m4_2_8_r;
wire signed [`CalcTempBus]          temp_m4_2_8_i;
wire signed [`CalcTempBus]          temp_m4_2_9_r;
wire signed [`CalcTempBus]          temp_m4_2_9_i;
wire signed [`CalcTempBus]          temp_m4_2_10_r;
wire signed [`CalcTempBus]          temp_m4_2_10_i;
wire signed [`CalcTempBus]          temp_m4_2_11_r;
wire signed [`CalcTempBus]          temp_m4_2_11_i;
wire signed [`CalcTempBus]          temp_m4_2_12_r;
wire signed [`CalcTempBus]          temp_m4_2_12_i;
wire signed [`CalcTempBus]          temp_m4_2_13_r;
wire signed [`CalcTempBus]          temp_m4_2_13_i;
wire signed [`CalcTempBus]          temp_m4_2_14_r;
wire signed [`CalcTempBus]          temp_m4_2_14_i;
wire signed [`CalcTempBus]          temp_m4_2_15_r;
wire signed [`CalcTempBus]          temp_m4_2_15_i;
wire signed [`CalcTempBus]          temp_m4_2_16_r;
wire signed [`CalcTempBus]          temp_m4_2_16_i;
wire signed [`CalcTempBus]          temp_m4_2_17_r;
wire signed [`CalcTempBus]          temp_m4_2_17_i;
wire signed [`CalcTempBus]          temp_m4_2_18_r;
wire signed [`CalcTempBus]          temp_m4_2_18_i;
wire signed [`CalcTempBus]          temp_m4_2_19_r;
wire signed [`CalcTempBus]          temp_m4_2_19_i;
wire signed [`CalcTempBus]          temp_m4_2_20_r;
wire signed [`CalcTempBus]          temp_m4_2_20_i;
wire signed [`CalcTempBus]          temp_m4_2_21_r;
wire signed [`CalcTempBus]          temp_m4_2_21_i;
wire signed [`CalcTempBus]          temp_m4_2_22_r;
wire signed [`CalcTempBus]          temp_m4_2_22_i;
wire signed [`CalcTempBus]          temp_m4_2_23_r;
wire signed [`CalcTempBus]          temp_m4_2_23_i;
wire signed [`CalcTempBus]          temp_m4_2_24_r;
wire signed [`CalcTempBus]          temp_m4_2_24_i;
wire signed [`CalcTempBus]          temp_m4_2_25_r;
wire signed [`CalcTempBus]          temp_m4_2_25_i;
wire signed [`CalcTempBus]          temp_m4_2_26_r;
wire signed [`CalcTempBus]          temp_m4_2_26_i;
wire signed [`CalcTempBus]          temp_m4_2_27_r;
wire signed [`CalcTempBus]          temp_m4_2_27_i;
wire signed [`CalcTempBus]          temp_m4_2_28_r;
wire signed [`CalcTempBus]          temp_m4_2_28_i;
wire signed [`CalcTempBus]          temp_m4_2_29_r;
wire signed [`CalcTempBus]          temp_m4_2_29_i;
wire signed [`CalcTempBus]          temp_m4_2_30_r;
wire signed [`CalcTempBus]          temp_m4_2_30_i;
wire signed [`CalcTempBus]          temp_m4_2_31_r;
wire signed [`CalcTempBus]          temp_m4_2_31_i;
wire signed [`CalcTempBus]          temp_m4_2_32_r;
wire signed [`CalcTempBus]          temp_m4_2_32_i;
wire signed [`CalcTempBus]          temp_m4_3_1_r;
wire signed [`CalcTempBus]          temp_m4_3_1_i;
wire signed [`CalcTempBus]          temp_m4_3_2_r;
wire signed [`CalcTempBus]          temp_m4_3_2_i;
wire signed [`CalcTempBus]          temp_m4_3_3_r;
wire signed [`CalcTempBus]          temp_m4_3_3_i;
wire signed [`CalcTempBus]          temp_m4_3_4_r;
wire signed [`CalcTempBus]          temp_m4_3_4_i;
wire signed [`CalcTempBus]          temp_m4_3_5_r;
wire signed [`CalcTempBus]          temp_m4_3_5_i;
wire signed [`CalcTempBus]          temp_m4_3_6_r;
wire signed [`CalcTempBus]          temp_m4_3_6_i;
wire signed [`CalcTempBus]          temp_m4_3_7_r;
wire signed [`CalcTempBus]          temp_m4_3_7_i;
wire signed [`CalcTempBus]          temp_m4_3_8_r;
wire signed [`CalcTempBus]          temp_m4_3_8_i;
wire signed [`CalcTempBus]          temp_m4_3_9_r;
wire signed [`CalcTempBus]          temp_m4_3_9_i;
wire signed [`CalcTempBus]          temp_m4_3_10_r;
wire signed [`CalcTempBus]          temp_m4_3_10_i;
wire signed [`CalcTempBus]          temp_m4_3_11_r;
wire signed [`CalcTempBus]          temp_m4_3_11_i;
wire signed [`CalcTempBus]          temp_m4_3_12_r;
wire signed [`CalcTempBus]          temp_m4_3_12_i;
wire signed [`CalcTempBus]          temp_m4_3_13_r;
wire signed [`CalcTempBus]          temp_m4_3_13_i;
wire signed [`CalcTempBus]          temp_m4_3_14_r;
wire signed [`CalcTempBus]          temp_m4_3_14_i;
wire signed [`CalcTempBus]          temp_m4_3_15_r;
wire signed [`CalcTempBus]          temp_m4_3_15_i;
wire signed [`CalcTempBus]          temp_m4_3_16_r;
wire signed [`CalcTempBus]          temp_m4_3_16_i;
wire signed [`CalcTempBus]          temp_m4_3_17_r;
wire signed [`CalcTempBus]          temp_m4_3_17_i;
wire signed [`CalcTempBus]          temp_m4_3_18_r;
wire signed [`CalcTempBus]          temp_m4_3_18_i;
wire signed [`CalcTempBus]          temp_m4_3_19_r;
wire signed [`CalcTempBus]          temp_m4_3_19_i;
wire signed [`CalcTempBus]          temp_m4_3_20_r;
wire signed [`CalcTempBus]          temp_m4_3_20_i;
wire signed [`CalcTempBus]          temp_m4_3_21_r;
wire signed [`CalcTempBus]          temp_m4_3_21_i;
wire signed [`CalcTempBus]          temp_m4_3_22_r;
wire signed [`CalcTempBus]          temp_m4_3_22_i;
wire signed [`CalcTempBus]          temp_m4_3_23_r;
wire signed [`CalcTempBus]          temp_m4_3_23_i;
wire signed [`CalcTempBus]          temp_m4_3_24_r;
wire signed [`CalcTempBus]          temp_m4_3_24_i;
wire signed [`CalcTempBus]          temp_m4_3_25_r;
wire signed [`CalcTempBus]          temp_m4_3_25_i;
wire signed [`CalcTempBus]          temp_m4_3_26_r;
wire signed [`CalcTempBus]          temp_m4_3_26_i;
wire signed [`CalcTempBus]          temp_m4_3_27_r;
wire signed [`CalcTempBus]          temp_m4_3_27_i;
wire signed [`CalcTempBus]          temp_m4_3_28_r;
wire signed [`CalcTempBus]          temp_m4_3_28_i;
wire signed [`CalcTempBus]          temp_m4_3_29_r;
wire signed [`CalcTempBus]          temp_m4_3_29_i;
wire signed [`CalcTempBus]          temp_m4_3_30_r;
wire signed [`CalcTempBus]          temp_m4_3_30_i;
wire signed [`CalcTempBus]          temp_m4_3_31_r;
wire signed [`CalcTempBus]          temp_m4_3_31_i;
wire signed [`CalcTempBus]          temp_m4_3_32_r;
wire signed [`CalcTempBus]          temp_m4_3_32_i;
wire signed [`CalcTempBus]          temp_m4_4_1_r;
wire signed [`CalcTempBus]          temp_m4_4_1_i;
wire signed [`CalcTempBus]          temp_m4_4_2_r;
wire signed [`CalcTempBus]          temp_m4_4_2_i;
wire signed [`CalcTempBus]          temp_m4_4_3_r;
wire signed [`CalcTempBus]          temp_m4_4_3_i;
wire signed [`CalcTempBus]          temp_m4_4_4_r;
wire signed [`CalcTempBus]          temp_m4_4_4_i;
wire signed [`CalcTempBus]          temp_m4_4_5_r;
wire signed [`CalcTempBus]          temp_m4_4_5_i;
wire signed [`CalcTempBus]          temp_m4_4_6_r;
wire signed [`CalcTempBus]          temp_m4_4_6_i;
wire signed [`CalcTempBus]          temp_m4_4_7_r;
wire signed [`CalcTempBus]          temp_m4_4_7_i;
wire signed [`CalcTempBus]          temp_m4_4_8_r;
wire signed [`CalcTempBus]          temp_m4_4_8_i;
wire signed [`CalcTempBus]          temp_m4_4_9_r;
wire signed [`CalcTempBus]          temp_m4_4_9_i;
wire signed [`CalcTempBus]          temp_m4_4_10_r;
wire signed [`CalcTempBus]          temp_m4_4_10_i;
wire signed [`CalcTempBus]          temp_m4_4_11_r;
wire signed [`CalcTempBus]          temp_m4_4_11_i;
wire signed [`CalcTempBus]          temp_m4_4_12_r;
wire signed [`CalcTempBus]          temp_m4_4_12_i;
wire signed [`CalcTempBus]          temp_m4_4_13_r;
wire signed [`CalcTempBus]          temp_m4_4_13_i;
wire signed [`CalcTempBus]          temp_m4_4_14_r;
wire signed [`CalcTempBus]          temp_m4_4_14_i;
wire signed [`CalcTempBus]          temp_m4_4_15_r;
wire signed [`CalcTempBus]          temp_m4_4_15_i;
wire signed [`CalcTempBus]          temp_m4_4_16_r;
wire signed [`CalcTempBus]          temp_m4_4_16_i;
wire signed [`CalcTempBus]          temp_m4_4_17_r;
wire signed [`CalcTempBus]          temp_m4_4_17_i;
wire signed [`CalcTempBus]          temp_m4_4_18_r;
wire signed [`CalcTempBus]          temp_m4_4_18_i;
wire signed [`CalcTempBus]          temp_m4_4_19_r;
wire signed [`CalcTempBus]          temp_m4_4_19_i;
wire signed [`CalcTempBus]          temp_m4_4_20_r;
wire signed [`CalcTempBus]          temp_m4_4_20_i;
wire signed [`CalcTempBus]          temp_m4_4_21_r;
wire signed [`CalcTempBus]          temp_m4_4_21_i;
wire signed [`CalcTempBus]          temp_m4_4_22_r;
wire signed [`CalcTempBus]          temp_m4_4_22_i;
wire signed [`CalcTempBus]          temp_m4_4_23_r;
wire signed [`CalcTempBus]          temp_m4_4_23_i;
wire signed [`CalcTempBus]          temp_m4_4_24_r;
wire signed [`CalcTempBus]          temp_m4_4_24_i;
wire signed [`CalcTempBus]          temp_m4_4_25_r;
wire signed [`CalcTempBus]          temp_m4_4_25_i;
wire signed [`CalcTempBus]          temp_m4_4_26_r;
wire signed [`CalcTempBus]          temp_m4_4_26_i;
wire signed [`CalcTempBus]          temp_m4_4_27_r;
wire signed [`CalcTempBus]          temp_m4_4_27_i;
wire signed [`CalcTempBus]          temp_m4_4_28_r;
wire signed [`CalcTempBus]          temp_m4_4_28_i;
wire signed [`CalcTempBus]          temp_m4_4_29_r;
wire signed [`CalcTempBus]          temp_m4_4_29_i;
wire signed [`CalcTempBus]          temp_m4_4_30_r;
wire signed [`CalcTempBus]          temp_m4_4_30_i;
wire signed [`CalcTempBus]          temp_m4_4_31_r;
wire signed [`CalcTempBus]          temp_m4_4_31_i;
wire signed [`CalcTempBus]          temp_m4_4_32_r;
wire signed [`CalcTempBus]          temp_m4_4_32_i;
wire signed [`CalcTempBus]          temp_m4_5_1_r;
wire signed [`CalcTempBus]          temp_m4_5_1_i;
wire signed [`CalcTempBus]          temp_m4_5_2_r;
wire signed [`CalcTempBus]          temp_m4_5_2_i;
wire signed [`CalcTempBus]          temp_m4_5_3_r;
wire signed [`CalcTempBus]          temp_m4_5_3_i;
wire signed [`CalcTempBus]          temp_m4_5_4_r;
wire signed [`CalcTempBus]          temp_m4_5_4_i;
wire signed [`CalcTempBus]          temp_m4_5_5_r;
wire signed [`CalcTempBus]          temp_m4_5_5_i;
wire signed [`CalcTempBus]          temp_m4_5_6_r;
wire signed [`CalcTempBus]          temp_m4_5_6_i;
wire signed [`CalcTempBus]          temp_m4_5_7_r;
wire signed [`CalcTempBus]          temp_m4_5_7_i;
wire signed [`CalcTempBus]          temp_m4_5_8_r;
wire signed [`CalcTempBus]          temp_m4_5_8_i;
wire signed [`CalcTempBus]          temp_m4_5_9_r;
wire signed [`CalcTempBus]          temp_m4_5_9_i;
wire signed [`CalcTempBus]          temp_m4_5_10_r;
wire signed [`CalcTempBus]          temp_m4_5_10_i;
wire signed [`CalcTempBus]          temp_m4_5_11_r;
wire signed [`CalcTempBus]          temp_m4_5_11_i;
wire signed [`CalcTempBus]          temp_m4_5_12_r;
wire signed [`CalcTempBus]          temp_m4_5_12_i;
wire signed [`CalcTempBus]          temp_m4_5_13_r;
wire signed [`CalcTempBus]          temp_m4_5_13_i;
wire signed [`CalcTempBus]          temp_m4_5_14_r;
wire signed [`CalcTempBus]          temp_m4_5_14_i;
wire signed [`CalcTempBus]          temp_m4_5_15_r;
wire signed [`CalcTempBus]          temp_m4_5_15_i;
wire signed [`CalcTempBus]          temp_m4_5_16_r;
wire signed [`CalcTempBus]          temp_m4_5_16_i;
wire signed [`CalcTempBus]          temp_m4_5_17_r;
wire signed [`CalcTempBus]          temp_m4_5_17_i;
wire signed [`CalcTempBus]          temp_m4_5_18_r;
wire signed [`CalcTempBus]          temp_m4_5_18_i;
wire signed [`CalcTempBus]          temp_m4_5_19_r;
wire signed [`CalcTempBus]          temp_m4_5_19_i;
wire signed [`CalcTempBus]          temp_m4_5_20_r;
wire signed [`CalcTempBus]          temp_m4_5_20_i;
wire signed [`CalcTempBus]          temp_m4_5_21_r;
wire signed [`CalcTempBus]          temp_m4_5_21_i;
wire signed [`CalcTempBus]          temp_m4_5_22_r;
wire signed [`CalcTempBus]          temp_m4_5_22_i;
wire signed [`CalcTempBus]          temp_m4_5_23_r;
wire signed [`CalcTempBus]          temp_m4_5_23_i;
wire signed [`CalcTempBus]          temp_m4_5_24_r;
wire signed [`CalcTempBus]          temp_m4_5_24_i;
wire signed [`CalcTempBus]          temp_m4_5_25_r;
wire signed [`CalcTempBus]          temp_m4_5_25_i;
wire signed [`CalcTempBus]          temp_m4_5_26_r;
wire signed [`CalcTempBus]          temp_m4_5_26_i;
wire signed [`CalcTempBus]          temp_m4_5_27_r;
wire signed [`CalcTempBus]          temp_m4_5_27_i;
wire signed [`CalcTempBus]          temp_m4_5_28_r;
wire signed [`CalcTempBus]          temp_m4_5_28_i;
wire signed [`CalcTempBus]          temp_m4_5_29_r;
wire signed [`CalcTempBus]          temp_m4_5_29_i;
wire signed [`CalcTempBus]          temp_m4_5_30_r;
wire signed [`CalcTempBus]          temp_m4_5_30_i;
wire signed [`CalcTempBus]          temp_m4_5_31_r;
wire signed [`CalcTempBus]          temp_m4_5_31_i;
wire signed [`CalcTempBus]          temp_m4_5_32_r;
wire signed [`CalcTempBus]          temp_m4_5_32_i;
wire signed [`CalcTempBus]          temp_m4_6_1_r;
wire signed [`CalcTempBus]          temp_m4_6_1_i;
wire signed [`CalcTempBus]          temp_m4_6_2_r;
wire signed [`CalcTempBus]          temp_m4_6_2_i;
wire signed [`CalcTempBus]          temp_m4_6_3_r;
wire signed [`CalcTempBus]          temp_m4_6_3_i;
wire signed [`CalcTempBus]          temp_m4_6_4_r;
wire signed [`CalcTempBus]          temp_m4_6_4_i;
wire signed [`CalcTempBus]          temp_m4_6_5_r;
wire signed [`CalcTempBus]          temp_m4_6_5_i;
wire signed [`CalcTempBus]          temp_m4_6_6_r;
wire signed [`CalcTempBus]          temp_m4_6_6_i;
wire signed [`CalcTempBus]          temp_m4_6_7_r;
wire signed [`CalcTempBus]          temp_m4_6_7_i;
wire signed [`CalcTempBus]          temp_m4_6_8_r;
wire signed [`CalcTempBus]          temp_m4_6_8_i;
wire signed [`CalcTempBus]          temp_m4_6_9_r;
wire signed [`CalcTempBus]          temp_m4_6_9_i;
wire signed [`CalcTempBus]          temp_m4_6_10_r;
wire signed [`CalcTempBus]          temp_m4_6_10_i;
wire signed [`CalcTempBus]          temp_m4_6_11_r;
wire signed [`CalcTempBus]          temp_m4_6_11_i;
wire signed [`CalcTempBus]          temp_m4_6_12_r;
wire signed [`CalcTempBus]          temp_m4_6_12_i;
wire signed [`CalcTempBus]          temp_m4_6_13_r;
wire signed [`CalcTempBus]          temp_m4_6_13_i;
wire signed [`CalcTempBus]          temp_m4_6_14_r;
wire signed [`CalcTempBus]          temp_m4_6_14_i;
wire signed [`CalcTempBus]          temp_m4_6_15_r;
wire signed [`CalcTempBus]          temp_m4_6_15_i;
wire signed [`CalcTempBus]          temp_m4_6_16_r;
wire signed [`CalcTempBus]          temp_m4_6_16_i;
wire signed [`CalcTempBus]          temp_m4_6_17_r;
wire signed [`CalcTempBus]          temp_m4_6_17_i;
wire signed [`CalcTempBus]          temp_m4_6_18_r;
wire signed [`CalcTempBus]          temp_m4_6_18_i;
wire signed [`CalcTempBus]          temp_m4_6_19_r;
wire signed [`CalcTempBus]          temp_m4_6_19_i;
wire signed [`CalcTempBus]          temp_m4_6_20_r;
wire signed [`CalcTempBus]          temp_m4_6_20_i;
wire signed [`CalcTempBus]          temp_m4_6_21_r;
wire signed [`CalcTempBus]          temp_m4_6_21_i;
wire signed [`CalcTempBus]          temp_m4_6_22_r;
wire signed [`CalcTempBus]          temp_m4_6_22_i;
wire signed [`CalcTempBus]          temp_m4_6_23_r;
wire signed [`CalcTempBus]          temp_m4_6_23_i;
wire signed [`CalcTempBus]          temp_m4_6_24_r;
wire signed [`CalcTempBus]          temp_m4_6_24_i;
wire signed [`CalcTempBus]          temp_m4_6_25_r;
wire signed [`CalcTempBus]          temp_m4_6_25_i;
wire signed [`CalcTempBus]          temp_m4_6_26_r;
wire signed [`CalcTempBus]          temp_m4_6_26_i;
wire signed [`CalcTempBus]          temp_m4_6_27_r;
wire signed [`CalcTempBus]          temp_m4_6_27_i;
wire signed [`CalcTempBus]          temp_m4_6_28_r;
wire signed [`CalcTempBus]          temp_m4_6_28_i;
wire signed [`CalcTempBus]          temp_m4_6_29_r;
wire signed [`CalcTempBus]          temp_m4_6_29_i;
wire signed [`CalcTempBus]          temp_m4_6_30_r;
wire signed [`CalcTempBus]          temp_m4_6_30_i;
wire signed [`CalcTempBus]          temp_m4_6_31_r;
wire signed [`CalcTempBus]          temp_m4_6_31_i;
wire signed [`CalcTempBus]          temp_m4_6_32_r;
wire signed [`CalcTempBus]          temp_m4_6_32_i;
wire signed [`CalcTempBus]          temp_m4_7_1_r;
wire signed [`CalcTempBus]          temp_m4_7_1_i;
wire signed [`CalcTempBus]          temp_m4_7_2_r;
wire signed [`CalcTempBus]          temp_m4_7_2_i;
wire signed [`CalcTempBus]          temp_m4_7_3_r;
wire signed [`CalcTempBus]          temp_m4_7_3_i;
wire signed [`CalcTempBus]          temp_m4_7_4_r;
wire signed [`CalcTempBus]          temp_m4_7_4_i;
wire signed [`CalcTempBus]          temp_m4_7_5_r;
wire signed [`CalcTempBus]          temp_m4_7_5_i;
wire signed [`CalcTempBus]          temp_m4_7_6_r;
wire signed [`CalcTempBus]          temp_m4_7_6_i;
wire signed [`CalcTempBus]          temp_m4_7_7_r;
wire signed [`CalcTempBus]          temp_m4_7_7_i;
wire signed [`CalcTempBus]          temp_m4_7_8_r;
wire signed [`CalcTempBus]          temp_m4_7_8_i;
wire signed [`CalcTempBus]          temp_m4_7_9_r;
wire signed [`CalcTempBus]          temp_m4_7_9_i;
wire signed [`CalcTempBus]          temp_m4_7_10_r;
wire signed [`CalcTempBus]          temp_m4_7_10_i;
wire signed [`CalcTempBus]          temp_m4_7_11_r;
wire signed [`CalcTempBus]          temp_m4_7_11_i;
wire signed [`CalcTempBus]          temp_m4_7_12_r;
wire signed [`CalcTempBus]          temp_m4_7_12_i;
wire signed [`CalcTempBus]          temp_m4_7_13_r;
wire signed [`CalcTempBus]          temp_m4_7_13_i;
wire signed [`CalcTempBus]          temp_m4_7_14_r;
wire signed [`CalcTempBus]          temp_m4_7_14_i;
wire signed [`CalcTempBus]          temp_m4_7_15_r;
wire signed [`CalcTempBus]          temp_m4_7_15_i;
wire signed [`CalcTempBus]          temp_m4_7_16_r;
wire signed [`CalcTempBus]          temp_m4_7_16_i;
wire signed [`CalcTempBus]          temp_m4_7_17_r;
wire signed [`CalcTempBus]          temp_m4_7_17_i;
wire signed [`CalcTempBus]          temp_m4_7_18_r;
wire signed [`CalcTempBus]          temp_m4_7_18_i;
wire signed [`CalcTempBus]          temp_m4_7_19_r;
wire signed [`CalcTempBus]          temp_m4_7_19_i;
wire signed [`CalcTempBus]          temp_m4_7_20_r;
wire signed [`CalcTempBus]          temp_m4_7_20_i;
wire signed [`CalcTempBus]          temp_m4_7_21_r;
wire signed [`CalcTempBus]          temp_m4_7_21_i;
wire signed [`CalcTempBus]          temp_m4_7_22_r;
wire signed [`CalcTempBus]          temp_m4_7_22_i;
wire signed [`CalcTempBus]          temp_m4_7_23_r;
wire signed [`CalcTempBus]          temp_m4_7_23_i;
wire signed [`CalcTempBus]          temp_m4_7_24_r;
wire signed [`CalcTempBus]          temp_m4_7_24_i;
wire signed [`CalcTempBus]          temp_m4_7_25_r;
wire signed [`CalcTempBus]          temp_m4_7_25_i;
wire signed [`CalcTempBus]          temp_m4_7_26_r;
wire signed [`CalcTempBus]          temp_m4_7_26_i;
wire signed [`CalcTempBus]          temp_m4_7_27_r;
wire signed [`CalcTempBus]          temp_m4_7_27_i;
wire signed [`CalcTempBus]          temp_m4_7_28_r;
wire signed [`CalcTempBus]          temp_m4_7_28_i;
wire signed [`CalcTempBus]          temp_m4_7_29_r;
wire signed [`CalcTempBus]          temp_m4_7_29_i;
wire signed [`CalcTempBus]          temp_m4_7_30_r;
wire signed [`CalcTempBus]          temp_m4_7_30_i;
wire signed [`CalcTempBus]          temp_m4_7_31_r;
wire signed [`CalcTempBus]          temp_m4_7_31_i;
wire signed [`CalcTempBus]          temp_m4_7_32_r;
wire signed [`CalcTempBus]          temp_m4_7_32_i;
wire signed [`CalcTempBus]          temp_m4_8_1_r;
wire signed [`CalcTempBus]          temp_m4_8_1_i;
wire signed [`CalcTempBus]          temp_m4_8_2_r;
wire signed [`CalcTempBus]          temp_m4_8_2_i;
wire signed [`CalcTempBus]          temp_m4_8_3_r;
wire signed [`CalcTempBus]          temp_m4_8_3_i;
wire signed [`CalcTempBus]          temp_m4_8_4_r;
wire signed [`CalcTempBus]          temp_m4_8_4_i;
wire signed [`CalcTempBus]          temp_m4_8_5_r;
wire signed [`CalcTempBus]          temp_m4_8_5_i;
wire signed [`CalcTempBus]          temp_m4_8_6_r;
wire signed [`CalcTempBus]          temp_m4_8_6_i;
wire signed [`CalcTempBus]          temp_m4_8_7_r;
wire signed [`CalcTempBus]          temp_m4_8_7_i;
wire signed [`CalcTempBus]          temp_m4_8_8_r;
wire signed [`CalcTempBus]          temp_m4_8_8_i;
wire signed [`CalcTempBus]          temp_m4_8_9_r;
wire signed [`CalcTempBus]          temp_m4_8_9_i;
wire signed [`CalcTempBus]          temp_m4_8_10_r;
wire signed [`CalcTempBus]          temp_m4_8_10_i;
wire signed [`CalcTempBus]          temp_m4_8_11_r;
wire signed [`CalcTempBus]          temp_m4_8_11_i;
wire signed [`CalcTempBus]          temp_m4_8_12_r;
wire signed [`CalcTempBus]          temp_m4_8_12_i;
wire signed [`CalcTempBus]          temp_m4_8_13_r;
wire signed [`CalcTempBus]          temp_m4_8_13_i;
wire signed [`CalcTempBus]          temp_m4_8_14_r;
wire signed [`CalcTempBus]          temp_m4_8_14_i;
wire signed [`CalcTempBus]          temp_m4_8_15_r;
wire signed [`CalcTempBus]          temp_m4_8_15_i;
wire signed [`CalcTempBus]          temp_m4_8_16_r;
wire signed [`CalcTempBus]          temp_m4_8_16_i;
wire signed [`CalcTempBus]          temp_m4_8_17_r;
wire signed [`CalcTempBus]          temp_m4_8_17_i;
wire signed [`CalcTempBus]          temp_m4_8_18_r;
wire signed [`CalcTempBus]          temp_m4_8_18_i;
wire signed [`CalcTempBus]          temp_m4_8_19_r;
wire signed [`CalcTempBus]          temp_m4_8_19_i;
wire signed [`CalcTempBus]          temp_m4_8_20_r;
wire signed [`CalcTempBus]          temp_m4_8_20_i;
wire signed [`CalcTempBus]          temp_m4_8_21_r;
wire signed [`CalcTempBus]          temp_m4_8_21_i;
wire signed [`CalcTempBus]          temp_m4_8_22_r;
wire signed [`CalcTempBus]          temp_m4_8_22_i;
wire signed [`CalcTempBus]          temp_m4_8_23_r;
wire signed [`CalcTempBus]          temp_m4_8_23_i;
wire signed [`CalcTempBus]          temp_m4_8_24_r;
wire signed [`CalcTempBus]          temp_m4_8_24_i;
wire signed [`CalcTempBus]          temp_m4_8_25_r;
wire signed [`CalcTempBus]          temp_m4_8_25_i;
wire signed [`CalcTempBus]          temp_m4_8_26_r;
wire signed [`CalcTempBus]          temp_m4_8_26_i;
wire signed [`CalcTempBus]          temp_m4_8_27_r;
wire signed [`CalcTempBus]          temp_m4_8_27_i;
wire signed [`CalcTempBus]          temp_m4_8_28_r;
wire signed [`CalcTempBus]          temp_m4_8_28_i;
wire signed [`CalcTempBus]          temp_m4_8_29_r;
wire signed [`CalcTempBus]          temp_m4_8_29_i;
wire signed [`CalcTempBus]          temp_m4_8_30_r;
wire signed [`CalcTempBus]          temp_m4_8_30_i;
wire signed [`CalcTempBus]          temp_m4_8_31_r;
wire signed [`CalcTempBus]          temp_m4_8_31_i;
wire signed [`CalcTempBus]          temp_m4_8_32_r;
wire signed [`CalcTempBus]          temp_m4_8_32_i;
wire signed [`CalcTempBus]          temp_m4_9_1_r;
wire signed [`CalcTempBus]          temp_m4_9_1_i;
wire signed [`CalcTempBus]          temp_m4_9_2_r;
wire signed [`CalcTempBus]          temp_m4_9_2_i;
wire signed [`CalcTempBus]          temp_m4_9_3_r;
wire signed [`CalcTempBus]          temp_m4_9_3_i;
wire signed [`CalcTempBus]          temp_m4_9_4_r;
wire signed [`CalcTempBus]          temp_m4_9_4_i;
wire signed [`CalcTempBus]          temp_m4_9_5_r;
wire signed [`CalcTempBus]          temp_m4_9_5_i;
wire signed [`CalcTempBus]          temp_m4_9_6_r;
wire signed [`CalcTempBus]          temp_m4_9_6_i;
wire signed [`CalcTempBus]          temp_m4_9_7_r;
wire signed [`CalcTempBus]          temp_m4_9_7_i;
wire signed [`CalcTempBus]          temp_m4_9_8_r;
wire signed [`CalcTempBus]          temp_m4_9_8_i;
wire signed [`CalcTempBus]          temp_m4_9_9_r;
wire signed [`CalcTempBus]          temp_m4_9_9_i;
wire signed [`CalcTempBus]          temp_m4_9_10_r;
wire signed [`CalcTempBus]          temp_m4_9_10_i;
wire signed [`CalcTempBus]          temp_m4_9_11_r;
wire signed [`CalcTempBus]          temp_m4_9_11_i;
wire signed [`CalcTempBus]          temp_m4_9_12_r;
wire signed [`CalcTempBus]          temp_m4_9_12_i;
wire signed [`CalcTempBus]          temp_m4_9_13_r;
wire signed [`CalcTempBus]          temp_m4_9_13_i;
wire signed [`CalcTempBus]          temp_m4_9_14_r;
wire signed [`CalcTempBus]          temp_m4_9_14_i;
wire signed [`CalcTempBus]          temp_m4_9_15_r;
wire signed [`CalcTempBus]          temp_m4_9_15_i;
wire signed [`CalcTempBus]          temp_m4_9_16_r;
wire signed [`CalcTempBus]          temp_m4_9_16_i;
wire signed [`CalcTempBus]          temp_m4_9_17_r;
wire signed [`CalcTempBus]          temp_m4_9_17_i;
wire signed [`CalcTempBus]          temp_m4_9_18_r;
wire signed [`CalcTempBus]          temp_m4_9_18_i;
wire signed [`CalcTempBus]          temp_m4_9_19_r;
wire signed [`CalcTempBus]          temp_m4_9_19_i;
wire signed [`CalcTempBus]          temp_m4_9_20_r;
wire signed [`CalcTempBus]          temp_m4_9_20_i;
wire signed [`CalcTempBus]          temp_m4_9_21_r;
wire signed [`CalcTempBus]          temp_m4_9_21_i;
wire signed [`CalcTempBus]          temp_m4_9_22_r;
wire signed [`CalcTempBus]          temp_m4_9_22_i;
wire signed [`CalcTempBus]          temp_m4_9_23_r;
wire signed [`CalcTempBus]          temp_m4_9_23_i;
wire signed [`CalcTempBus]          temp_m4_9_24_r;
wire signed [`CalcTempBus]          temp_m4_9_24_i;
wire signed [`CalcTempBus]          temp_m4_9_25_r;
wire signed [`CalcTempBus]          temp_m4_9_25_i;
wire signed [`CalcTempBus]          temp_m4_9_26_r;
wire signed [`CalcTempBus]          temp_m4_9_26_i;
wire signed [`CalcTempBus]          temp_m4_9_27_r;
wire signed [`CalcTempBus]          temp_m4_9_27_i;
wire signed [`CalcTempBus]          temp_m4_9_28_r;
wire signed [`CalcTempBus]          temp_m4_9_28_i;
wire signed [`CalcTempBus]          temp_m4_9_29_r;
wire signed [`CalcTempBus]          temp_m4_9_29_i;
wire signed [`CalcTempBus]          temp_m4_9_30_r;
wire signed [`CalcTempBus]          temp_m4_9_30_i;
wire signed [`CalcTempBus]          temp_m4_9_31_r;
wire signed [`CalcTempBus]          temp_m4_9_31_i;
wire signed [`CalcTempBus]          temp_m4_9_32_r;
wire signed [`CalcTempBus]          temp_m4_9_32_i;
wire signed [`CalcTempBus]          temp_m4_10_1_r;
wire signed [`CalcTempBus]          temp_m4_10_1_i;
wire signed [`CalcTempBus]          temp_m4_10_2_r;
wire signed [`CalcTempBus]          temp_m4_10_2_i;
wire signed [`CalcTempBus]          temp_m4_10_3_r;
wire signed [`CalcTempBus]          temp_m4_10_3_i;
wire signed [`CalcTempBus]          temp_m4_10_4_r;
wire signed [`CalcTempBus]          temp_m4_10_4_i;
wire signed [`CalcTempBus]          temp_m4_10_5_r;
wire signed [`CalcTempBus]          temp_m4_10_5_i;
wire signed [`CalcTempBus]          temp_m4_10_6_r;
wire signed [`CalcTempBus]          temp_m4_10_6_i;
wire signed [`CalcTempBus]          temp_m4_10_7_r;
wire signed [`CalcTempBus]          temp_m4_10_7_i;
wire signed [`CalcTempBus]          temp_m4_10_8_r;
wire signed [`CalcTempBus]          temp_m4_10_8_i;
wire signed [`CalcTempBus]          temp_m4_10_9_r;
wire signed [`CalcTempBus]          temp_m4_10_9_i;
wire signed [`CalcTempBus]          temp_m4_10_10_r;
wire signed [`CalcTempBus]          temp_m4_10_10_i;
wire signed [`CalcTempBus]          temp_m4_10_11_r;
wire signed [`CalcTempBus]          temp_m4_10_11_i;
wire signed [`CalcTempBus]          temp_m4_10_12_r;
wire signed [`CalcTempBus]          temp_m4_10_12_i;
wire signed [`CalcTempBus]          temp_m4_10_13_r;
wire signed [`CalcTempBus]          temp_m4_10_13_i;
wire signed [`CalcTempBus]          temp_m4_10_14_r;
wire signed [`CalcTempBus]          temp_m4_10_14_i;
wire signed [`CalcTempBus]          temp_m4_10_15_r;
wire signed [`CalcTempBus]          temp_m4_10_15_i;
wire signed [`CalcTempBus]          temp_m4_10_16_r;
wire signed [`CalcTempBus]          temp_m4_10_16_i;
wire signed [`CalcTempBus]          temp_m4_10_17_r;
wire signed [`CalcTempBus]          temp_m4_10_17_i;
wire signed [`CalcTempBus]          temp_m4_10_18_r;
wire signed [`CalcTempBus]          temp_m4_10_18_i;
wire signed [`CalcTempBus]          temp_m4_10_19_r;
wire signed [`CalcTempBus]          temp_m4_10_19_i;
wire signed [`CalcTempBus]          temp_m4_10_20_r;
wire signed [`CalcTempBus]          temp_m4_10_20_i;
wire signed [`CalcTempBus]          temp_m4_10_21_r;
wire signed [`CalcTempBus]          temp_m4_10_21_i;
wire signed [`CalcTempBus]          temp_m4_10_22_r;
wire signed [`CalcTempBus]          temp_m4_10_22_i;
wire signed [`CalcTempBus]          temp_m4_10_23_r;
wire signed [`CalcTempBus]          temp_m4_10_23_i;
wire signed [`CalcTempBus]          temp_m4_10_24_r;
wire signed [`CalcTempBus]          temp_m4_10_24_i;
wire signed [`CalcTempBus]          temp_m4_10_25_r;
wire signed [`CalcTempBus]          temp_m4_10_25_i;
wire signed [`CalcTempBus]          temp_m4_10_26_r;
wire signed [`CalcTempBus]          temp_m4_10_26_i;
wire signed [`CalcTempBus]          temp_m4_10_27_r;
wire signed [`CalcTempBus]          temp_m4_10_27_i;
wire signed [`CalcTempBus]          temp_m4_10_28_r;
wire signed [`CalcTempBus]          temp_m4_10_28_i;
wire signed [`CalcTempBus]          temp_m4_10_29_r;
wire signed [`CalcTempBus]          temp_m4_10_29_i;
wire signed [`CalcTempBus]          temp_m4_10_30_r;
wire signed [`CalcTempBus]          temp_m4_10_30_i;
wire signed [`CalcTempBus]          temp_m4_10_31_r;
wire signed [`CalcTempBus]          temp_m4_10_31_i;
wire signed [`CalcTempBus]          temp_m4_10_32_r;
wire signed [`CalcTempBus]          temp_m4_10_32_i;
wire signed [`CalcTempBus]          temp_m4_11_1_r;
wire signed [`CalcTempBus]          temp_m4_11_1_i;
wire signed [`CalcTempBus]          temp_m4_11_2_r;
wire signed [`CalcTempBus]          temp_m4_11_2_i;
wire signed [`CalcTempBus]          temp_m4_11_3_r;
wire signed [`CalcTempBus]          temp_m4_11_3_i;
wire signed [`CalcTempBus]          temp_m4_11_4_r;
wire signed [`CalcTempBus]          temp_m4_11_4_i;
wire signed [`CalcTempBus]          temp_m4_11_5_r;
wire signed [`CalcTempBus]          temp_m4_11_5_i;
wire signed [`CalcTempBus]          temp_m4_11_6_r;
wire signed [`CalcTempBus]          temp_m4_11_6_i;
wire signed [`CalcTempBus]          temp_m4_11_7_r;
wire signed [`CalcTempBus]          temp_m4_11_7_i;
wire signed [`CalcTempBus]          temp_m4_11_8_r;
wire signed [`CalcTempBus]          temp_m4_11_8_i;
wire signed [`CalcTempBus]          temp_m4_11_9_r;
wire signed [`CalcTempBus]          temp_m4_11_9_i;
wire signed [`CalcTempBus]          temp_m4_11_10_r;
wire signed [`CalcTempBus]          temp_m4_11_10_i;
wire signed [`CalcTempBus]          temp_m4_11_11_r;
wire signed [`CalcTempBus]          temp_m4_11_11_i;
wire signed [`CalcTempBus]          temp_m4_11_12_r;
wire signed [`CalcTempBus]          temp_m4_11_12_i;
wire signed [`CalcTempBus]          temp_m4_11_13_r;
wire signed [`CalcTempBus]          temp_m4_11_13_i;
wire signed [`CalcTempBus]          temp_m4_11_14_r;
wire signed [`CalcTempBus]          temp_m4_11_14_i;
wire signed [`CalcTempBus]          temp_m4_11_15_r;
wire signed [`CalcTempBus]          temp_m4_11_15_i;
wire signed [`CalcTempBus]          temp_m4_11_16_r;
wire signed [`CalcTempBus]          temp_m4_11_16_i;
wire signed [`CalcTempBus]          temp_m4_11_17_r;
wire signed [`CalcTempBus]          temp_m4_11_17_i;
wire signed [`CalcTempBus]          temp_m4_11_18_r;
wire signed [`CalcTempBus]          temp_m4_11_18_i;
wire signed [`CalcTempBus]          temp_m4_11_19_r;
wire signed [`CalcTempBus]          temp_m4_11_19_i;
wire signed [`CalcTempBus]          temp_m4_11_20_r;
wire signed [`CalcTempBus]          temp_m4_11_20_i;
wire signed [`CalcTempBus]          temp_m4_11_21_r;
wire signed [`CalcTempBus]          temp_m4_11_21_i;
wire signed [`CalcTempBus]          temp_m4_11_22_r;
wire signed [`CalcTempBus]          temp_m4_11_22_i;
wire signed [`CalcTempBus]          temp_m4_11_23_r;
wire signed [`CalcTempBus]          temp_m4_11_23_i;
wire signed [`CalcTempBus]          temp_m4_11_24_r;
wire signed [`CalcTempBus]          temp_m4_11_24_i;
wire signed [`CalcTempBus]          temp_m4_11_25_r;
wire signed [`CalcTempBus]          temp_m4_11_25_i;
wire signed [`CalcTempBus]          temp_m4_11_26_r;
wire signed [`CalcTempBus]          temp_m4_11_26_i;
wire signed [`CalcTempBus]          temp_m4_11_27_r;
wire signed [`CalcTempBus]          temp_m4_11_27_i;
wire signed [`CalcTempBus]          temp_m4_11_28_r;
wire signed [`CalcTempBus]          temp_m4_11_28_i;
wire signed [`CalcTempBus]          temp_m4_11_29_r;
wire signed [`CalcTempBus]          temp_m4_11_29_i;
wire signed [`CalcTempBus]          temp_m4_11_30_r;
wire signed [`CalcTempBus]          temp_m4_11_30_i;
wire signed [`CalcTempBus]          temp_m4_11_31_r;
wire signed [`CalcTempBus]          temp_m4_11_31_i;
wire signed [`CalcTempBus]          temp_m4_11_32_r;
wire signed [`CalcTempBus]          temp_m4_11_32_i;
wire signed [`CalcTempBus]          temp_m4_12_1_r;
wire signed [`CalcTempBus]          temp_m4_12_1_i;
wire signed [`CalcTempBus]          temp_m4_12_2_r;
wire signed [`CalcTempBus]          temp_m4_12_2_i;
wire signed [`CalcTempBus]          temp_m4_12_3_r;
wire signed [`CalcTempBus]          temp_m4_12_3_i;
wire signed [`CalcTempBus]          temp_m4_12_4_r;
wire signed [`CalcTempBus]          temp_m4_12_4_i;
wire signed [`CalcTempBus]          temp_m4_12_5_r;
wire signed [`CalcTempBus]          temp_m4_12_5_i;
wire signed [`CalcTempBus]          temp_m4_12_6_r;
wire signed [`CalcTempBus]          temp_m4_12_6_i;
wire signed [`CalcTempBus]          temp_m4_12_7_r;
wire signed [`CalcTempBus]          temp_m4_12_7_i;
wire signed [`CalcTempBus]          temp_m4_12_8_r;
wire signed [`CalcTempBus]          temp_m4_12_8_i;
wire signed [`CalcTempBus]          temp_m4_12_9_r;
wire signed [`CalcTempBus]          temp_m4_12_9_i;
wire signed [`CalcTempBus]          temp_m4_12_10_r;
wire signed [`CalcTempBus]          temp_m4_12_10_i;
wire signed [`CalcTempBus]          temp_m4_12_11_r;
wire signed [`CalcTempBus]          temp_m4_12_11_i;
wire signed [`CalcTempBus]          temp_m4_12_12_r;
wire signed [`CalcTempBus]          temp_m4_12_12_i;
wire signed [`CalcTempBus]          temp_m4_12_13_r;
wire signed [`CalcTempBus]          temp_m4_12_13_i;
wire signed [`CalcTempBus]          temp_m4_12_14_r;
wire signed [`CalcTempBus]          temp_m4_12_14_i;
wire signed [`CalcTempBus]          temp_m4_12_15_r;
wire signed [`CalcTempBus]          temp_m4_12_15_i;
wire signed [`CalcTempBus]          temp_m4_12_16_r;
wire signed [`CalcTempBus]          temp_m4_12_16_i;
wire signed [`CalcTempBus]          temp_m4_12_17_r;
wire signed [`CalcTempBus]          temp_m4_12_17_i;
wire signed [`CalcTempBus]          temp_m4_12_18_r;
wire signed [`CalcTempBus]          temp_m4_12_18_i;
wire signed [`CalcTempBus]          temp_m4_12_19_r;
wire signed [`CalcTempBus]          temp_m4_12_19_i;
wire signed [`CalcTempBus]          temp_m4_12_20_r;
wire signed [`CalcTempBus]          temp_m4_12_20_i;
wire signed [`CalcTempBus]          temp_m4_12_21_r;
wire signed [`CalcTempBus]          temp_m4_12_21_i;
wire signed [`CalcTempBus]          temp_m4_12_22_r;
wire signed [`CalcTempBus]          temp_m4_12_22_i;
wire signed [`CalcTempBus]          temp_m4_12_23_r;
wire signed [`CalcTempBus]          temp_m4_12_23_i;
wire signed [`CalcTempBus]          temp_m4_12_24_r;
wire signed [`CalcTempBus]          temp_m4_12_24_i;
wire signed [`CalcTempBus]          temp_m4_12_25_r;
wire signed [`CalcTempBus]          temp_m4_12_25_i;
wire signed [`CalcTempBus]          temp_m4_12_26_r;
wire signed [`CalcTempBus]          temp_m4_12_26_i;
wire signed [`CalcTempBus]          temp_m4_12_27_r;
wire signed [`CalcTempBus]          temp_m4_12_27_i;
wire signed [`CalcTempBus]          temp_m4_12_28_r;
wire signed [`CalcTempBus]          temp_m4_12_28_i;
wire signed [`CalcTempBus]          temp_m4_12_29_r;
wire signed [`CalcTempBus]          temp_m4_12_29_i;
wire signed [`CalcTempBus]          temp_m4_12_30_r;
wire signed [`CalcTempBus]          temp_m4_12_30_i;
wire signed [`CalcTempBus]          temp_m4_12_31_r;
wire signed [`CalcTempBus]          temp_m4_12_31_i;
wire signed [`CalcTempBus]          temp_m4_12_32_r;
wire signed [`CalcTempBus]          temp_m4_12_32_i;
wire signed [`CalcTempBus]          temp_m4_13_1_r;
wire signed [`CalcTempBus]          temp_m4_13_1_i;
wire signed [`CalcTempBus]          temp_m4_13_2_r;
wire signed [`CalcTempBus]          temp_m4_13_2_i;
wire signed [`CalcTempBus]          temp_m4_13_3_r;
wire signed [`CalcTempBus]          temp_m4_13_3_i;
wire signed [`CalcTempBus]          temp_m4_13_4_r;
wire signed [`CalcTempBus]          temp_m4_13_4_i;
wire signed [`CalcTempBus]          temp_m4_13_5_r;
wire signed [`CalcTempBus]          temp_m4_13_5_i;
wire signed [`CalcTempBus]          temp_m4_13_6_r;
wire signed [`CalcTempBus]          temp_m4_13_6_i;
wire signed [`CalcTempBus]          temp_m4_13_7_r;
wire signed [`CalcTempBus]          temp_m4_13_7_i;
wire signed [`CalcTempBus]          temp_m4_13_8_r;
wire signed [`CalcTempBus]          temp_m4_13_8_i;
wire signed [`CalcTempBus]          temp_m4_13_9_r;
wire signed [`CalcTempBus]          temp_m4_13_9_i;
wire signed [`CalcTempBus]          temp_m4_13_10_r;
wire signed [`CalcTempBus]          temp_m4_13_10_i;
wire signed [`CalcTempBus]          temp_m4_13_11_r;
wire signed [`CalcTempBus]          temp_m4_13_11_i;
wire signed [`CalcTempBus]          temp_m4_13_12_r;
wire signed [`CalcTempBus]          temp_m4_13_12_i;
wire signed [`CalcTempBus]          temp_m4_13_13_r;
wire signed [`CalcTempBus]          temp_m4_13_13_i;
wire signed [`CalcTempBus]          temp_m4_13_14_r;
wire signed [`CalcTempBus]          temp_m4_13_14_i;
wire signed [`CalcTempBus]          temp_m4_13_15_r;
wire signed [`CalcTempBus]          temp_m4_13_15_i;
wire signed [`CalcTempBus]          temp_m4_13_16_r;
wire signed [`CalcTempBus]          temp_m4_13_16_i;
wire signed [`CalcTempBus]          temp_m4_13_17_r;
wire signed [`CalcTempBus]          temp_m4_13_17_i;
wire signed [`CalcTempBus]          temp_m4_13_18_r;
wire signed [`CalcTempBus]          temp_m4_13_18_i;
wire signed [`CalcTempBus]          temp_m4_13_19_r;
wire signed [`CalcTempBus]          temp_m4_13_19_i;
wire signed [`CalcTempBus]          temp_m4_13_20_r;
wire signed [`CalcTempBus]          temp_m4_13_20_i;
wire signed [`CalcTempBus]          temp_m4_13_21_r;
wire signed [`CalcTempBus]          temp_m4_13_21_i;
wire signed [`CalcTempBus]          temp_m4_13_22_r;
wire signed [`CalcTempBus]          temp_m4_13_22_i;
wire signed [`CalcTempBus]          temp_m4_13_23_r;
wire signed [`CalcTempBus]          temp_m4_13_23_i;
wire signed [`CalcTempBus]          temp_m4_13_24_r;
wire signed [`CalcTempBus]          temp_m4_13_24_i;
wire signed [`CalcTempBus]          temp_m4_13_25_r;
wire signed [`CalcTempBus]          temp_m4_13_25_i;
wire signed [`CalcTempBus]          temp_m4_13_26_r;
wire signed [`CalcTempBus]          temp_m4_13_26_i;
wire signed [`CalcTempBus]          temp_m4_13_27_r;
wire signed [`CalcTempBus]          temp_m4_13_27_i;
wire signed [`CalcTempBus]          temp_m4_13_28_r;
wire signed [`CalcTempBus]          temp_m4_13_28_i;
wire signed [`CalcTempBus]          temp_m4_13_29_r;
wire signed [`CalcTempBus]          temp_m4_13_29_i;
wire signed [`CalcTempBus]          temp_m4_13_30_r;
wire signed [`CalcTempBus]          temp_m4_13_30_i;
wire signed [`CalcTempBus]          temp_m4_13_31_r;
wire signed [`CalcTempBus]          temp_m4_13_31_i;
wire signed [`CalcTempBus]          temp_m4_13_32_r;
wire signed [`CalcTempBus]          temp_m4_13_32_i;
wire signed [`CalcTempBus]          temp_m4_14_1_r;
wire signed [`CalcTempBus]          temp_m4_14_1_i;
wire signed [`CalcTempBus]          temp_m4_14_2_r;
wire signed [`CalcTempBus]          temp_m4_14_2_i;
wire signed [`CalcTempBus]          temp_m4_14_3_r;
wire signed [`CalcTempBus]          temp_m4_14_3_i;
wire signed [`CalcTempBus]          temp_m4_14_4_r;
wire signed [`CalcTempBus]          temp_m4_14_4_i;
wire signed [`CalcTempBus]          temp_m4_14_5_r;
wire signed [`CalcTempBus]          temp_m4_14_5_i;
wire signed [`CalcTempBus]          temp_m4_14_6_r;
wire signed [`CalcTempBus]          temp_m4_14_6_i;
wire signed [`CalcTempBus]          temp_m4_14_7_r;
wire signed [`CalcTempBus]          temp_m4_14_7_i;
wire signed [`CalcTempBus]          temp_m4_14_8_r;
wire signed [`CalcTempBus]          temp_m4_14_8_i;
wire signed [`CalcTempBus]          temp_m4_14_9_r;
wire signed [`CalcTempBus]          temp_m4_14_9_i;
wire signed [`CalcTempBus]          temp_m4_14_10_r;
wire signed [`CalcTempBus]          temp_m4_14_10_i;
wire signed [`CalcTempBus]          temp_m4_14_11_r;
wire signed [`CalcTempBus]          temp_m4_14_11_i;
wire signed [`CalcTempBus]          temp_m4_14_12_r;
wire signed [`CalcTempBus]          temp_m4_14_12_i;
wire signed [`CalcTempBus]          temp_m4_14_13_r;
wire signed [`CalcTempBus]          temp_m4_14_13_i;
wire signed [`CalcTempBus]          temp_m4_14_14_r;
wire signed [`CalcTempBus]          temp_m4_14_14_i;
wire signed [`CalcTempBus]          temp_m4_14_15_r;
wire signed [`CalcTempBus]          temp_m4_14_15_i;
wire signed [`CalcTempBus]          temp_m4_14_16_r;
wire signed [`CalcTempBus]          temp_m4_14_16_i;
wire signed [`CalcTempBus]          temp_m4_14_17_r;
wire signed [`CalcTempBus]          temp_m4_14_17_i;
wire signed [`CalcTempBus]          temp_m4_14_18_r;
wire signed [`CalcTempBus]          temp_m4_14_18_i;
wire signed [`CalcTempBus]          temp_m4_14_19_r;
wire signed [`CalcTempBus]          temp_m4_14_19_i;
wire signed [`CalcTempBus]          temp_m4_14_20_r;
wire signed [`CalcTempBus]          temp_m4_14_20_i;
wire signed [`CalcTempBus]          temp_m4_14_21_r;
wire signed [`CalcTempBus]          temp_m4_14_21_i;
wire signed [`CalcTempBus]          temp_m4_14_22_r;
wire signed [`CalcTempBus]          temp_m4_14_22_i;
wire signed [`CalcTempBus]          temp_m4_14_23_r;
wire signed [`CalcTempBus]          temp_m4_14_23_i;
wire signed [`CalcTempBus]          temp_m4_14_24_r;
wire signed [`CalcTempBus]          temp_m4_14_24_i;
wire signed [`CalcTempBus]          temp_m4_14_25_r;
wire signed [`CalcTempBus]          temp_m4_14_25_i;
wire signed [`CalcTempBus]          temp_m4_14_26_r;
wire signed [`CalcTempBus]          temp_m4_14_26_i;
wire signed [`CalcTempBus]          temp_m4_14_27_r;
wire signed [`CalcTempBus]          temp_m4_14_27_i;
wire signed [`CalcTempBus]          temp_m4_14_28_r;
wire signed [`CalcTempBus]          temp_m4_14_28_i;
wire signed [`CalcTempBus]          temp_m4_14_29_r;
wire signed [`CalcTempBus]          temp_m4_14_29_i;
wire signed [`CalcTempBus]          temp_m4_14_30_r;
wire signed [`CalcTempBus]          temp_m4_14_30_i;
wire signed [`CalcTempBus]          temp_m4_14_31_r;
wire signed [`CalcTempBus]          temp_m4_14_31_i;
wire signed [`CalcTempBus]          temp_m4_14_32_r;
wire signed [`CalcTempBus]          temp_m4_14_32_i;
wire signed [`CalcTempBus]          temp_m4_15_1_r;
wire signed [`CalcTempBus]          temp_m4_15_1_i;
wire signed [`CalcTempBus]          temp_m4_15_2_r;
wire signed [`CalcTempBus]          temp_m4_15_2_i;
wire signed [`CalcTempBus]          temp_m4_15_3_r;
wire signed [`CalcTempBus]          temp_m4_15_3_i;
wire signed [`CalcTempBus]          temp_m4_15_4_r;
wire signed [`CalcTempBus]          temp_m4_15_4_i;
wire signed [`CalcTempBus]          temp_m4_15_5_r;
wire signed [`CalcTempBus]          temp_m4_15_5_i;
wire signed [`CalcTempBus]          temp_m4_15_6_r;
wire signed [`CalcTempBus]          temp_m4_15_6_i;
wire signed [`CalcTempBus]          temp_m4_15_7_r;
wire signed [`CalcTempBus]          temp_m4_15_7_i;
wire signed [`CalcTempBus]          temp_m4_15_8_r;
wire signed [`CalcTempBus]          temp_m4_15_8_i;
wire signed [`CalcTempBus]          temp_m4_15_9_r;
wire signed [`CalcTempBus]          temp_m4_15_9_i;
wire signed [`CalcTempBus]          temp_m4_15_10_r;
wire signed [`CalcTempBus]          temp_m4_15_10_i;
wire signed [`CalcTempBus]          temp_m4_15_11_r;
wire signed [`CalcTempBus]          temp_m4_15_11_i;
wire signed [`CalcTempBus]          temp_m4_15_12_r;
wire signed [`CalcTempBus]          temp_m4_15_12_i;
wire signed [`CalcTempBus]          temp_m4_15_13_r;
wire signed [`CalcTempBus]          temp_m4_15_13_i;
wire signed [`CalcTempBus]          temp_m4_15_14_r;
wire signed [`CalcTempBus]          temp_m4_15_14_i;
wire signed [`CalcTempBus]          temp_m4_15_15_r;
wire signed [`CalcTempBus]          temp_m4_15_15_i;
wire signed [`CalcTempBus]          temp_m4_15_16_r;
wire signed [`CalcTempBus]          temp_m4_15_16_i;
wire signed [`CalcTempBus]          temp_m4_15_17_r;
wire signed [`CalcTempBus]          temp_m4_15_17_i;
wire signed [`CalcTempBus]          temp_m4_15_18_r;
wire signed [`CalcTempBus]          temp_m4_15_18_i;
wire signed [`CalcTempBus]          temp_m4_15_19_r;
wire signed [`CalcTempBus]          temp_m4_15_19_i;
wire signed [`CalcTempBus]          temp_m4_15_20_r;
wire signed [`CalcTempBus]          temp_m4_15_20_i;
wire signed [`CalcTempBus]          temp_m4_15_21_r;
wire signed [`CalcTempBus]          temp_m4_15_21_i;
wire signed [`CalcTempBus]          temp_m4_15_22_r;
wire signed [`CalcTempBus]          temp_m4_15_22_i;
wire signed [`CalcTempBus]          temp_m4_15_23_r;
wire signed [`CalcTempBus]          temp_m4_15_23_i;
wire signed [`CalcTempBus]          temp_m4_15_24_r;
wire signed [`CalcTempBus]          temp_m4_15_24_i;
wire signed [`CalcTempBus]          temp_m4_15_25_r;
wire signed [`CalcTempBus]          temp_m4_15_25_i;
wire signed [`CalcTempBus]          temp_m4_15_26_r;
wire signed [`CalcTempBus]          temp_m4_15_26_i;
wire signed [`CalcTempBus]          temp_m4_15_27_r;
wire signed [`CalcTempBus]          temp_m4_15_27_i;
wire signed [`CalcTempBus]          temp_m4_15_28_r;
wire signed [`CalcTempBus]          temp_m4_15_28_i;
wire signed [`CalcTempBus]          temp_m4_15_29_r;
wire signed [`CalcTempBus]          temp_m4_15_29_i;
wire signed [`CalcTempBus]          temp_m4_15_30_r;
wire signed [`CalcTempBus]          temp_m4_15_30_i;
wire signed [`CalcTempBus]          temp_m4_15_31_r;
wire signed [`CalcTempBus]          temp_m4_15_31_i;
wire signed [`CalcTempBus]          temp_m4_15_32_r;
wire signed [`CalcTempBus]          temp_m4_15_32_i;
wire signed [`CalcTempBus]          temp_m4_16_1_r;
wire signed [`CalcTempBus]          temp_m4_16_1_i;
wire signed [`CalcTempBus]          temp_m4_16_2_r;
wire signed [`CalcTempBus]          temp_m4_16_2_i;
wire signed [`CalcTempBus]          temp_m4_16_3_r;
wire signed [`CalcTempBus]          temp_m4_16_3_i;
wire signed [`CalcTempBus]          temp_m4_16_4_r;
wire signed [`CalcTempBus]          temp_m4_16_4_i;
wire signed [`CalcTempBus]          temp_m4_16_5_r;
wire signed [`CalcTempBus]          temp_m4_16_5_i;
wire signed [`CalcTempBus]          temp_m4_16_6_r;
wire signed [`CalcTempBus]          temp_m4_16_6_i;
wire signed [`CalcTempBus]          temp_m4_16_7_r;
wire signed [`CalcTempBus]          temp_m4_16_7_i;
wire signed [`CalcTempBus]          temp_m4_16_8_r;
wire signed [`CalcTempBus]          temp_m4_16_8_i;
wire signed [`CalcTempBus]          temp_m4_16_9_r;
wire signed [`CalcTempBus]          temp_m4_16_9_i;
wire signed [`CalcTempBus]          temp_m4_16_10_r;
wire signed [`CalcTempBus]          temp_m4_16_10_i;
wire signed [`CalcTempBus]          temp_m4_16_11_r;
wire signed [`CalcTempBus]          temp_m4_16_11_i;
wire signed [`CalcTempBus]          temp_m4_16_12_r;
wire signed [`CalcTempBus]          temp_m4_16_12_i;
wire signed [`CalcTempBus]          temp_m4_16_13_r;
wire signed [`CalcTempBus]          temp_m4_16_13_i;
wire signed [`CalcTempBus]          temp_m4_16_14_r;
wire signed [`CalcTempBus]          temp_m4_16_14_i;
wire signed [`CalcTempBus]          temp_m4_16_15_r;
wire signed [`CalcTempBus]          temp_m4_16_15_i;
wire signed [`CalcTempBus]          temp_m4_16_16_r;
wire signed [`CalcTempBus]          temp_m4_16_16_i;
wire signed [`CalcTempBus]          temp_m4_16_17_r;
wire signed [`CalcTempBus]          temp_m4_16_17_i;
wire signed [`CalcTempBus]          temp_m4_16_18_r;
wire signed [`CalcTempBus]          temp_m4_16_18_i;
wire signed [`CalcTempBus]          temp_m4_16_19_r;
wire signed [`CalcTempBus]          temp_m4_16_19_i;
wire signed [`CalcTempBus]          temp_m4_16_20_r;
wire signed [`CalcTempBus]          temp_m4_16_20_i;
wire signed [`CalcTempBus]          temp_m4_16_21_r;
wire signed [`CalcTempBus]          temp_m4_16_21_i;
wire signed [`CalcTempBus]          temp_m4_16_22_r;
wire signed [`CalcTempBus]          temp_m4_16_22_i;
wire signed [`CalcTempBus]          temp_m4_16_23_r;
wire signed [`CalcTempBus]          temp_m4_16_23_i;
wire signed [`CalcTempBus]          temp_m4_16_24_r;
wire signed [`CalcTempBus]          temp_m4_16_24_i;
wire signed [`CalcTempBus]          temp_m4_16_25_r;
wire signed [`CalcTempBus]          temp_m4_16_25_i;
wire signed [`CalcTempBus]          temp_m4_16_26_r;
wire signed [`CalcTempBus]          temp_m4_16_26_i;
wire signed [`CalcTempBus]          temp_m4_16_27_r;
wire signed [`CalcTempBus]          temp_m4_16_27_i;
wire signed [`CalcTempBus]          temp_m4_16_28_r;
wire signed [`CalcTempBus]          temp_m4_16_28_i;
wire signed [`CalcTempBus]          temp_m4_16_29_r;
wire signed [`CalcTempBus]          temp_m4_16_29_i;
wire signed [`CalcTempBus]          temp_m4_16_30_r;
wire signed [`CalcTempBus]          temp_m4_16_30_i;
wire signed [`CalcTempBus]          temp_m4_16_31_r;
wire signed [`CalcTempBus]          temp_m4_16_31_i;
wire signed [`CalcTempBus]          temp_m4_16_32_r;
wire signed [`CalcTempBus]          temp_m4_16_32_i;
wire signed [`CalcTempBus]          temp_m4_17_1_r;
wire signed [`CalcTempBus]          temp_m4_17_1_i;
wire signed [`CalcTempBus]          temp_m4_17_2_r;
wire signed [`CalcTempBus]          temp_m4_17_2_i;
wire signed [`CalcTempBus]          temp_m4_17_3_r;
wire signed [`CalcTempBus]          temp_m4_17_3_i;
wire signed [`CalcTempBus]          temp_m4_17_4_r;
wire signed [`CalcTempBus]          temp_m4_17_4_i;
wire signed [`CalcTempBus]          temp_m4_17_5_r;
wire signed [`CalcTempBus]          temp_m4_17_5_i;
wire signed [`CalcTempBus]          temp_m4_17_6_r;
wire signed [`CalcTempBus]          temp_m4_17_6_i;
wire signed [`CalcTempBus]          temp_m4_17_7_r;
wire signed [`CalcTempBus]          temp_m4_17_7_i;
wire signed [`CalcTempBus]          temp_m4_17_8_r;
wire signed [`CalcTempBus]          temp_m4_17_8_i;
wire signed [`CalcTempBus]          temp_m4_17_9_r;
wire signed [`CalcTempBus]          temp_m4_17_9_i;
wire signed [`CalcTempBus]          temp_m4_17_10_r;
wire signed [`CalcTempBus]          temp_m4_17_10_i;
wire signed [`CalcTempBus]          temp_m4_17_11_r;
wire signed [`CalcTempBus]          temp_m4_17_11_i;
wire signed [`CalcTempBus]          temp_m4_17_12_r;
wire signed [`CalcTempBus]          temp_m4_17_12_i;
wire signed [`CalcTempBus]          temp_m4_17_13_r;
wire signed [`CalcTempBus]          temp_m4_17_13_i;
wire signed [`CalcTempBus]          temp_m4_17_14_r;
wire signed [`CalcTempBus]          temp_m4_17_14_i;
wire signed [`CalcTempBus]          temp_m4_17_15_r;
wire signed [`CalcTempBus]          temp_m4_17_15_i;
wire signed [`CalcTempBus]          temp_m4_17_16_r;
wire signed [`CalcTempBus]          temp_m4_17_16_i;
wire signed [`CalcTempBus]          temp_m4_17_17_r;
wire signed [`CalcTempBus]          temp_m4_17_17_i;
wire signed [`CalcTempBus]          temp_m4_17_18_r;
wire signed [`CalcTempBus]          temp_m4_17_18_i;
wire signed [`CalcTempBus]          temp_m4_17_19_r;
wire signed [`CalcTempBus]          temp_m4_17_19_i;
wire signed [`CalcTempBus]          temp_m4_17_20_r;
wire signed [`CalcTempBus]          temp_m4_17_20_i;
wire signed [`CalcTempBus]          temp_m4_17_21_r;
wire signed [`CalcTempBus]          temp_m4_17_21_i;
wire signed [`CalcTempBus]          temp_m4_17_22_r;
wire signed [`CalcTempBus]          temp_m4_17_22_i;
wire signed [`CalcTempBus]          temp_m4_17_23_r;
wire signed [`CalcTempBus]          temp_m4_17_23_i;
wire signed [`CalcTempBus]          temp_m4_17_24_r;
wire signed [`CalcTempBus]          temp_m4_17_24_i;
wire signed [`CalcTempBus]          temp_m4_17_25_r;
wire signed [`CalcTempBus]          temp_m4_17_25_i;
wire signed [`CalcTempBus]          temp_m4_17_26_r;
wire signed [`CalcTempBus]          temp_m4_17_26_i;
wire signed [`CalcTempBus]          temp_m4_17_27_r;
wire signed [`CalcTempBus]          temp_m4_17_27_i;
wire signed [`CalcTempBus]          temp_m4_17_28_r;
wire signed [`CalcTempBus]          temp_m4_17_28_i;
wire signed [`CalcTempBus]          temp_m4_17_29_r;
wire signed [`CalcTempBus]          temp_m4_17_29_i;
wire signed [`CalcTempBus]          temp_m4_17_30_r;
wire signed [`CalcTempBus]          temp_m4_17_30_i;
wire signed [`CalcTempBus]          temp_m4_17_31_r;
wire signed [`CalcTempBus]          temp_m4_17_31_i;
wire signed [`CalcTempBus]          temp_m4_17_32_r;
wire signed [`CalcTempBus]          temp_m4_17_32_i;
wire signed [`CalcTempBus]          temp_m4_18_1_r;
wire signed [`CalcTempBus]          temp_m4_18_1_i;
wire signed [`CalcTempBus]          temp_m4_18_2_r;
wire signed [`CalcTempBus]          temp_m4_18_2_i;
wire signed [`CalcTempBus]          temp_m4_18_3_r;
wire signed [`CalcTempBus]          temp_m4_18_3_i;
wire signed [`CalcTempBus]          temp_m4_18_4_r;
wire signed [`CalcTempBus]          temp_m4_18_4_i;
wire signed [`CalcTempBus]          temp_m4_18_5_r;
wire signed [`CalcTempBus]          temp_m4_18_5_i;
wire signed [`CalcTempBus]          temp_m4_18_6_r;
wire signed [`CalcTempBus]          temp_m4_18_6_i;
wire signed [`CalcTempBus]          temp_m4_18_7_r;
wire signed [`CalcTempBus]          temp_m4_18_7_i;
wire signed [`CalcTempBus]          temp_m4_18_8_r;
wire signed [`CalcTempBus]          temp_m4_18_8_i;
wire signed [`CalcTempBus]          temp_m4_18_9_r;
wire signed [`CalcTempBus]          temp_m4_18_9_i;
wire signed [`CalcTempBus]          temp_m4_18_10_r;
wire signed [`CalcTempBus]          temp_m4_18_10_i;
wire signed [`CalcTempBus]          temp_m4_18_11_r;
wire signed [`CalcTempBus]          temp_m4_18_11_i;
wire signed [`CalcTempBus]          temp_m4_18_12_r;
wire signed [`CalcTempBus]          temp_m4_18_12_i;
wire signed [`CalcTempBus]          temp_m4_18_13_r;
wire signed [`CalcTempBus]          temp_m4_18_13_i;
wire signed [`CalcTempBus]          temp_m4_18_14_r;
wire signed [`CalcTempBus]          temp_m4_18_14_i;
wire signed [`CalcTempBus]          temp_m4_18_15_r;
wire signed [`CalcTempBus]          temp_m4_18_15_i;
wire signed [`CalcTempBus]          temp_m4_18_16_r;
wire signed [`CalcTempBus]          temp_m4_18_16_i;
wire signed [`CalcTempBus]          temp_m4_18_17_r;
wire signed [`CalcTempBus]          temp_m4_18_17_i;
wire signed [`CalcTempBus]          temp_m4_18_18_r;
wire signed [`CalcTempBus]          temp_m4_18_18_i;
wire signed [`CalcTempBus]          temp_m4_18_19_r;
wire signed [`CalcTempBus]          temp_m4_18_19_i;
wire signed [`CalcTempBus]          temp_m4_18_20_r;
wire signed [`CalcTempBus]          temp_m4_18_20_i;
wire signed [`CalcTempBus]          temp_m4_18_21_r;
wire signed [`CalcTempBus]          temp_m4_18_21_i;
wire signed [`CalcTempBus]          temp_m4_18_22_r;
wire signed [`CalcTempBus]          temp_m4_18_22_i;
wire signed [`CalcTempBus]          temp_m4_18_23_r;
wire signed [`CalcTempBus]          temp_m4_18_23_i;
wire signed [`CalcTempBus]          temp_m4_18_24_r;
wire signed [`CalcTempBus]          temp_m4_18_24_i;
wire signed [`CalcTempBus]          temp_m4_18_25_r;
wire signed [`CalcTempBus]          temp_m4_18_25_i;
wire signed [`CalcTempBus]          temp_m4_18_26_r;
wire signed [`CalcTempBus]          temp_m4_18_26_i;
wire signed [`CalcTempBus]          temp_m4_18_27_r;
wire signed [`CalcTempBus]          temp_m4_18_27_i;
wire signed [`CalcTempBus]          temp_m4_18_28_r;
wire signed [`CalcTempBus]          temp_m4_18_28_i;
wire signed [`CalcTempBus]          temp_m4_18_29_r;
wire signed [`CalcTempBus]          temp_m4_18_29_i;
wire signed [`CalcTempBus]          temp_m4_18_30_r;
wire signed [`CalcTempBus]          temp_m4_18_30_i;
wire signed [`CalcTempBus]          temp_m4_18_31_r;
wire signed [`CalcTempBus]          temp_m4_18_31_i;
wire signed [`CalcTempBus]          temp_m4_18_32_r;
wire signed [`CalcTempBus]          temp_m4_18_32_i;
wire signed [`CalcTempBus]          temp_m4_19_1_r;
wire signed [`CalcTempBus]          temp_m4_19_1_i;
wire signed [`CalcTempBus]          temp_m4_19_2_r;
wire signed [`CalcTempBus]          temp_m4_19_2_i;
wire signed [`CalcTempBus]          temp_m4_19_3_r;
wire signed [`CalcTempBus]          temp_m4_19_3_i;
wire signed [`CalcTempBus]          temp_m4_19_4_r;
wire signed [`CalcTempBus]          temp_m4_19_4_i;
wire signed [`CalcTempBus]          temp_m4_19_5_r;
wire signed [`CalcTempBus]          temp_m4_19_5_i;
wire signed [`CalcTempBus]          temp_m4_19_6_r;
wire signed [`CalcTempBus]          temp_m4_19_6_i;
wire signed [`CalcTempBus]          temp_m4_19_7_r;
wire signed [`CalcTempBus]          temp_m4_19_7_i;
wire signed [`CalcTempBus]          temp_m4_19_8_r;
wire signed [`CalcTempBus]          temp_m4_19_8_i;
wire signed [`CalcTempBus]          temp_m4_19_9_r;
wire signed [`CalcTempBus]          temp_m4_19_9_i;
wire signed [`CalcTempBus]          temp_m4_19_10_r;
wire signed [`CalcTempBus]          temp_m4_19_10_i;
wire signed [`CalcTempBus]          temp_m4_19_11_r;
wire signed [`CalcTempBus]          temp_m4_19_11_i;
wire signed [`CalcTempBus]          temp_m4_19_12_r;
wire signed [`CalcTempBus]          temp_m4_19_12_i;
wire signed [`CalcTempBus]          temp_m4_19_13_r;
wire signed [`CalcTempBus]          temp_m4_19_13_i;
wire signed [`CalcTempBus]          temp_m4_19_14_r;
wire signed [`CalcTempBus]          temp_m4_19_14_i;
wire signed [`CalcTempBus]          temp_m4_19_15_r;
wire signed [`CalcTempBus]          temp_m4_19_15_i;
wire signed [`CalcTempBus]          temp_m4_19_16_r;
wire signed [`CalcTempBus]          temp_m4_19_16_i;
wire signed [`CalcTempBus]          temp_m4_19_17_r;
wire signed [`CalcTempBus]          temp_m4_19_17_i;
wire signed [`CalcTempBus]          temp_m4_19_18_r;
wire signed [`CalcTempBus]          temp_m4_19_18_i;
wire signed [`CalcTempBus]          temp_m4_19_19_r;
wire signed [`CalcTempBus]          temp_m4_19_19_i;
wire signed [`CalcTempBus]          temp_m4_19_20_r;
wire signed [`CalcTempBus]          temp_m4_19_20_i;
wire signed [`CalcTempBus]          temp_m4_19_21_r;
wire signed [`CalcTempBus]          temp_m4_19_21_i;
wire signed [`CalcTempBus]          temp_m4_19_22_r;
wire signed [`CalcTempBus]          temp_m4_19_22_i;
wire signed [`CalcTempBus]          temp_m4_19_23_r;
wire signed [`CalcTempBus]          temp_m4_19_23_i;
wire signed [`CalcTempBus]          temp_m4_19_24_r;
wire signed [`CalcTempBus]          temp_m4_19_24_i;
wire signed [`CalcTempBus]          temp_m4_19_25_r;
wire signed [`CalcTempBus]          temp_m4_19_25_i;
wire signed [`CalcTempBus]          temp_m4_19_26_r;
wire signed [`CalcTempBus]          temp_m4_19_26_i;
wire signed [`CalcTempBus]          temp_m4_19_27_r;
wire signed [`CalcTempBus]          temp_m4_19_27_i;
wire signed [`CalcTempBus]          temp_m4_19_28_r;
wire signed [`CalcTempBus]          temp_m4_19_28_i;
wire signed [`CalcTempBus]          temp_m4_19_29_r;
wire signed [`CalcTempBus]          temp_m4_19_29_i;
wire signed [`CalcTempBus]          temp_m4_19_30_r;
wire signed [`CalcTempBus]          temp_m4_19_30_i;
wire signed [`CalcTempBus]          temp_m4_19_31_r;
wire signed [`CalcTempBus]          temp_m4_19_31_i;
wire signed [`CalcTempBus]          temp_m4_19_32_r;
wire signed [`CalcTempBus]          temp_m4_19_32_i;
wire signed [`CalcTempBus]          temp_m4_20_1_r;
wire signed [`CalcTempBus]          temp_m4_20_1_i;
wire signed [`CalcTempBus]          temp_m4_20_2_r;
wire signed [`CalcTempBus]          temp_m4_20_2_i;
wire signed [`CalcTempBus]          temp_m4_20_3_r;
wire signed [`CalcTempBus]          temp_m4_20_3_i;
wire signed [`CalcTempBus]          temp_m4_20_4_r;
wire signed [`CalcTempBus]          temp_m4_20_4_i;
wire signed [`CalcTempBus]          temp_m4_20_5_r;
wire signed [`CalcTempBus]          temp_m4_20_5_i;
wire signed [`CalcTempBus]          temp_m4_20_6_r;
wire signed [`CalcTempBus]          temp_m4_20_6_i;
wire signed [`CalcTempBus]          temp_m4_20_7_r;
wire signed [`CalcTempBus]          temp_m4_20_7_i;
wire signed [`CalcTempBus]          temp_m4_20_8_r;
wire signed [`CalcTempBus]          temp_m4_20_8_i;
wire signed [`CalcTempBus]          temp_m4_20_9_r;
wire signed [`CalcTempBus]          temp_m4_20_9_i;
wire signed [`CalcTempBus]          temp_m4_20_10_r;
wire signed [`CalcTempBus]          temp_m4_20_10_i;
wire signed [`CalcTempBus]          temp_m4_20_11_r;
wire signed [`CalcTempBus]          temp_m4_20_11_i;
wire signed [`CalcTempBus]          temp_m4_20_12_r;
wire signed [`CalcTempBus]          temp_m4_20_12_i;
wire signed [`CalcTempBus]          temp_m4_20_13_r;
wire signed [`CalcTempBus]          temp_m4_20_13_i;
wire signed [`CalcTempBus]          temp_m4_20_14_r;
wire signed [`CalcTempBus]          temp_m4_20_14_i;
wire signed [`CalcTempBus]          temp_m4_20_15_r;
wire signed [`CalcTempBus]          temp_m4_20_15_i;
wire signed [`CalcTempBus]          temp_m4_20_16_r;
wire signed [`CalcTempBus]          temp_m4_20_16_i;
wire signed [`CalcTempBus]          temp_m4_20_17_r;
wire signed [`CalcTempBus]          temp_m4_20_17_i;
wire signed [`CalcTempBus]          temp_m4_20_18_r;
wire signed [`CalcTempBus]          temp_m4_20_18_i;
wire signed [`CalcTempBus]          temp_m4_20_19_r;
wire signed [`CalcTempBus]          temp_m4_20_19_i;
wire signed [`CalcTempBus]          temp_m4_20_20_r;
wire signed [`CalcTempBus]          temp_m4_20_20_i;
wire signed [`CalcTempBus]          temp_m4_20_21_r;
wire signed [`CalcTempBus]          temp_m4_20_21_i;
wire signed [`CalcTempBus]          temp_m4_20_22_r;
wire signed [`CalcTempBus]          temp_m4_20_22_i;
wire signed [`CalcTempBus]          temp_m4_20_23_r;
wire signed [`CalcTempBus]          temp_m4_20_23_i;
wire signed [`CalcTempBus]          temp_m4_20_24_r;
wire signed [`CalcTempBus]          temp_m4_20_24_i;
wire signed [`CalcTempBus]          temp_m4_20_25_r;
wire signed [`CalcTempBus]          temp_m4_20_25_i;
wire signed [`CalcTempBus]          temp_m4_20_26_r;
wire signed [`CalcTempBus]          temp_m4_20_26_i;
wire signed [`CalcTempBus]          temp_m4_20_27_r;
wire signed [`CalcTempBus]          temp_m4_20_27_i;
wire signed [`CalcTempBus]          temp_m4_20_28_r;
wire signed [`CalcTempBus]          temp_m4_20_28_i;
wire signed [`CalcTempBus]          temp_m4_20_29_r;
wire signed [`CalcTempBus]          temp_m4_20_29_i;
wire signed [`CalcTempBus]          temp_m4_20_30_r;
wire signed [`CalcTempBus]          temp_m4_20_30_i;
wire signed [`CalcTempBus]          temp_m4_20_31_r;
wire signed [`CalcTempBus]          temp_m4_20_31_i;
wire signed [`CalcTempBus]          temp_m4_20_32_r;
wire signed [`CalcTempBus]          temp_m4_20_32_i;
wire signed [`CalcTempBus]          temp_m4_21_1_r;
wire signed [`CalcTempBus]          temp_m4_21_1_i;
wire signed [`CalcTempBus]          temp_m4_21_2_r;
wire signed [`CalcTempBus]          temp_m4_21_2_i;
wire signed [`CalcTempBus]          temp_m4_21_3_r;
wire signed [`CalcTempBus]          temp_m4_21_3_i;
wire signed [`CalcTempBus]          temp_m4_21_4_r;
wire signed [`CalcTempBus]          temp_m4_21_4_i;
wire signed [`CalcTempBus]          temp_m4_21_5_r;
wire signed [`CalcTempBus]          temp_m4_21_5_i;
wire signed [`CalcTempBus]          temp_m4_21_6_r;
wire signed [`CalcTempBus]          temp_m4_21_6_i;
wire signed [`CalcTempBus]          temp_m4_21_7_r;
wire signed [`CalcTempBus]          temp_m4_21_7_i;
wire signed [`CalcTempBus]          temp_m4_21_8_r;
wire signed [`CalcTempBus]          temp_m4_21_8_i;
wire signed [`CalcTempBus]          temp_m4_21_9_r;
wire signed [`CalcTempBus]          temp_m4_21_9_i;
wire signed [`CalcTempBus]          temp_m4_21_10_r;
wire signed [`CalcTempBus]          temp_m4_21_10_i;
wire signed [`CalcTempBus]          temp_m4_21_11_r;
wire signed [`CalcTempBus]          temp_m4_21_11_i;
wire signed [`CalcTempBus]          temp_m4_21_12_r;
wire signed [`CalcTempBus]          temp_m4_21_12_i;
wire signed [`CalcTempBus]          temp_m4_21_13_r;
wire signed [`CalcTempBus]          temp_m4_21_13_i;
wire signed [`CalcTempBus]          temp_m4_21_14_r;
wire signed [`CalcTempBus]          temp_m4_21_14_i;
wire signed [`CalcTempBus]          temp_m4_21_15_r;
wire signed [`CalcTempBus]          temp_m4_21_15_i;
wire signed [`CalcTempBus]          temp_m4_21_16_r;
wire signed [`CalcTempBus]          temp_m4_21_16_i;
wire signed [`CalcTempBus]          temp_m4_21_17_r;
wire signed [`CalcTempBus]          temp_m4_21_17_i;
wire signed [`CalcTempBus]          temp_m4_21_18_r;
wire signed [`CalcTempBus]          temp_m4_21_18_i;
wire signed [`CalcTempBus]          temp_m4_21_19_r;
wire signed [`CalcTempBus]          temp_m4_21_19_i;
wire signed [`CalcTempBus]          temp_m4_21_20_r;
wire signed [`CalcTempBus]          temp_m4_21_20_i;
wire signed [`CalcTempBus]          temp_m4_21_21_r;
wire signed [`CalcTempBus]          temp_m4_21_21_i;
wire signed [`CalcTempBus]          temp_m4_21_22_r;
wire signed [`CalcTempBus]          temp_m4_21_22_i;
wire signed [`CalcTempBus]          temp_m4_21_23_r;
wire signed [`CalcTempBus]          temp_m4_21_23_i;
wire signed [`CalcTempBus]          temp_m4_21_24_r;
wire signed [`CalcTempBus]          temp_m4_21_24_i;
wire signed [`CalcTempBus]          temp_m4_21_25_r;
wire signed [`CalcTempBus]          temp_m4_21_25_i;
wire signed [`CalcTempBus]          temp_m4_21_26_r;
wire signed [`CalcTempBus]          temp_m4_21_26_i;
wire signed [`CalcTempBus]          temp_m4_21_27_r;
wire signed [`CalcTempBus]          temp_m4_21_27_i;
wire signed [`CalcTempBus]          temp_m4_21_28_r;
wire signed [`CalcTempBus]          temp_m4_21_28_i;
wire signed [`CalcTempBus]          temp_m4_21_29_r;
wire signed [`CalcTempBus]          temp_m4_21_29_i;
wire signed [`CalcTempBus]          temp_m4_21_30_r;
wire signed [`CalcTempBus]          temp_m4_21_30_i;
wire signed [`CalcTempBus]          temp_m4_21_31_r;
wire signed [`CalcTempBus]          temp_m4_21_31_i;
wire signed [`CalcTempBus]          temp_m4_21_32_r;
wire signed [`CalcTempBus]          temp_m4_21_32_i;
wire signed [`CalcTempBus]          temp_m4_22_1_r;
wire signed [`CalcTempBus]          temp_m4_22_1_i;
wire signed [`CalcTempBus]          temp_m4_22_2_r;
wire signed [`CalcTempBus]          temp_m4_22_2_i;
wire signed [`CalcTempBus]          temp_m4_22_3_r;
wire signed [`CalcTempBus]          temp_m4_22_3_i;
wire signed [`CalcTempBus]          temp_m4_22_4_r;
wire signed [`CalcTempBus]          temp_m4_22_4_i;
wire signed [`CalcTempBus]          temp_m4_22_5_r;
wire signed [`CalcTempBus]          temp_m4_22_5_i;
wire signed [`CalcTempBus]          temp_m4_22_6_r;
wire signed [`CalcTempBus]          temp_m4_22_6_i;
wire signed [`CalcTempBus]          temp_m4_22_7_r;
wire signed [`CalcTempBus]          temp_m4_22_7_i;
wire signed [`CalcTempBus]          temp_m4_22_8_r;
wire signed [`CalcTempBus]          temp_m4_22_8_i;
wire signed [`CalcTempBus]          temp_m4_22_9_r;
wire signed [`CalcTempBus]          temp_m4_22_9_i;
wire signed [`CalcTempBus]          temp_m4_22_10_r;
wire signed [`CalcTempBus]          temp_m4_22_10_i;
wire signed [`CalcTempBus]          temp_m4_22_11_r;
wire signed [`CalcTempBus]          temp_m4_22_11_i;
wire signed [`CalcTempBus]          temp_m4_22_12_r;
wire signed [`CalcTempBus]          temp_m4_22_12_i;
wire signed [`CalcTempBus]          temp_m4_22_13_r;
wire signed [`CalcTempBus]          temp_m4_22_13_i;
wire signed [`CalcTempBus]          temp_m4_22_14_r;
wire signed [`CalcTempBus]          temp_m4_22_14_i;
wire signed [`CalcTempBus]          temp_m4_22_15_r;
wire signed [`CalcTempBus]          temp_m4_22_15_i;
wire signed [`CalcTempBus]          temp_m4_22_16_r;
wire signed [`CalcTempBus]          temp_m4_22_16_i;
wire signed [`CalcTempBus]          temp_m4_22_17_r;
wire signed [`CalcTempBus]          temp_m4_22_17_i;
wire signed [`CalcTempBus]          temp_m4_22_18_r;
wire signed [`CalcTempBus]          temp_m4_22_18_i;
wire signed [`CalcTempBus]          temp_m4_22_19_r;
wire signed [`CalcTempBus]          temp_m4_22_19_i;
wire signed [`CalcTempBus]          temp_m4_22_20_r;
wire signed [`CalcTempBus]          temp_m4_22_20_i;
wire signed [`CalcTempBus]          temp_m4_22_21_r;
wire signed [`CalcTempBus]          temp_m4_22_21_i;
wire signed [`CalcTempBus]          temp_m4_22_22_r;
wire signed [`CalcTempBus]          temp_m4_22_22_i;
wire signed [`CalcTempBus]          temp_m4_22_23_r;
wire signed [`CalcTempBus]          temp_m4_22_23_i;
wire signed [`CalcTempBus]          temp_m4_22_24_r;
wire signed [`CalcTempBus]          temp_m4_22_24_i;
wire signed [`CalcTempBus]          temp_m4_22_25_r;
wire signed [`CalcTempBus]          temp_m4_22_25_i;
wire signed [`CalcTempBus]          temp_m4_22_26_r;
wire signed [`CalcTempBus]          temp_m4_22_26_i;
wire signed [`CalcTempBus]          temp_m4_22_27_r;
wire signed [`CalcTempBus]          temp_m4_22_27_i;
wire signed [`CalcTempBus]          temp_m4_22_28_r;
wire signed [`CalcTempBus]          temp_m4_22_28_i;
wire signed [`CalcTempBus]          temp_m4_22_29_r;
wire signed [`CalcTempBus]          temp_m4_22_29_i;
wire signed [`CalcTempBus]          temp_m4_22_30_r;
wire signed [`CalcTempBus]          temp_m4_22_30_i;
wire signed [`CalcTempBus]          temp_m4_22_31_r;
wire signed [`CalcTempBus]          temp_m4_22_31_i;
wire signed [`CalcTempBus]          temp_m4_22_32_r;
wire signed [`CalcTempBus]          temp_m4_22_32_i;
wire signed [`CalcTempBus]          temp_m4_23_1_r;
wire signed [`CalcTempBus]          temp_m4_23_1_i;
wire signed [`CalcTempBus]          temp_m4_23_2_r;
wire signed [`CalcTempBus]          temp_m4_23_2_i;
wire signed [`CalcTempBus]          temp_m4_23_3_r;
wire signed [`CalcTempBus]          temp_m4_23_3_i;
wire signed [`CalcTempBus]          temp_m4_23_4_r;
wire signed [`CalcTempBus]          temp_m4_23_4_i;
wire signed [`CalcTempBus]          temp_m4_23_5_r;
wire signed [`CalcTempBus]          temp_m4_23_5_i;
wire signed [`CalcTempBus]          temp_m4_23_6_r;
wire signed [`CalcTempBus]          temp_m4_23_6_i;
wire signed [`CalcTempBus]          temp_m4_23_7_r;
wire signed [`CalcTempBus]          temp_m4_23_7_i;
wire signed [`CalcTempBus]          temp_m4_23_8_r;
wire signed [`CalcTempBus]          temp_m4_23_8_i;
wire signed [`CalcTempBus]          temp_m4_23_9_r;
wire signed [`CalcTempBus]          temp_m4_23_9_i;
wire signed [`CalcTempBus]          temp_m4_23_10_r;
wire signed [`CalcTempBus]          temp_m4_23_10_i;
wire signed [`CalcTempBus]          temp_m4_23_11_r;
wire signed [`CalcTempBus]          temp_m4_23_11_i;
wire signed [`CalcTempBus]          temp_m4_23_12_r;
wire signed [`CalcTempBus]          temp_m4_23_12_i;
wire signed [`CalcTempBus]          temp_m4_23_13_r;
wire signed [`CalcTempBus]          temp_m4_23_13_i;
wire signed [`CalcTempBus]          temp_m4_23_14_r;
wire signed [`CalcTempBus]          temp_m4_23_14_i;
wire signed [`CalcTempBus]          temp_m4_23_15_r;
wire signed [`CalcTempBus]          temp_m4_23_15_i;
wire signed [`CalcTempBus]          temp_m4_23_16_r;
wire signed [`CalcTempBus]          temp_m4_23_16_i;
wire signed [`CalcTempBus]          temp_m4_23_17_r;
wire signed [`CalcTempBus]          temp_m4_23_17_i;
wire signed [`CalcTempBus]          temp_m4_23_18_r;
wire signed [`CalcTempBus]          temp_m4_23_18_i;
wire signed [`CalcTempBus]          temp_m4_23_19_r;
wire signed [`CalcTempBus]          temp_m4_23_19_i;
wire signed [`CalcTempBus]          temp_m4_23_20_r;
wire signed [`CalcTempBus]          temp_m4_23_20_i;
wire signed [`CalcTempBus]          temp_m4_23_21_r;
wire signed [`CalcTempBus]          temp_m4_23_21_i;
wire signed [`CalcTempBus]          temp_m4_23_22_r;
wire signed [`CalcTempBus]          temp_m4_23_22_i;
wire signed [`CalcTempBus]          temp_m4_23_23_r;
wire signed [`CalcTempBus]          temp_m4_23_23_i;
wire signed [`CalcTempBus]          temp_m4_23_24_r;
wire signed [`CalcTempBus]          temp_m4_23_24_i;
wire signed [`CalcTempBus]          temp_m4_23_25_r;
wire signed [`CalcTempBus]          temp_m4_23_25_i;
wire signed [`CalcTempBus]          temp_m4_23_26_r;
wire signed [`CalcTempBus]          temp_m4_23_26_i;
wire signed [`CalcTempBus]          temp_m4_23_27_r;
wire signed [`CalcTempBus]          temp_m4_23_27_i;
wire signed [`CalcTempBus]          temp_m4_23_28_r;
wire signed [`CalcTempBus]          temp_m4_23_28_i;
wire signed [`CalcTempBus]          temp_m4_23_29_r;
wire signed [`CalcTempBus]          temp_m4_23_29_i;
wire signed [`CalcTempBus]          temp_m4_23_30_r;
wire signed [`CalcTempBus]          temp_m4_23_30_i;
wire signed [`CalcTempBus]          temp_m4_23_31_r;
wire signed [`CalcTempBus]          temp_m4_23_31_i;
wire signed [`CalcTempBus]          temp_m4_23_32_r;
wire signed [`CalcTempBus]          temp_m4_23_32_i;
wire signed [`CalcTempBus]          temp_m4_24_1_r;
wire signed [`CalcTempBus]          temp_m4_24_1_i;
wire signed [`CalcTempBus]          temp_m4_24_2_r;
wire signed [`CalcTempBus]          temp_m4_24_2_i;
wire signed [`CalcTempBus]          temp_m4_24_3_r;
wire signed [`CalcTempBus]          temp_m4_24_3_i;
wire signed [`CalcTempBus]          temp_m4_24_4_r;
wire signed [`CalcTempBus]          temp_m4_24_4_i;
wire signed [`CalcTempBus]          temp_m4_24_5_r;
wire signed [`CalcTempBus]          temp_m4_24_5_i;
wire signed [`CalcTempBus]          temp_m4_24_6_r;
wire signed [`CalcTempBus]          temp_m4_24_6_i;
wire signed [`CalcTempBus]          temp_m4_24_7_r;
wire signed [`CalcTempBus]          temp_m4_24_7_i;
wire signed [`CalcTempBus]          temp_m4_24_8_r;
wire signed [`CalcTempBus]          temp_m4_24_8_i;
wire signed [`CalcTempBus]          temp_m4_24_9_r;
wire signed [`CalcTempBus]          temp_m4_24_9_i;
wire signed [`CalcTempBus]          temp_m4_24_10_r;
wire signed [`CalcTempBus]          temp_m4_24_10_i;
wire signed [`CalcTempBus]          temp_m4_24_11_r;
wire signed [`CalcTempBus]          temp_m4_24_11_i;
wire signed [`CalcTempBus]          temp_m4_24_12_r;
wire signed [`CalcTempBus]          temp_m4_24_12_i;
wire signed [`CalcTempBus]          temp_m4_24_13_r;
wire signed [`CalcTempBus]          temp_m4_24_13_i;
wire signed [`CalcTempBus]          temp_m4_24_14_r;
wire signed [`CalcTempBus]          temp_m4_24_14_i;
wire signed [`CalcTempBus]          temp_m4_24_15_r;
wire signed [`CalcTempBus]          temp_m4_24_15_i;
wire signed [`CalcTempBus]          temp_m4_24_16_r;
wire signed [`CalcTempBus]          temp_m4_24_16_i;
wire signed [`CalcTempBus]          temp_m4_24_17_r;
wire signed [`CalcTempBus]          temp_m4_24_17_i;
wire signed [`CalcTempBus]          temp_m4_24_18_r;
wire signed [`CalcTempBus]          temp_m4_24_18_i;
wire signed [`CalcTempBus]          temp_m4_24_19_r;
wire signed [`CalcTempBus]          temp_m4_24_19_i;
wire signed [`CalcTempBus]          temp_m4_24_20_r;
wire signed [`CalcTempBus]          temp_m4_24_20_i;
wire signed [`CalcTempBus]          temp_m4_24_21_r;
wire signed [`CalcTempBus]          temp_m4_24_21_i;
wire signed [`CalcTempBus]          temp_m4_24_22_r;
wire signed [`CalcTempBus]          temp_m4_24_22_i;
wire signed [`CalcTempBus]          temp_m4_24_23_r;
wire signed [`CalcTempBus]          temp_m4_24_23_i;
wire signed [`CalcTempBus]          temp_m4_24_24_r;
wire signed [`CalcTempBus]          temp_m4_24_24_i;
wire signed [`CalcTempBus]          temp_m4_24_25_r;
wire signed [`CalcTempBus]          temp_m4_24_25_i;
wire signed [`CalcTempBus]          temp_m4_24_26_r;
wire signed [`CalcTempBus]          temp_m4_24_26_i;
wire signed [`CalcTempBus]          temp_m4_24_27_r;
wire signed [`CalcTempBus]          temp_m4_24_27_i;
wire signed [`CalcTempBus]          temp_m4_24_28_r;
wire signed [`CalcTempBus]          temp_m4_24_28_i;
wire signed [`CalcTempBus]          temp_m4_24_29_r;
wire signed [`CalcTempBus]          temp_m4_24_29_i;
wire signed [`CalcTempBus]          temp_m4_24_30_r;
wire signed [`CalcTempBus]          temp_m4_24_30_i;
wire signed [`CalcTempBus]          temp_m4_24_31_r;
wire signed [`CalcTempBus]          temp_m4_24_31_i;
wire signed [`CalcTempBus]          temp_m4_24_32_r;
wire signed [`CalcTempBus]          temp_m4_24_32_i;
wire signed [`CalcTempBus]          temp_m4_25_1_r;
wire signed [`CalcTempBus]          temp_m4_25_1_i;
wire signed [`CalcTempBus]          temp_m4_25_2_r;
wire signed [`CalcTempBus]          temp_m4_25_2_i;
wire signed [`CalcTempBus]          temp_m4_25_3_r;
wire signed [`CalcTempBus]          temp_m4_25_3_i;
wire signed [`CalcTempBus]          temp_m4_25_4_r;
wire signed [`CalcTempBus]          temp_m4_25_4_i;
wire signed [`CalcTempBus]          temp_m4_25_5_r;
wire signed [`CalcTempBus]          temp_m4_25_5_i;
wire signed [`CalcTempBus]          temp_m4_25_6_r;
wire signed [`CalcTempBus]          temp_m4_25_6_i;
wire signed [`CalcTempBus]          temp_m4_25_7_r;
wire signed [`CalcTempBus]          temp_m4_25_7_i;
wire signed [`CalcTempBus]          temp_m4_25_8_r;
wire signed [`CalcTempBus]          temp_m4_25_8_i;
wire signed [`CalcTempBus]          temp_m4_25_9_r;
wire signed [`CalcTempBus]          temp_m4_25_9_i;
wire signed [`CalcTempBus]          temp_m4_25_10_r;
wire signed [`CalcTempBus]          temp_m4_25_10_i;
wire signed [`CalcTempBus]          temp_m4_25_11_r;
wire signed [`CalcTempBus]          temp_m4_25_11_i;
wire signed [`CalcTempBus]          temp_m4_25_12_r;
wire signed [`CalcTempBus]          temp_m4_25_12_i;
wire signed [`CalcTempBus]          temp_m4_25_13_r;
wire signed [`CalcTempBus]          temp_m4_25_13_i;
wire signed [`CalcTempBus]          temp_m4_25_14_r;
wire signed [`CalcTempBus]          temp_m4_25_14_i;
wire signed [`CalcTempBus]          temp_m4_25_15_r;
wire signed [`CalcTempBus]          temp_m4_25_15_i;
wire signed [`CalcTempBus]          temp_m4_25_16_r;
wire signed [`CalcTempBus]          temp_m4_25_16_i;
wire signed [`CalcTempBus]          temp_m4_25_17_r;
wire signed [`CalcTempBus]          temp_m4_25_17_i;
wire signed [`CalcTempBus]          temp_m4_25_18_r;
wire signed [`CalcTempBus]          temp_m4_25_18_i;
wire signed [`CalcTempBus]          temp_m4_25_19_r;
wire signed [`CalcTempBus]          temp_m4_25_19_i;
wire signed [`CalcTempBus]          temp_m4_25_20_r;
wire signed [`CalcTempBus]          temp_m4_25_20_i;
wire signed [`CalcTempBus]          temp_m4_25_21_r;
wire signed [`CalcTempBus]          temp_m4_25_21_i;
wire signed [`CalcTempBus]          temp_m4_25_22_r;
wire signed [`CalcTempBus]          temp_m4_25_22_i;
wire signed [`CalcTempBus]          temp_m4_25_23_r;
wire signed [`CalcTempBus]          temp_m4_25_23_i;
wire signed [`CalcTempBus]          temp_m4_25_24_r;
wire signed [`CalcTempBus]          temp_m4_25_24_i;
wire signed [`CalcTempBus]          temp_m4_25_25_r;
wire signed [`CalcTempBus]          temp_m4_25_25_i;
wire signed [`CalcTempBus]          temp_m4_25_26_r;
wire signed [`CalcTempBus]          temp_m4_25_26_i;
wire signed [`CalcTempBus]          temp_m4_25_27_r;
wire signed [`CalcTempBus]          temp_m4_25_27_i;
wire signed [`CalcTempBus]          temp_m4_25_28_r;
wire signed [`CalcTempBus]          temp_m4_25_28_i;
wire signed [`CalcTempBus]          temp_m4_25_29_r;
wire signed [`CalcTempBus]          temp_m4_25_29_i;
wire signed [`CalcTempBus]          temp_m4_25_30_r;
wire signed [`CalcTempBus]          temp_m4_25_30_i;
wire signed [`CalcTempBus]          temp_m4_25_31_r;
wire signed [`CalcTempBus]          temp_m4_25_31_i;
wire signed [`CalcTempBus]          temp_m4_25_32_r;
wire signed [`CalcTempBus]          temp_m4_25_32_i;
wire signed [`CalcTempBus]          temp_m4_26_1_r;
wire signed [`CalcTempBus]          temp_m4_26_1_i;
wire signed [`CalcTempBus]          temp_m4_26_2_r;
wire signed [`CalcTempBus]          temp_m4_26_2_i;
wire signed [`CalcTempBus]          temp_m4_26_3_r;
wire signed [`CalcTempBus]          temp_m4_26_3_i;
wire signed [`CalcTempBus]          temp_m4_26_4_r;
wire signed [`CalcTempBus]          temp_m4_26_4_i;
wire signed [`CalcTempBus]          temp_m4_26_5_r;
wire signed [`CalcTempBus]          temp_m4_26_5_i;
wire signed [`CalcTempBus]          temp_m4_26_6_r;
wire signed [`CalcTempBus]          temp_m4_26_6_i;
wire signed [`CalcTempBus]          temp_m4_26_7_r;
wire signed [`CalcTempBus]          temp_m4_26_7_i;
wire signed [`CalcTempBus]          temp_m4_26_8_r;
wire signed [`CalcTempBus]          temp_m4_26_8_i;
wire signed [`CalcTempBus]          temp_m4_26_9_r;
wire signed [`CalcTempBus]          temp_m4_26_9_i;
wire signed [`CalcTempBus]          temp_m4_26_10_r;
wire signed [`CalcTempBus]          temp_m4_26_10_i;
wire signed [`CalcTempBus]          temp_m4_26_11_r;
wire signed [`CalcTempBus]          temp_m4_26_11_i;
wire signed [`CalcTempBus]          temp_m4_26_12_r;
wire signed [`CalcTempBus]          temp_m4_26_12_i;
wire signed [`CalcTempBus]          temp_m4_26_13_r;
wire signed [`CalcTempBus]          temp_m4_26_13_i;
wire signed [`CalcTempBus]          temp_m4_26_14_r;
wire signed [`CalcTempBus]          temp_m4_26_14_i;
wire signed [`CalcTempBus]          temp_m4_26_15_r;
wire signed [`CalcTempBus]          temp_m4_26_15_i;
wire signed [`CalcTempBus]          temp_m4_26_16_r;
wire signed [`CalcTempBus]          temp_m4_26_16_i;
wire signed [`CalcTempBus]          temp_m4_26_17_r;
wire signed [`CalcTempBus]          temp_m4_26_17_i;
wire signed [`CalcTempBus]          temp_m4_26_18_r;
wire signed [`CalcTempBus]          temp_m4_26_18_i;
wire signed [`CalcTempBus]          temp_m4_26_19_r;
wire signed [`CalcTempBus]          temp_m4_26_19_i;
wire signed [`CalcTempBus]          temp_m4_26_20_r;
wire signed [`CalcTempBus]          temp_m4_26_20_i;
wire signed [`CalcTempBus]          temp_m4_26_21_r;
wire signed [`CalcTempBus]          temp_m4_26_21_i;
wire signed [`CalcTempBus]          temp_m4_26_22_r;
wire signed [`CalcTempBus]          temp_m4_26_22_i;
wire signed [`CalcTempBus]          temp_m4_26_23_r;
wire signed [`CalcTempBus]          temp_m4_26_23_i;
wire signed [`CalcTempBus]          temp_m4_26_24_r;
wire signed [`CalcTempBus]          temp_m4_26_24_i;
wire signed [`CalcTempBus]          temp_m4_26_25_r;
wire signed [`CalcTempBus]          temp_m4_26_25_i;
wire signed [`CalcTempBus]          temp_m4_26_26_r;
wire signed [`CalcTempBus]          temp_m4_26_26_i;
wire signed [`CalcTempBus]          temp_m4_26_27_r;
wire signed [`CalcTempBus]          temp_m4_26_27_i;
wire signed [`CalcTempBus]          temp_m4_26_28_r;
wire signed [`CalcTempBus]          temp_m4_26_28_i;
wire signed [`CalcTempBus]          temp_m4_26_29_r;
wire signed [`CalcTempBus]          temp_m4_26_29_i;
wire signed [`CalcTempBus]          temp_m4_26_30_r;
wire signed [`CalcTempBus]          temp_m4_26_30_i;
wire signed [`CalcTempBus]          temp_m4_26_31_r;
wire signed [`CalcTempBus]          temp_m4_26_31_i;
wire signed [`CalcTempBus]          temp_m4_26_32_r;
wire signed [`CalcTempBus]          temp_m4_26_32_i;
wire signed [`CalcTempBus]          temp_m4_27_1_r;
wire signed [`CalcTempBus]          temp_m4_27_1_i;
wire signed [`CalcTempBus]          temp_m4_27_2_r;
wire signed [`CalcTempBus]          temp_m4_27_2_i;
wire signed [`CalcTempBus]          temp_m4_27_3_r;
wire signed [`CalcTempBus]          temp_m4_27_3_i;
wire signed [`CalcTempBus]          temp_m4_27_4_r;
wire signed [`CalcTempBus]          temp_m4_27_4_i;
wire signed [`CalcTempBus]          temp_m4_27_5_r;
wire signed [`CalcTempBus]          temp_m4_27_5_i;
wire signed [`CalcTempBus]          temp_m4_27_6_r;
wire signed [`CalcTempBus]          temp_m4_27_6_i;
wire signed [`CalcTempBus]          temp_m4_27_7_r;
wire signed [`CalcTempBus]          temp_m4_27_7_i;
wire signed [`CalcTempBus]          temp_m4_27_8_r;
wire signed [`CalcTempBus]          temp_m4_27_8_i;
wire signed [`CalcTempBus]          temp_m4_27_9_r;
wire signed [`CalcTempBus]          temp_m4_27_9_i;
wire signed [`CalcTempBus]          temp_m4_27_10_r;
wire signed [`CalcTempBus]          temp_m4_27_10_i;
wire signed [`CalcTempBus]          temp_m4_27_11_r;
wire signed [`CalcTempBus]          temp_m4_27_11_i;
wire signed [`CalcTempBus]          temp_m4_27_12_r;
wire signed [`CalcTempBus]          temp_m4_27_12_i;
wire signed [`CalcTempBus]          temp_m4_27_13_r;
wire signed [`CalcTempBus]          temp_m4_27_13_i;
wire signed [`CalcTempBus]          temp_m4_27_14_r;
wire signed [`CalcTempBus]          temp_m4_27_14_i;
wire signed [`CalcTempBus]          temp_m4_27_15_r;
wire signed [`CalcTempBus]          temp_m4_27_15_i;
wire signed [`CalcTempBus]          temp_m4_27_16_r;
wire signed [`CalcTempBus]          temp_m4_27_16_i;
wire signed [`CalcTempBus]          temp_m4_27_17_r;
wire signed [`CalcTempBus]          temp_m4_27_17_i;
wire signed [`CalcTempBus]          temp_m4_27_18_r;
wire signed [`CalcTempBus]          temp_m4_27_18_i;
wire signed [`CalcTempBus]          temp_m4_27_19_r;
wire signed [`CalcTempBus]          temp_m4_27_19_i;
wire signed [`CalcTempBus]          temp_m4_27_20_r;
wire signed [`CalcTempBus]          temp_m4_27_20_i;
wire signed [`CalcTempBus]          temp_m4_27_21_r;
wire signed [`CalcTempBus]          temp_m4_27_21_i;
wire signed [`CalcTempBus]          temp_m4_27_22_r;
wire signed [`CalcTempBus]          temp_m4_27_22_i;
wire signed [`CalcTempBus]          temp_m4_27_23_r;
wire signed [`CalcTempBus]          temp_m4_27_23_i;
wire signed [`CalcTempBus]          temp_m4_27_24_r;
wire signed [`CalcTempBus]          temp_m4_27_24_i;
wire signed [`CalcTempBus]          temp_m4_27_25_r;
wire signed [`CalcTempBus]          temp_m4_27_25_i;
wire signed [`CalcTempBus]          temp_m4_27_26_r;
wire signed [`CalcTempBus]          temp_m4_27_26_i;
wire signed [`CalcTempBus]          temp_m4_27_27_r;
wire signed [`CalcTempBus]          temp_m4_27_27_i;
wire signed [`CalcTempBus]          temp_m4_27_28_r;
wire signed [`CalcTempBus]          temp_m4_27_28_i;
wire signed [`CalcTempBus]          temp_m4_27_29_r;
wire signed [`CalcTempBus]          temp_m4_27_29_i;
wire signed [`CalcTempBus]          temp_m4_27_30_r;
wire signed [`CalcTempBus]          temp_m4_27_30_i;
wire signed [`CalcTempBus]          temp_m4_27_31_r;
wire signed [`CalcTempBus]          temp_m4_27_31_i;
wire signed [`CalcTempBus]          temp_m4_27_32_r;
wire signed [`CalcTempBus]          temp_m4_27_32_i;
wire signed [`CalcTempBus]          temp_m4_28_1_r;
wire signed [`CalcTempBus]          temp_m4_28_1_i;
wire signed [`CalcTempBus]          temp_m4_28_2_r;
wire signed [`CalcTempBus]          temp_m4_28_2_i;
wire signed [`CalcTempBus]          temp_m4_28_3_r;
wire signed [`CalcTempBus]          temp_m4_28_3_i;
wire signed [`CalcTempBus]          temp_m4_28_4_r;
wire signed [`CalcTempBus]          temp_m4_28_4_i;
wire signed [`CalcTempBus]          temp_m4_28_5_r;
wire signed [`CalcTempBus]          temp_m4_28_5_i;
wire signed [`CalcTempBus]          temp_m4_28_6_r;
wire signed [`CalcTempBus]          temp_m4_28_6_i;
wire signed [`CalcTempBus]          temp_m4_28_7_r;
wire signed [`CalcTempBus]          temp_m4_28_7_i;
wire signed [`CalcTempBus]          temp_m4_28_8_r;
wire signed [`CalcTempBus]          temp_m4_28_8_i;
wire signed [`CalcTempBus]          temp_m4_28_9_r;
wire signed [`CalcTempBus]          temp_m4_28_9_i;
wire signed [`CalcTempBus]          temp_m4_28_10_r;
wire signed [`CalcTempBus]          temp_m4_28_10_i;
wire signed [`CalcTempBus]          temp_m4_28_11_r;
wire signed [`CalcTempBus]          temp_m4_28_11_i;
wire signed [`CalcTempBus]          temp_m4_28_12_r;
wire signed [`CalcTempBus]          temp_m4_28_12_i;
wire signed [`CalcTempBus]          temp_m4_28_13_r;
wire signed [`CalcTempBus]          temp_m4_28_13_i;
wire signed [`CalcTempBus]          temp_m4_28_14_r;
wire signed [`CalcTempBus]          temp_m4_28_14_i;
wire signed [`CalcTempBus]          temp_m4_28_15_r;
wire signed [`CalcTempBus]          temp_m4_28_15_i;
wire signed [`CalcTempBus]          temp_m4_28_16_r;
wire signed [`CalcTempBus]          temp_m4_28_16_i;
wire signed [`CalcTempBus]          temp_m4_28_17_r;
wire signed [`CalcTempBus]          temp_m4_28_17_i;
wire signed [`CalcTempBus]          temp_m4_28_18_r;
wire signed [`CalcTempBus]          temp_m4_28_18_i;
wire signed [`CalcTempBus]          temp_m4_28_19_r;
wire signed [`CalcTempBus]          temp_m4_28_19_i;
wire signed [`CalcTempBus]          temp_m4_28_20_r;
wire signed [`CalcTempBus]          temp_m4_28_20_i;
wire signed [`CalcTempBus]          temp_m4_28_21_r;
wire signed [`CalcTempBus]          temp_m4_28_21_i;
wire signed [`CalcTempBus]          temp_m4_28_22_r;
wire signed [`CalcTempBus]          temp_m4_28_22_i;
wire signed [`CalcTempBus]          temp_m4_28_23_r;
wire signed [`CalcTempBus]          temp_m4_28_23_i;
wire signed [`CalcTempBus]          temp_m4_28_24_r;
wire signed [`CalcTempBus]          temp_m4_28_24_i;
wire signed [`CalcTempBus]          temp_m4_28_25_r;
wire signed [`CalcTempBus]          temp_m4_28_25_i;
wire signed [`CalcTempBus]          temp_m4_28_26_r;
wire signed [`CalcTempBus]          temp_m4_28_26_i;
wire signed [`CalcTempBus]          temp_m4_28_27_r;
wire signed [`CalcTempBus]          temp_m4_28_27_i;
wire signed [`CalcTempBus]          temp_m4_28_28_r;
wire signed [`CalcTempBus]          temp_m4_28_28_i;
wire signed [`CalcTempBus]          temp_m4_28_29_r;
wire signed [`CalcTempBus]          temp_m4_28_29_i;
wire signed [`CalcTempBus]          temp_m4_28_30_r;
wire signed [`CalcTempBus]          temp_m4_28_30_i;
wire signed [`CalcTempBus]          temp_m4_28_31_r;
wire signed [`CalcTempBus]          temp_m4_28_31_i;
wire signed [`CalcTempBus]          temp_m4_28_32_r;
wire signed [`CalcTempBus]          temp_m4_28_32_i;
wire signed [`CalcTempBus]          temp_m4_29_1_r;
wire signed [`CalcTempBus]          temp_m4_29_1_i;
wire signed [`CalcTempBus]          temp_m4_29_2_r;
wire signed [`CalcTempBus]          temp_m4_29_2_i;
wire signed [`CalcTempBus]          temp_m4_29_3_r;
wire signed [`CalcTempBus]          temp_m4_29_3_i;
wire signed [`CalcTempBus]          temp_m4_29_4_r;
wire signed [`CalcTempBus]          temp_m4_29_4_i;
wire signed [`CalcTempBus]          temp_m4_29_5_r;
wire signed [`CalcTempBus]          temp_m4_29_5_i;
wire signed [`CalcTempBus]          temp_m4_29_6_r;
wire signed [`CalcTempBus]          temp_m4_29_6_i;
wire signed [`CalcTempBus]          temp_m4_29_7_r;
wire signed [`CalcTempBus]          temp_m4_29_7_i;
wire signed [`CalcTempBus]          temp_m4_29_8_r;
wire signed [`CalcTempBus]          temp_m4_29_8_i;
wire signed [`CalcTempBus]          temp_m4_29_9_r;
wire signed [`CalcTempBus]          temp_m4_29_9_i;
wire signed [`CalcTempBus]          temp_m4_29_10_r;
wire signed [`CalcTempBus]          temp_m4_29_10_i;
wire signed [`CalcTempBus]          temp_m4_29_11_r;
wire signed [`CalcTempBus]          temp_m4_29_11_i;
wire signed [`CalcTempBus]          temp_m4_29_12_r;
wire signed [`CalcTempBus]          temp_m4_29_12_i;
wire signed [`CalcTempBus]          temp_m4_29_13_r;
wire signed [`CalcTempBus]          temp_m4_29_13_i;
wire signed [`CalcTempBus]          temp_m4_29_14_r;
wire signed [`CalcTempBus]          temp_m4_29_14_i;
wire signed [`CalcTempBus]          temp_m4_29_15_r;
wire signed [`CalcTempBus]          temp_m4_29_15_i;
wire signed [`CalcTempBus]          temp_m4_29_16_r;
wire signed [`CalcTempBus]          temp_m4_29_16_i;
wire signed [`CalcTempBus]          temp_m4_29_17_r;
wire signed [`CalcTempBus]          temp_m4_29_17_i;
wire signed [`CalcTempBus]          temp_m4_29_18_r;
wire signed [`CalcTempBus]          temp_m4_29_18_i;
wire signed [`CalcTempBus]          temp_m4_29_19_r;
wire signed [`CalcTempBus]          temp_m4_29_19_i;
wire signed [`CalcTempBus]          temp_m4_29_20_r;
wire signed [`CalcTempBus]          temp_m4_29_20_i;
wire signed [`CalcTempBus]          temp_m4_29_21_r;
wire signed [`CalcTempBus]          temp_m4_29_21_i;
wire signed [`CalcTempBus]          temp_m4_29_22_r;
wire signed [`CalcTempBus]          temp_m4_29_22_i;
wire signed [`CalcTempBus]          temp_m4_29_23_r;
wire signed [`CalcTempBus]          temp_m4_29_23_i;
wire signed [`CalcTempBus]          temp_m4_29_24_r;
wire signed [`CalcTempBus]          temp_m4_29_24_i;
wire signed [`CalcTempBus]          temp_m4_29_25_r;
wire signed [`CalcTempBus]          temp_m4_29_25_i;
wire signed [`CalcTempBus]          temp_m4_29_26_r;
wire signed [`CalcTempBus]          temp_m4_29_26_i;
wire signed [`CalcTempBus]          temp_m4_29_27_r;
wire signed [`CalcTempBus]          temp_m4_29_27_i;
wire signed [`CalcTempBus]          temp_m4_29_28_r;
wire signed [`CalcTempBus]          temp_m4_29_28_i;
wire signed [`CalcTempBus]          temp_m4_29_29_r;
wire signed [`CalcTempBus]          temp_m4_29_29_i;
wire signed [`CalcTempBus]          temp_m4_29_30_r;
wire signed [`CalcTempBus]          temp_m4_29_30_i;
wire signed [`CalcTempBus]          temp_m4_29_31_r;
wire signed [`CalcTempBus]          temp_m4_29_31_i;
wire signed [`CalcTempBus]          temp_m4_29_32_r;
wire signed [`CalcTempBus]          temp_m4_29_32_i;
wire signed [`CalcTempBus]          temp_m4_30_1_r;
wire signed [`CalcTempBus]          temp_m4_30_1_i;
wire signed [`CalcTempBus]          temp_m4_30_2_r;
wire signed [`CalcTempBus]          temp_m4_30_2_i;
wire signed [`CalcTempBus]          temp_m4_30_3_r;
wire signed [`CalcTempBus]          temp_m4_30_3_i;
wire signed [`CalcTempBus]          temp_m4_30_4_r;
wire signed [`CalcTempBus]          temp_m4_30_4_i;
wire signed [`CalcTempBus]          temp_m4_30_5_r;
wire signed [`CalcTempBus]          temp_m4_30_5_i;
wire signed [`CalcTempBus]          temp_m4_30_6_r;
wire signed [`CalcTempBus]          temp_m4_30_6_i;
wire signed [`CalcTempBus]          temp_m4_30_7_r;
wire signed [`CalcTempBus]          temp_m4_30_7_i;
wire signed [`CalcTempBus]          temp_m4_30_8_r;
wire signed [`CalcTempBus]          temp_m4_30_8_i;
wire signed [`CalcTempBus]          temp_m4_30_9_r;
wire signed [`CalcTempBus]          temp_m4_30_9_i;
wire signed [`CalcTempBus]          temp_m4_30_10_r;
wire signed [`CalcTempBus]          temp_m4_30_10_i;
wire signed [`CalcTempBus]          temp_m4_30_11_r;
wire signed [`CalcTempBus]          temp_m4_30_11_i;
wire signed [`CalcTempBus]          temp_m4_30_12_r;
wire signed [`CalcTempBus]          temp_m4_30_12_i;
wire signed [`CalcTempBus]          temp_m4_30_13_r;
wire signed [`CalcTempBus]          temp_m4_30_13_i;
wire signed [`CalcTempBus]          temp_m4_30_14_r;
wire signed [`CalcTempBus]          temp_m4_30_14_i;
wire signed [`CalcTempBus]          temp_m4_30_15_r;
wire signed [`CalcTempBus]          temp_m4_30_15_i;
wire signed [`CalcTempBus]          temp_m4_30_16_r;
wire signed [`CalcTempBus]          temp_m4_30_16_i;
wire signed [`CalcTempBus]          temp_m4_30_17_r;
wire signed [`CalcTempBus]          temp_m4_30_17_i;
wire signed [`CalcTempBus]          temp_m4_30_18_r;
wire signed [`CalcTempBus]          temp_m4_30_18_i;
wire signed [`CalcTempBus]          temp_m4_30_19_r;
wire signed [`CalcTempBus]          temp_m4_30_19_i;
wire signed [`CalcTempBus]          temp_m4_30_20_r;
wire signed [`CalcTempBus]          temp_m4_30_20_i;
wire signed [`CalcTempBus]          temp_m4_30_21_r;
wire signed [`CalcTempBus]          temp_m4_30_21_i;
wire signed [`CalcTempBus]          temp_m4_30_22_r;
wire signed [`CalcTempBus]          temp_m4_30_22_i;
wire signed [`CalcTempBus]          temp_m4_30_23_r;
wire signed [`CalcTempBus]          temp_m4_30_23_i;
wire signed [`CalcTempBus]          temp_m4_30_24_r;
wire signed [`CalcTempBus]          temp_m4_30_24_i;
wire signed [`CalcTempBus]          temp_m4_30_25_r;
wire signed [`CalcTempBus]          temp_m4_30_25_i;
wire signed [`CalcTempBus]          temp_m4_30_26_r;
wire signed [`CalcTempBus]          temp_m4_30_26_i;
wire signed [`CalcTempBus]          temp_m4_30_27_r;
wire signed [`CalcTempBus]          temp_m4_30_27_i;
wire signed [`CalcTempBus]          temp_m4_30_28_r;
wire signed [`CalcTempBus]          temp_m4_30_28_i;
wire signed [`CalcTempBus]          temp_m4_30_29_r;
wire signed [`CalcTempBus]          temp_m4_30_29_i;
wire signed [`CalcTempBus]          temp_m4_30_30_r;
wire signed [`CalcTempBus]          temp_m4_30_30_i;
wire signed [`CalcTempBus]          temp_m4_30_31_r;
wire signed [`CalcTempBus]          temp_m4_30_31_i;
wire signed [`CalcTempBus]          temp_m4_30_32_r;
wire signed [`CalcTempBus]          temp_m4_30_32_i;
wire signed [`CalcTempBus]          temp_m4_31_1_r;
wire signed [`CalcTempBus]          temp_m4_31_1_i;
wire signed [`CalcTempBus]          temp_m4_31_2_r;
wire signed [`CalcTempBus]          temp_m4_31_2_i;
wire signed [`CalcTempBus]          temp_m4_31_3_r;
wire signed [`CalcTempBus]          temp_m4_31_3_i;
wire signed [`CalcTempBus]          temp_m4_31_4_r;
wire signed [`CalcTempBus]          temp_m4_31_4_i;
wire signed [`CalcTempBus]          temp_m4_31_5_r;
wire signed [`CalcTempBus]          temp_m4_31_5_i;
wire signed [`CalcTempBus]          temp_m4_31_6_r;
wire signed [`CalcTempBus]          temp_m4_31_6_i;
wire signed [`CalcTempBus]          temp_m4_31_7_r;
wire signed [`CalcTempBus]          temp_m4_31_7_i;
wire signed [`CalcTempBus]          temp_m4_31_8_r;
wire signed [`CalcTempBus]          temp_m4_31_8_i;
wire signed [`CalcTempBus]          temp_m4_31_9_r;
wire signed [`CalcTempBus]          temp_m4_31_9_i;
wire signed [`CalcTempBus]          temp_m4_31_10_r;
wire signed [`CalcTempBus]          temp_m4_31_10_i;
wire signed [`CalcTempBus]          temp_m4_31_11_r;
wire signed [`CalcTempBus]          temp_m4_31_11_i;
wire signed [`CalcTempBus]          temp_m4_31_12_r;
wire signed [`CalcTempBus]          temp_m4_31_12_i;
wire signed [`CalcTempBus]          temp_m4_31_13_r;
wire signed [`CalcTempBus]          temp_m4_31_13_i;
wire signed [`CalcTempBus]          temp_m4_31_14_r;
wire signed [`CalcTempBus]          temp_m4_31_14_i;
wire signed [`CalcTempBus]          temp_m4_31_15_r;
wire signed [`CalcTempBus]          temp_m4_31_15_i;
wire signed [`CalcTempBus]          temp_m4_31_16_r;
wire signed [`CalcTempBus]          temp_m4_31_16_i;
wire signed [`CalcTempBus]          temp_m4_31_17_r;
wire signed [`CalcTempBus]          temp_m4_31_17_i;
wire signed [`CalcTempBus]          temp_m4_31_18_r;
wire signed [`CalcTempBus]          temp_m4_31_18_i;
wire signed [`CalcTempBus]          temp_m4_31_19_r;
wire signed [`CalcTempBus]          temp_m4_31_19_i;
wire signed [`CalcTempBus]          temp_m4_31_20_r;
wire signed [`CalcTempBus]          temp_m4_31_20_i;
wire signed [`CalcTempBus]          temp_m4_31_21_r;
wire signed [`CalcTempBus]          temp_m4_31_21_i;
wire signed [`CalcTempBus]          temp_m4_31_22_r;
wire signed [`CalcTempBus]          temp_m4_31_22_i;
wire signed [`CalcTempBus]          temp_m4_31_23_r;
wire signed [`CalcTempBus]          temp_m4_31_23_i;
wire signed [`CalcTempBus]          temp_m4_31_24_r;
wire signed [`CalcTempBus]          temp_m4_31_24_i;
wire signed [`CalcTempBus]          temp_m4_31_25_r;
wire signed [`CalcTempBus]          temp_m4_31_25_i;
wire signed [`CalcTempBus]          temp_m4_31_26_r;
wire signed [`CalcTempBus]          temp_m4_31_26_i;
wire signed [`CalcTempBus]          temp_m4_31_27_r;
wire signed [`CalcTempBus]          temp_m4_31_27_i;
wire signed [`CalcTempBus]          temp_m4_31_28_r;
wire signed [`CalcTempBus]          temp_m4_31_28_i;
wire signed [`CalcTempBus]          temp_m4_31_29_r;
wire signed [`CalcTempBus]          temp_m4_31_29_i;
wire signed [`CalcTempBus]          temp_m4_31_30_r;
wire signed [`CalcTempBus]          temp_m4_31_30_i;
wire signed [`CalcTempBus]          temp_m4_31_31_r;
wire signed [`CalcTempBus]          temp_m4_31_31_i;
wire signed [`CalcTempBus]          temp_m4_31_32_r;
wire signed [`CalcTempBus]          temp_m4_31_32_i;
wire signed [`CalcTempBus]          temp_m4_32_1_r;
wire signed [`CalcTempBus]          temp_m4_32_1_i;
wire signed [`CalcTempBus]          temp_m4_32_2_r;
wire signed [`CalcTempBus]          temp_m4_32_2_i;
wire signed [`CalcTempBus]          temp_m4_32_3_r;
wire signed [`CalcTempBus]          temp_m4_32_3_i;
wire signed [`CalcTempBus]          temp_m4_32_4_r;
wire signed [`CalcTempBus]          temp_m4_32_4_i;
wire signed [`CalcTempBus]          temp_m4_32_5_r;
wire signed [`CalcTempBus]          temp_m4_32_5_i;
wire signed [`CalcTempBus]          temp_m4_32_6_r;
wire signed [`CalcTempBus]          temp_m4_32_6_i;
wire signed [`CalcTempBus]          temp_m4_32_7_r;
wire signed [`CalcTempBus]          temp_m4_32_7_i;
wire signed [`CalcTempBus]          temp_m4_32_8_r;
wire signed [`CalcTempBus]          temp_m4_32_8_i;
wire signed [`CalcTempBus]          temp_m4_32_9_r;
wire signed [`CalcTempBus]          temp_m4_32_9_i;
wire signed [`CalcTempBus]          temp_m4_32_10_r;
wire signed [`CalcTempBus]          temp_m4_32_10_i;
wire signed [`CalcTempBus]          temp_m4_32_11_r;
wire signed [`CalcTempBus]          temp_m4_32_11_i;
wire signed [`CalcTempBus]          temp_m4_32_12_r;
wire signed [`CalcTempBus]          temp_m4_32_12_i;
wire signed [`CalcTempBus]          temp_m4_32_13_r;
wire signed [`CalcTempBus]          temp_m4_32_13_i;
wire signed [`CalcTempBus]          temp_m4_32_14_r;
wire signed [`CalcTempBus]          temp_m4_32_14_i;
wire signed [`CalcTempBus]          temp_m4_32_15_r;
wire signed [`CalcTempBus]          temp_m4_32_15_i;
wire signed [`CalcTempBus]          temp_m4_32_16_r;
wire signed [`CalcTempBus]          temp_m4_32_16_i;
wire signed [`CalcTempBus]          temp_m4_32_17_r;
wire signed [`CalcTempBus]          temp_m4_32_17_i;
wire signed [`CalcTempBus]          temp_m4_32_18_r;
wire signed [`CalcTempBus]          temp_m4_32_18_i;
wire signed [`CalcTempBus]          temp_m4_32_19_r;
wire signed [`CalcTempBus]          temp_m4_32_19_i;
wire signed [`CalcTempBus]          temp_m4_32_20_r;
wire signed [`CalcTempBus]          temp_m4_32_20_i;
wire signed [`CalcTempBus]          temp_m4_32_21_r;
wire signed [`CalcTempBus]          temp_m4_32_21_i;
wire signed [`CalcTempBus]          temp_m4_32_22_r;
wire signed [`CalcTempBus]          temp_m4_32_22_i;
wire signed [`CalcTempBus]          temp_m4_32_23_r;
wire signed [`CalcTempBus]          temp_m4_32_23_i;
wire signed [`CalcTempBus]          temp_m4_32_24_r;
wire signed [`CalcTempBus]          temp_m4_32_24_i;
wire signed [`CalcTempBus]          temp_m4_32_25_r;
wire signed [`CalcTempBus]          temp_m4_32_25_i;
wire signed [`CalcTempBus]          temp_m4_32_26_r;
wire signed [`CalcTempBus]          temp_m4_32_26_i;
wire signed [`CalcTempBus]          temp_m4_32_27_r;
wire signed [`CalcTempBus]          temp_m4_32_27_i;
wire signed [`CalcTempBus]          temp_m4_32_28_r;
wire signed [`CalcTempBus]          temp_m4_32_28_i;
wire signed [`CalcTempBus]          temp_m4_32_29_r;
wire signed [`CalcTempBus]          temp_m4_32_29_i;
wire signed [`CalcTempBus]          temp_m4_32_30_r;
wire signed [`CalcTempBus]          temp_m4_32_30_i;
wire signed [`CalcTempBus]          temp_m4_32_31_r;
wire signed [`CalcTempBus]          temp_m4_32_31_i;
wire signed [`CalcTempBus]          temp_m4_32_32_r;
wire signed [`CalcTempBus]          temp_m4_32_32_i;
wire signed [`CalcTempBus]          temp_m5_1_1_r;
wire signed [`CalcTempBus]          temp_m5_1_1_i;
wire signed [`CalcTempBus]          temp_m5_1_2_r;
wire signed [`CalcTempBus]          temp_m5_1_2_i;
wire signed [`CalcTempBus]          temp_m5_1_3_r;
wire signed [`CalcTempBus]          temp_m5_1_3_i;
wire signed [`CalcTempBus]          temp_m5_1_4_r;
wire signed [`CalcTempBus]          temp_m5_1_4_i;
wire signed [`CalcTempBus]          temp_m5_1_5_r;
wire signed [`CalcTempBus]          temp_m5_1_5_i;
wire signed [`CalcTempBus]          temp_m5_1_6_r;
wire signed [`CalcTempBus]          temp_m5_1_6_i;
wire signed [`CalcTempBus]          temp_m5_1_7_r;
wire signed [`CalcTempBus]          temp_m5_1_7_i;
wire signed [`CalcTempBus]          temp_m5_1_8_r;
wire signed [`CalcTempBus]          temp_m5_1_8_i;
wire signed [`CalcTempBus]          temp_m5_1_9_r;
wire signed [`CalcTempBus]          temp_m5_1_9_i;
wire signed [`CalcTempBus]          temp_m5_1_10_r;
wire signed [`CalcTempBus]          temp_m5_1_10_i;
wire signed [`CalcTempBus]          temp_m5_1_11_r;
wire signed [`CalcTempBus]          temp_m5_1_11_i;
wire signed [`CalcTempBus]          temp_m5_1_12_r;
wire signed [`CalcTempBus]          temp_m5_1_12_i;
wire signed [`CalcTempBus]          temp_m5_1_13_r;
wire signed [`CalcTempBus]          temp_m5_1_13_i;
wire signed [`CalcTempBus]          temp_m5_1_14_r;
wire signed [`CalcTempBus]          temp_m5_1_14_i;
wire signed [`CalcTempBus]          temp_m5_1_15_r;
wire signed [`CalcTempBus]          temp_m5_1_15_i;
wire signed [`CalcTempBus]          temp_m5_1_16_r;
wire signed [`CalcTempBus]          temp_m5_1_16_i;
wire signed [`CalcTempBus]          temp_m5_1_17_r;
wire signed [`CalcTempBus]          temp_m5_1_17_i;
wire signed [`CalcTempBus]          temp_m5_1_18_r;
wire signed [`CalcTempBus]          temp_m5_1_18_i;
wire signed [`CalcTempBus]          temp_m5_1_19_r;
wire signed [`CalcTempBus]          temp_m5_1_19_i;
wire signed [`CalcTempBus]          temp_m5_1_20_r;
wire signed [`CalcTempBus]          temp_m5_1_20_i;
wire signed [`CalcTempBus]          temp_m5_1_21_r;
wire signed [`CalcTempBus]          temp_m5_1_21_i;
wire signed [`CalcTempBus]          temp_m5_1_22_r;
wire signed [`CalcTempBus]          temp_m5_1_22_i;
wire signed [`CalcTempBus]          temp_m5_1_23_r;
wire signed [`CalcTempBus]          temp_m5_1_23_i;
wire signed [`CalcTempBus]          temp_m5_1_24_r;
wire signed [`CalcTempBus]          temp_m5_1_24_i;
wire signed [`CalcTempBus]          temp_m5_1_25_r;
wire signed [`CalcTempBus]          temp_m5_1_25_i;
wire signed [`CalcTempBus]          temp_m5_1_26_r;
wire signed [`CalcTempBus]          temp_m5_1_26_i;
wire signed [`CalcTempBus]          temp_m5_1_27_r;
wire signed [`CalcTempBus]          temp_m5_1_27_i;
wire signed [`CalcTempBus]          temp_m5_1_28_r;
wire signed [`CalcTempBus]          temp_m5_1_28_i;
wire signed [`CalcTempBus]          temp_m5_1_29_r;
wire signed [`CalcTempBus]          temp_m5_1_29_i;
wire signed [`CalcTempBus]          temp_m5_1_30_r;
wire signed [`CalcTempBus]          temp_m5_1_30_i;
wire signed [`CalcTempBus]          temp_m5_1_31_r;
wire signed [`CalcTempBus]          temp_m5_1_31_i;
wire signed [`CalcTempBus]          temp_m5_1_32_r;
wire signed [`CalcTempBus]          temp_m5_1_32_i;
wire signed [`CalcTempBus]          temp_m5_2_1_r;
wire signed [`CalcTempBus]          temp_m5_2_1_i;
wire signed [`CalcTempBus]          temp_m5_2_2_r;
wire signed [`CalcTempBus]          temp_m5_2_2_i;
wire signed [`CalcTempBus]          temp_m5_2_3_r;
wire signed [`CalcTempBus]          temp_m5_2_3_i;
wire signed [`CalcTempBus]          temp_m5_2_4_r;
wire signed [`CalcTempBus]          temp_m5_2_4_i;
wire signed [`CalcTempBus]          temp_m5_2_5_r;
wire signed [`CalcTempBus]          temp_m5_2_5_i;
wire signed [`CalcTempBus]          temp_m5_2_6_r;
wire signed [`CalcTempBus]          temp_m5_2_6_i;
wire signed [`CalcTempBus]          temp_m5_2_7_r;
wire signed [`CalcTempBus]          temp_m5_2_7_i;
wire signed [`CalcTempBus]          temp_m5_2_8_r;
wire signed [`CalcTempBus]          temp_m5_2_8_i;
wire signed [`CalcTempBus]          temp_m5_2_9_r;
wire signed [`CalcTempBus]          temp_m5_2_9_i;
wire signed [`CalcTempBus]          temp_m5_2_10_r;
wire signed [`CalcTempBus]          temp_m5_2_10_i;
wire signed [`CalcTempBus]          temp_m5_2_11_r;
wire signed [`CalcTempBus]          temp_m5_2_11_i;
wire signed [`CalcTempBus]          temp_m5_2_12_r;
wire signed [`CalcTempBus]          temp_m5_2_12_i;
wire signed [`CalcTempBus]          temp_m5_2_13_r;
wire signed [`CalcTempBus]          temp_m5_2_13_i;
wire signed [`CalcTempBus]          temp_m5_2_14_r;
wire signed [`CalcTempBus]          temp_m5_2_14_i;
wire signed [`CalcTempBus]          temp_m5_2_15_r;
wire signed [`CalcTempBus]          temp_m5_2_15_i;
wire signed [`CalcTempBus]          temp_m5_2_16_r;
wire signed [`CalcTempBus]          temp_m5_2_16_i;
wire signed [`CalcTempBus]          temp_m5_2_17_r;
wire signed [`CalcTempBus]          temp_m5_2_17_i;
wire signed [`CalcTempBus]          temp_m5_2_18_r;
wire signed [`CalcTempBus]          temp_m5_2_18_i;
wire signed [`CalcTempBus]          temp_m5_2_19_r;
wire signed [`CalcTempBus]          temp_m5_2_19_i;
wire signed [`CalcTempBus]          temp_m5_2_20_r;
wire signed [`CalcTempBus]          temp_m5_2_20_i;
wire signed [`CalcTempBus]          temp_m5_2_21_r;
wire signed [`CalcTempBus]          temp_m5_2_21_i;
wire signed [`CalcTempBus]          temp_m5_2_22_r;
wire signed [`CalcTempBus]          temp_m5_2_22_i;
wire signed [`CalcTempBus]          temp_m5_2_23_r;
wire signed [`CalcTempBus]          temp_m5_2_23_i;
wire signed [`CalcTempBus]          temp_m5_2_24_r;
wire signed [`CalcTempBus]          temp_m5_2_24_i;
wire signed [`CalcTempBus]          temp_m5_2_25_r;
wire signed [`CalcTempBus]          temp_m5_2_25_i;
wire signed [`CalcTempBus]          temp_m5_2_26_r;
wire signed [`CalcTempBus]          temp_m5_2_26_i;
wire signed [`CalcTempBus]          temp_m5_2_27_r;
wire signed [`CalcTempBus]          temp_m5_2_27_i;
wire signed [`CalcTempBus]          temp_m5_2_28_r;
wire signed [`CalcTempBus]          temp_m5_2_28_i;
wire signed [`CalcTempBus]          temp_m5_2_29_r;
wire signed [`CalcTempBus]          temp_m5_2_29_i;
wire signed [`CalcTempBus]          temp_m5_2_30_r;
wire signed [`CalcTempBus]          temp_m5_2_30_i;
wire signed [`CalcTempBus]          temp_m5_2_31_r;
wire signed [`CalcTempBus]          temp_m5_2_31_i;
wire signed [`CalcTempBus]          temp_m5_2_32_r;
wire signed [`CalcTempBus]          temp_m5_2_32_i;
wire signed [`CalcTempBus]          temp_m5_3_1_r;
wire signed [`CalcTempBus]          temp_m5_3_1_i;
wire signed [`CalcTempBus]          temp_m5_3_2_r;
wire signed [`CalcTempBus]          temp_m5_3_2_i;
wire signed [`CalcTempBus]          temp_m5_3_3_r;
wire signed [`CalcTempBus]          temp_m5_3_3_i;
wire signed [`CalcTempBus]          temp_m5_3_4_r;
wire signed [`CalcTempBus]          temp_m5_3_4_i;
wire signed [`CalcTempBus]          temp_m5_3_5_r;
wire signed [`CalcTempBus]          temp_m5_3_5_i;
wire signed [`CalcTempBus]          temp_m5_3_6_r;
wire signed [`CalcTempBus]          temp_m5_3_6_i;
wire signed [`CalcTempBus]          temp_m5_3_7_r;
wire signed [`CalcTempBus]          temp_m5_3_7_i;
wire signed [`CalcTempBus]          temp_m5_3_8_r;
wire signed [`CalcTempBus]          temp_m5_3_8_i;
wire signed [`CalcTempBus]          temp_m5_3_9_r;
wire signed [`CalcTempBus]          temp_m5_3_9_i;
wire signed [`CalcTempBus]          temp_m5_3_10_r;
wire signed [`CalcTempBus]          temp_m5_3_10_i;
wire signed [`CalcTempBus]          temp_m5_3_11_r;
wire signed [`CalcTempBus]          temp_m5_3_11_i;
wire signed [`CalcTempBus]          temp_m5_3_12_r;
wire signed [`CalcTempBus]          temp_m5_3_12_i;
wire signed [`CalcTempBus]          temp_m5_3_13_r;
wire signed [`CalcTempBus]          temp_m5_3_13_i;
wire signed [`CalcTempBus]          temp_m5_3_14_r;
wire signed [`CalcTempBus]          temp_m5_3_14_i;
wire signed [`CalcTempBus]          temp_m5_3_15_r;
wire signed [`CalcTempBus]          temp_m5_3_15_i;
wire signed [`CalcTempBus]          temp_m5_3_16_r;
wire signed [`CalcTempBus]          temp_m5_3_16_i;
wire signed [`CalcTempBus]          temp_m5_3_17_r;
wire signed [`CalcTempBus]          temp_m5_3_17_i;
wire signed [`CalcTempBus]          temp_m5_3_18_r;
wire signed [`CalcTempBus]          temp_m5_3_18_i;
wire signed [`CalcTempBus]          temp_m5_3_19_r;
wire signed [`CalcTempBus]          temp_m5_3_19_i;
wire signed [`CalcTempBus]          temp_m5_3_20_r;
wire signed [`CalcTempBus]          temp_m5_3_20_i;
wire signed [`CalcTempBus]          temp_m5_3_21_r;
wire signed [`CalcTempBus]          temp_m5_3_21_i;
wire signed [`CalcTempBus]          temp_m5_3_22_r;
wire signed [`CalcTempBus]          temp_m5_3_22_i;
wire signed [`CalcTempBus]          temp_m5_3_23_r;
wire signed [`CalcTempBus]          temp_m5_3_23_i;
wire signed [`CalcTempBus]          temp_m5_3_24_r;
wire signed [`CalcTempBus]          temp_m5_3_24_i;
wire signed [`CalcTempBus]          temp_m5_3_25_r;
wire signed [`CalcTempBus]          temp_m5_3_25_i;
wire signed [`CalcTempBus]          temp_m5_3_26_r;
wire signed [`CalcTempBus]          temp_m5_3_26_i;
wire signed [`CalcTempBus]          temp_m5_3_27_r;
wire signed [`CalcTempBus]          temp_m5_3_27_i;
wire signed [`CalcTempBus]          temp_m5_3_28_r;
wire signed [`CalcTempBus]          temp_m5_3_28_i;
wire signed [`CalcTempBus]          temp_m5_3_29_r;
wire signed [`CalcTempBus]          temp_m5_3_29_i;
wire signed [`CalcTempBus]          temp_m5_3_30_r;
wire signed [`CalcTempBus]          temp_m5_3_30_i;
wire signed [`CalcTempBus]          temp_m5_3_31_r;
wire signed [`CalcTempBus]          temp_m5_3_31_i;
wire signed [`CalcTempBus]          temp_m5_3_32_r;
wire signed [`CalcTempBus]          temp_m5_3_32_i;
wire signed [`CalcTempBus]          temp_m5_4_1_r;
wire signed [`CalcTempBus]          temp_m5_4_1_i;
wire signed [`CalcTempBus]          temp_m5_4_2_r;
wire signed [`CalcTempBus]          temp_m5_4_2_i;
wire signed [`CalcTempBus]          temp_m5_4_3_r;
wire signed [`CalcTempBus]          temp_m5_4_3_i;
wire signed [`CalcTempBus]          temp_m5_4_4_r;
wire signed [`CalcTempBus]          temp_m5_4_4_i;
wire signed [`CalcTempBus]          temp_m5_4_5_r;
wire signed [`CalcTempBus]          temp_m5_4_5_i;
wire signed [`CalcTempBus]          temp_m5_4_6_r;
wire signed [`CalcTempBus]          temp_m5_4_6_i;
wire signed [`CalcTempBus]          temp_m5_4_7_r;
wire signed [`CalcTempBus]          temp_m5_4_7_i;
wire signed [`CalcTempBus]          temp_m5_4_8_r;
wire signed [`CalcTempBus]          temp_m5_4_8_i;
wire signed [`CalcTempBus]          temp_m5_4_9_r;
wire signed [`CalcTempBus]          temp_m5_4_9_i;
wire signed [`CalcTempBus]          temp_m5_4_10_r;
wire signed [`CalcTempBus]          temp_m5_4_10_i;
wire signed [`CalcTempBus]          temp_m5_4_11_r;
wire signed [`CalcTempBus]          temp_m5_4_11_i;
wire signed [`CalcTempBus]          temp_m5_4_12_r;
wire signed [`CalcTempBus]          temp_m5_4_12_i;
wire signed [`CalcTempBus]          temp_m5_4_13_r;
wire signed [`CalcTempBus]          temp_m5_4_13_i;
wire signed [`CalcTempBus]          temp_m5_4_14_r;
wire signed [`CalcTempBus]          temp_m5_4_14_i;
wire signed [`CalcTempBus]          temp_m5_4_15_r;
wire signed [`CalcTempBus]          temp_m5_4_15_i;
wire signed [`CalcTempBus]          temp_m5_4_16_r;
wire signed [`CalcTempBus]          temp_m5_4_16_i;
wire signed [`CalcTempBus]          temp_m5_4_17_r;
wire signed [`CalcTempBus]          temp_m5_4_17_i;
wire signed [`CalcTempBus]          temp_m5_4_18_r;
wire signed [`CalcTempBus]          temp_m5_4_18_i;
wire signed [`CalcTempBus]          temp_m5_4_19_r;
wire signed [`CalcTempBus]          temp_m5_4_19_i;
wire signed [`CalcTempBus]          temp_m5_4_20_r;
wire signed [`CalcTempBus]          temp_m5_4_20_i;
wire signed [`CalcTempBus]          temp_m5_4_21_r;
wire signed [`CalcTempBus]          temp_m5_4_21_i;
wire signed [`CalcTempBus]          temp_m5_4_22_r;
wire signed [`CalcTempBus]          temp_m5_4_22_i;
wire signed [`CalcTempBus]          temp_m5_4_23_r;
wire signed [`CalcTempBus]          temp_m5_4_23_i;
wire signed [`CalcTempBus]          temp_m5_4_24_r;
wire signed [`CalcTempBus]          temp_m5_4_24_i;
wire signed [`CalcTempBus]          temp_m5_4_25_r;
wire signed [`CalcTempBus]          temp_m5_4_25_i;
wire signed [`CalcTempBus]          temp_m5_4_26_r;
wire signed [`CalcTempBus]          temp_m5_4_26_i;
wire signed [`CalcTempBus]          temp_m5_4_27_r;
wire signed [`CalcTempBus]          temp_m5_4_27_i;
wire signed [`CalcTempBus]          temp_m5_4_28_r;
wire signed [`CalcTempBus]          temp_m5_4_28_i;
wire signed [`CalcTempBus]          temp_m5_4_29_r;
wire signed [`CalcTempBus]          temp_m5_4_29_i;
wire signed [`CalcTempBus]          temp_m5_4_30_r;
wire signed [`CalcTempBus]          temp_m5_4_30_i;
wire signed [`CalcTempBus]          temp_m5_4_31_r;
wire signed [`CalcTempBus]          temp_m5_4_31_i;
wire signed [`CalcTempBus]          temp_m5_4_32_r;
wire signed [`CalcTempBus]          temp_m5_4_32_i;
wire signed [`CalcTempBus]          temp_m5_5_1_r;
wire signed [`CalcTempBus]          temp_m5_5_1_i;
wire signed [`CalcTempBus]          temp_m5_5_2_r;
wire signed [`CalcTempBus]          temp_m5_5_2_i;
wire signed [`CalcTempBus]          temp_m5_5_3_r;
wire signed [`CalcTempBus]          temp_m5_5_3_i;
wire signed [`CalcTempBus]          temp_m5_5_4_r;
wire signed [`CalcTempBus]          temp_m5_5_4_i;
wire signed [`CalcTempBus]          temp_m5_5_5_r;
wire signed [`CalcTempBus]          temp_m5_5_5_i;
wire signed [`CalcTempBus]          temp_m5_5_6_r;
wire signed [`CalcTempBus]          temp_m5_5_6_i;
wire signed [`CalcTempBus]          temp_m5_5_7_r;
wire signed [`CalcTempBus]          temp_m5_5_7_i;
wire signed [`CalcTempBus]          temp_m5_5_8_r;
wire signed [`CalcTempBus]          temp_m5_5_8_i;
wire signed [`CalcTempBus]          temp_m5_5_9_r;
wire signed [`CalcTempBus]          temp_m5_5_9_i;
wire signed [`CalcTempBus]          temp_m5_5_10_r;
wire signed [`CalcTempBus]          temp_m5_5_10_i;
wire signed [`CalcTempBus]          temp_m5_5_11_r;
wire signed [`CalcTempBus]          temp_m5_5_11_i;
wire signed [`CalcTempBus]          temp_m5_5_12_r;
wire signed [`CalcTempBus]          temp_m5_5_12_i;
wire signed [`CalcTempBus]          temp_m5_5_13_r;
wire signed [`CalcTempBus]          temp_m5_5_13_i;
wire signed [`CalcTempBus]          temp_m5_5_14_r;
wire signed [`CalcTempBus]          temp_m5_5_14_i;
wire signed [`CalcTempBus]          temp_m5_5_15_r;
wire signed [`CalcTempBus]          temp_m5_5_15_i;
wire signed [`CalcTempBus]          temp_m5_5_16_r;
wire signed [`CalcTempBus]          temp_m5_5_16_i;
wire signed [`CalcTempBus]          temp_m5_5_17_r;
wire signed [`CalcTempBus]          temp_m5_5_17_i;
wire signed [`CalcTempBus]          temp_m5_5_18_r;
wire signed [`CalcTempBus]          temp_m5_5_18_i;
wire signed [`CalcTempBus]          temp_m5_5_19_r;
wire signed [`CalcTempBus]          temp_m5_5_19_i;
wire signed [`CalcTempBus]          temp_m5_5_20_r;
wire signed [`CalcTempBus]          temp_m5_5_20_i;
wire signed [`CalcTempBus]          temp_m5_5_21_r;
wire signed [`CalcTempBus]          temp_m5_5_21_i;
wire signed [`CalcTempBus]          temp_m5_5_22_r;
wire signed [`CalcTempBus]          temp_m5_5_22_i;
wire signed [`CalcTempBus]          temp_m5_5_23_r;
wire signed [`CalcTempBus]          temp_m5_5_23_i;
wire signed [`CalcTempBus]          temp_m5_5_24_r;
wire signed [`CalcTempBus]          temp_m5_5_24_i;
wire signed [`CalcTempBus]          temp_m5_5_25_r;
wire signed [`CalcTempBus]          temp_m5_5_25_i;
wire signed [`CalcTempBus]          temp_m5_5_26_r;
wire signed [`CalcTempBus]          temp_m5_5_26_i;
wire signed [`CalcTempBus]          temp_m5_5_27_r;
wire signed [`CalcTempBus]          temp_m5_5_27_i;
wire signed [`CalcTempBus]          temp_m5_5_28_r;
wire signed [`CalcTempBus]          temp_m5_5_28_i;
wire signed [`CalcTempBus]          temp_m5_5_29_r;
wire signed [`CalcTempBus]          temp_m5_5_29_i;
wire signed [`CalcTempBus]          temp_m5_5_30_r;
wire signed [`CalcTempBus]          temp_m5_5_30_i;
wire signed [`CalcTempBus]          temp_m5_5_31_r;
wire signed [`CalcTempBus]          temp_m5_5_31_i;
wire signed [`CalcTempBus]          temp_m5_5_32_r;
wire signed [`CalcTempBus]          temp_m5_5_32_i;
wire signed [`CalcTempBus]          temp_m5_6_1_r;
wire signed [`CalcTempBus]          temp_m5_6_1_i;
wire signed [`CalcTempBus]          temp_m5_6_2_r;
wire signed [`CalcTempBus]          temp_m5_6_2_i;
wire signed [`CalcTempBus]          temp_m5_6_3_r;
wire signed [`CalcTempBus]          temp_m5_6_3_i;
wire signed [`CalcTempBus]          temp_m5_6_4_r;
wire signed [`CalcTempBus]          temp_m5_6_4_i;
wire signed [`CalcTempBus]          temp_m5_6_5_r;
wire signed [`CalcTempBus]          temp_m5_6_5_i;
wire signed [`CalcTempBus]          temp_m5_6_6_r;
wire signed [`CalcTempBus]          temp_m5_6_6_i;
wire signed [`CalcTempBus]          temp_m5_6_7_r;
wire signed [`CalcTempBus]          temp_m5_6_7_i;
wire signed [`CalcTempBus]          temp_m5_6_8_r;
wire signed [`CalcTempBus]          temp_m5_6_8_i;
wire signed [`CalcTempBus]          temp_m5_6_9_r;
wire signed [`CalcTempBus]          temp_m5_6_9_i;
wire signed [`CalcTempBus]          temp_m5_6_10_r;
wire signed [`CalcTempBus]          temp_m5_6_10_i;
wire signed [`CalcTempBus]          temp_m5_6_11_r;
wire signed [`CalcTempBus]          temp_m5_6_11_i;
wire signed [`CalcTempBus]          temp_m5_6_12_r;
wire signed [`CalcTempBus]          temp_m5_6_12_i;
wire signed [`CalcTempBus]          temp_m5_6_13_r;
wire signed [`CalcTempBus]          temp_m5_6_13_i;
wire signed [`CalcTempBus]          temp_m5_6_14_r;
wire signed [`CalcTempBus]          temp_m5_6_14_i;
wire signed [`CalcTempBus]          temp_m5_6_15_r;
wire signed [`CalcTempBus]          temp_m5_6_15_i;
wire signed [`CalcTempBus]          temp_m5_6_16_r;
wire signed [`CalcTempBus]          temp_m5_6_16_i;
wire signed [`CalcTempBus]          temp_m5_6_17_r;
wire signed [`CalcTempBus]          temp_m5_6_17_i;
wire signed [`CalcTempBus]          temp_m5_6_18_r;
wire signed [`CalcTempBus]          temp_m5_6_18_i;
wire signed [`CalcTempBus]          temp_m5_6_19_r;
wire signed [`CalcTempBus]          temp_m5_6_19_i;
wire signed [`CalcTempBus]          temp_m5_6_20_r;
wire signed [`CalcTempBus]          temp_m5_6_20_i;
wire signed [`CalcTempBus]          temp_m5_6_21_r;
wire signed [`CalcTempBus]          temp_m5_6_21_i;
wire signed [`CalcTempBus]          temp_m5_6_22_r;
wire signed [`CalcTempBus]          temp_m5_6_22_i;
wire signed [`CalcTempBus]          temp_m5_6_23_r;
wire signed [`CalcTempBus]          temp_m5_6_23_i;
wire signed [`CalcTempBus]          temp_m5_6_24_r;
wire signed [`CalcTempBus]          temp_m5_6_24_i;
wire signed [`CalcTempBus]          temp_m5_6_25_r;
wire signed [`CalcTempBus]          temp_m5_6_25_i;
wire signed [`CalcTempBus]          temp_m5_6_26_r;
wire signed [`CalcTempBus]          temp_m5_6_26_i;
wire signed [`CalcTempBus]          temp_m5_6_27_r;
wire signed [`CalcTempBus]          temp_m5_6_27_i;
wire signed [`CalcTempBus]          temp_m5_6_28_r;
wire signed [`CalcTempBus]          temp_m5_6_28_i;
wire signed [`CalcTempBus]          temp_m5_6_29_r;
wire signed [`CalcTempBus]          temp_m5_6_29_i;
wire signed [`CalcTempBus]          temp_m5_6_30_r;
wire signed [`CalcTempBus]          temp_m5_6_30_i;
wire signed [`CalcTempBus]          temp_m5_6_31_r;
wire signed [`CalcTempBus]          temp_m5_6_31_i;
wire signed [`CalcTempBus]          temp_m5_6_32_r;
wire signed [`CalcTempBus]          temp_m5_6_32_i;
wire signed [`CalcTempBus]          temp_m5_7_1_r;
wire signed [`CalcTempBus]          temp_m5_7_1_i;
wire signed [`CalcTempBus]          temp_m5_7_2_r;
wire signed [`CalcTempBus]          temp_m5_7_2_i;
wire signed [`CalcTempBus]          temp_m5_7_3_r;
wire signed [`CalcTempBus]          temp_m5_7_3_i;
wire signed [`CalcTempBus]          temp_m5_7_4_r;
wire signed [`CalcTempBus]          temp_m5_7_4_i;
wire signed [`CalcTempBus]          temp_m5_7_5_r;
wire signed [`CalcTempBus]          temp_m5_7_5_i;
wire signed [`CalcTempBus]          temp_m5_7_6_r;
wire signed [`CalcTempBus]          temp_m5_7_6_i;
wire signed [`CalcTempBus]          temp_m5_7_7_r;
wire signed [`CalcTempBus]          temp_m5_7_7_i;
wire signed [`CalcTempBus]          temp_m5_7_8_r;
wire signed [`CalcTempBus]          temp_m5_7_8_i;
wire signed [`CalcTempBus]          temp_m5_7_9_r;
wire signed [`CalcTempBus]          temp_m5_7_9_i;
wire signed [`CalcTempBus]          temp_m5_7_10_r;
wire signed [`CalcTempBus]          temp_m5_7_10_i;
wire signed [`CalcTempBus]          temp_m5_7_11_r;
wire signed [`CalcTempBus]          temp_m5_7_11_i;
wire signed [`CalcTempBus]          temp_m5_7_12_r;
wire signed [`CalcTempBus]          temp_m5_7_12_i;
wire signed [`CalcTempBus]          temp_m5_7_13_r;
wire signed [`CalcTempBus]          temp_m5_7_13_i;
wire signed [`CalcTempBus]          temp_m5_7_14_r;
wire signed [`CalcTempBus]          temp_m5_7_14_i;
wire signed [`CalcTempBus]          temp_m5_7_15_r;
wire signed [`CalcTempBus]          temp_m5_7_15_i;
wire signed [`CalcTempBus]          temp_m5_7_16_r;
wire signed [`CalcTempBus]          temp_m5_7_16_i;
wire signed [`CalcTempBus]          temp_m5_7_17_r;
wire signed [`CalcTempBus]          temp_m5_7_17_i;
wire signed [`CalcTempBus]          temp_m5_7_18_r;
wire signed [`CalcTempBus]          temp_m5_7_18_i;
wire signed [`CalcTempBus]          temp_m5_7_19_r;
wire signed [`CalcTempBus]          temp_m5_7_19_i;
wire signed [`CalcTempBus]          temp_m5_7_20_r;
wire signed [`CalcTempBus]          temp_m5_7_20_i;
wire signed [`CalcTempBus]          temp_m5_7_21_r;
wire signed [`CalcTempBus]          temp_m5_7_21_i;
wire signed [`CalcTempBus]          temp_m5_7_22_r;
wire signed [`CalcTempBus]          temp_m5_7_22_i;
wire signed [`CalcTempBus]          temp_m5_7_23_r;
wire signed [`CalcTempBus]          temp_m5_7_23_i;
wire signed [`CalcTempBus]          temp_m5_7_24_r;
wire signed [`CalcTempBus]          temp_m5_7_24_i;
wire signed [`CalcTempBus]          temp_m5_7_25_r;
wire signed [`CalcTempBus]          temp_m5_7_25_i;
wire signed [`CalcTempBus]          temp_m5_7_26_r;
wire signed [`CalcTempBus]          temp_m5_7_26_i;
wire signed [`CalcTempBus]          temp_m5_7_27_r;
wire signed [`CalcTempBus]          temp_m5_7_27_i;
wire signed [`CalcTempBus]          temp_m5_7_28_r;
wire signed [`CalcTempBus]          temp_m5_7_28_i;
wire signed [`CalcTempBus]          temp_m5_7_29_r;
wire signed [`CalcTempBus]          temp_m5_7_29_i;
wire signed [`CalcTempBus]          temp_m5_7_30_r;
wire signed [`CalcTempBus]          temp_m5_7_30_i;
wire signed [`CalcTempBus]          temp_m5_7_31_r;
wire signed [`CalcTempBus]          temp_m5_7_31_i;
wire signed [`CalcTempBus]          temp_m5_7_32_r;
wire signed [`CalcTempBus]          temp_m5_7_32_i;
wire signed [`CalcTempBus]          temp_m5_8_1_r;
wire signed [`CalcTempBus]          temp_m5_8_1_i;
wire signed [`CalcTempBus]          temp_m5_8_2_r;
wire signed [`CalcTempBus]          temp_m5_8_2_i;
wire signed [`CalcTempBus]          temp_m5_8_3_r;
wire signed [`CalcTempBus]          temp_m5_8_3_i;
wire signed [`CalcTempBus]          temp_m5_8_4_r;
wire signed [`CalcTempBus]          temp_m5_8_4_i;
wire signed [`CalcTempBus]          temp_m5_8_5_r;
wire signed [`CalcTempBus]          temp_m5_8_5_i;
wire signed [`CalcTempBus]          temp_m5_8_6_r;
wire signed [`CalcTempBus]          temp_m5_8_6_i;
wire signed [`CalcTempBus]          temp_m5_8_7_r;
wire signed [`CalcTempBus]          temp_m5_8_7_i;
wire signed [`CalcTempBus]          temp_m5_8_8_r;
wire signed [`CalcTempBus]          temp_m5_8_8_i;
wire signed [`CalcTempBus]          temp_m5_8_9_r;
wire signed [`CalcTempBus]          temp_m5_8_9_i;
wire signed [`CalcTempBus]          temp_m5_8_10_r;
wire signed [`CalcTempBus]          temp_m5_8_10_i;
wire signed [`CalcTempBus]          temp_m5_8_11_r;
wire signed [`CalcTempBus]          temp_m5_8_11_i;
wire signed [`CalcTempBus]          temp_m5_8_12_r;
wire signed [`CalcTempBus]          temp_m5_8_12_i;
wire signed [`CalcTempBus]          temp_m5_8_13_r;
wire signed [`CalcTempBus]          temp_m5_8_13_i;
wire signed [`CalcTempBus]          temp_m5_8_14_r;
wire signed [`CalcTempBus]          temp_m5_8_14_i;
wire signed [`CalcTempBus]          temp_m5_8_15_r;
wire signed [`CalcTempBus]          temp_m5_8_15_i;
wire signed [`CalcTempBus]          temp_m5_8_16_r;
wire signed [`CalcTempBus]          temp_m5_8_16_i;
wire signed [`CalcTempBus]          temp_m5_8_17_r;
wire signed [`CalcTempBus]          temp_m5_8_17_i;
wire signed [`CalcTempBus]          temp_m5_8_18_r;
wire signed [`CalcTempBus]          temp_m5_8_18_i;
wire signed [`CalcTempBus]          temp_m5_8_19_r;
wire signed [`CalcTempBus]          temp_m5_8_19_i;
wire signed [`CalcTempBus]          temp_m5_8_20_r;
wire signed [`CalcTempBus]          temp_m5_8_20_i;
wire signed [`CalcTempBus]          temp_m5_8_21_r;
wire signed [`CalcTempBus]          temp_m5_8_21_i;
wire signed [`CalcTempBus]          temp_m5_8_22_r;
wire signed [`CalcTempBus]          temp_m5_8_22_i;
wire signed [`CalcTempBus]          temp_m5_8_23_r;
wire signed [`CalcTempBus]          temp_m5_8_23_i;
wire signed [`CalcTempBus]          temp_m5_8_24_r;
wire signed [`CalcTempBus]          temp_m5_8_24_i;
wire signed [`CalcTempBus]          temp_m5_8_25_r;
wire signed [`CalcTempBus]          temp_m5_8_25_i;
wire signed [`CalcTempBus]          temp_m5_8_26_r;
wire signed [`CalcTempBus]          temp_m5_8_26_i;
wire signed [`CalcTempBus]          temp_m5_8_27_r;
wire signed [`CalcTempBus]          temp_m5_8_27_i;
wire signed [`CalcTempBus]          temp_m5_8_28_r;
wire signed [`CalcTempBus]          temp_m5_8_28_i;
wire signed [`CalcTempBus]          temp_m5_8_29_r;
wire signed [`CalcTempBus]          temp_m5_8_29_i;
wire signed [`CalcTempBus]          temp_m5_8_30_r;
wire signed [`CalcTempBus]          temp_m5_8_30_i;
wire signed [`CalcTempBus]          temp_m5_8_31_r;
wire signed [`CalcTempBus]          temp_m5_8_31_i;
wire signed [`CalcTempBus]          temp_m5_8_32_r;
wire signed [`CalcTempBus]          temp_m5_8_32_i;
wire signed [`CalcTempBus]          temp_m5_9_1_r;
wire signed [`CalcTempBus]          temp_m5_9_1_i;
wire signed [`CalcTempBus]          temp_m5_9_2_r;
wire signed [`CalcTempBus]          temp_m5_9_2_i;
wire signed [`CalcTempBus]          temp_m5_9_3_r;
wire signed [`CalcTempBus]          temp_m5_9_3_i;
wire signed [`CalcTempBus]          temp_m5_9_4_r;
wire signed [`CalcTempBus]          temp_m5_9_4_i;
wire signed [`CalcTempBus]          temp_m5_9_5_r;
wire signed [`CalcTempBus]          temp_m5_9_5_i;
wire signed [`CalcTempBus]          temp_m5_9_6_r;
wire signed [`CalcTempBus]          temp_m5_9_6_i;
wire signed [`CalcTempBus]          temp_m5_9_7_r;
wire signed [`CalcTempBus]          temp_m5_9_7_i;
wire signed [`CalcTempBus]          temp_m5_9_8_r;
wire signed [`CalcTempBus]          temp_m5_9_8_i;
wire signed [`CalcTempBus]          temp_m5_9_9_r;
wire signed [`CalcTempBus]          temp_m5_9_9_i;
wire signed [`CalcTempBus]          temp_m5_9_10_r;
wire signed [`CalcTempBus]          temp_m5_9_10_i;
wire signed [`CalcTempBus]          temp_m5_9_11_r;
wire signed [`CalcTempBus]          temp_m5_9_11_i;
wire signed [`CalcTempBus]          temp_m5_9_12_r;
wire signed [`CalcTempBus]          temp_m5_9_12_i;
wire signed [`CalcTempBus]          temp_m5_9_13_r;
wire signed [`CalcTempBus]          temp_m5_9_13_i;
wire signed [`CalcTempBus]          temp_m5_9_14_r;
wire signed [`CalcTempBus]          temp_m5_9_14_i;
wire signed [`CalcTempBus]          temp_m5_9_15_r;
wire signed [`CalcTempBus]          temp_m5_9_15_i;
wire signed [`CalcTempBus]          temp_m5_9_16_r;
wire signed [`CalcTempBus]          temp_m5_9_16_i;
wire signed [`CalcTempBus]          temp_m5_9_17_r;
wire signed [`CalcTempBus]          temp_m5_9_17_i;
wire signed [`CalcTempBus]          temp_m5_9_18_r;
wire signed [`CalcTempBus]          temp_m5_9_18_i;
wire signed [`CalcTempBus]          temp_m5_9_19_r;
wire signed [`CalcTempBus]          temp_m5_9_19_i;
wire signed [`CalcTempBus]          temp_m5_9_20_r;
wire signed [`CalcTempBus]          temp_m5_9_20_i;
wire signed [`CalcTempBus]          temp_m5_9_21_r;
wire signed [`CalcTempBus]          temp_m5_9_21_i;
wire signed [`CalcTempBus]          temp_m5_9_22_r;
wire signed [`CalcTempBus]          temp_m5_9_22_i;
wire signed [`CalcTempBus]          temp_m5_9_23_r;
wire signed [`CalcTempBus]          temp_m5_9_23_i;
wire signed [`CalcTempBus]          temp_m5_9_24_r;
wire signed [`CalcTempBus]          temp_m5_9_24_i;
wire signed [`CalcTempBus]          temp_m5_9_25_r;
wire signed [`CalcTempBus]          temp_m5_9_25_i;
wire signed [`CalcTempBus]          temp_m5_9_26_r;
wire signed [`CalcTempBus]          temp_m5_9_26_i;
wire signed [`CalcTempBus]          temp_m5_9_27_r;
wire signed [`CalcTempBus]          temp_m5_9_27_i;
wire signed [`CalcTempBus]          temp_m5_9_28_r;
wire signed [`CalcTempBus]          temp_m5_9_28_i;
wire signed [`CalcTempBus]          temp_m5_9_29_r;
wire signed [`CalcTempBus]          temp_m5_9_29_i;
wire signed [`CalcTempBus]          temp_m5_9_30_r;
wire signed [`CalcTempBus]          temp_m5_9_30_i;
wire signed [`CalcTempBus]          temp_m5_9_31_r;
wire signed [`CalcTempBus]          temp_m5_9_31_i;
wire signed [`CalcTempBus]          temp_m5_9_32_r;
wire signed [`CalcTempBus]          temp_m5_9_32_i;
wire signed [`CalcTempBus]          temp_m5_10_1_r;
wire signed [`CalcTempBus]          temp_m5_10_1_i;
wire signed [`CalcTempBus]          temp_m5_10_2_r;
wire signed [`CalcTempBus]          temp_m5_10_2_i;
wire signed [`CalcTempBus]          temp_m5_10_3_r;
wire signed [`CalcTempBus]          temp_m5_10_3_i;
wire signed [`CalcTempBus]          temp_m5_10_4_r;
wire signed [`CalcTempBus]          temp_m5_10_4_i;
wire signed [`CalcTempBus]          temp_m5_10_5_r;
wire signed [`CalcTempBus]          temp_m5_10_5_i;
wire signed [`CalcTempBus]          temp_m5_10_6_r;
wire signed [`CalcTempBus]          temp_m5_10_6_i;
wire signed [`CalcTempBus]          temp_m5_10_7_r;
wire signed [`CalcTempBus]          temp_m5_10_7_i;
wire signed [`CalcTempBus]          temp_m5_10_8_r;
wire signed [`CalcTempBus]          temp_m5_10_8_i;
wire signed [`CalcTempBus]          temp_m5_10_9_r;
wire signed [`CalcTempBus]          temp_m5_10_9_i;
wire signed [`CalcTempBus]          temp_m5_10_10_r;
wire signed [`CalcTempBus]          temp_m5_10_10_i;
wire signed [`CalcTempBus]          temp_m5_10_11_r;
wire signed [`CalcTempBus]          temp_m5_10_11_i;
wire signed [`CalcTempBus]          temp_m5_10_12_r;
wire signed [`CalcTempBus]          temp_m5_10_12_i;
wire signed [`CalcTempBus]          temp_m5_10_13_r;
wire signed [`CalcTempBus]          temp_m5_10_13_i;
wire signed [`CalcTempBus]          temp_m5_10_14_r;
wire signed [`CalcTempBus]          temp_m5_10_14_i;
wire signed [`CalcTempBus]          temp_m5_10_15_r;
wire signed [`CalcTempBus]          temp_m5_10_15_i;
wire signed [`CalcTempBus]          temp_m5_10_16_r;
wire signed [`CalcTempBus]          temp_m5_10_16_i;
wire signed [`CalcTempBus]          temp_m5_10_17_r;
wire signed [`CalcTempBus]          temp_m5_10_17_i;
wire signed [`CalcTempBus]          temp_m5_10_18_r;
wire signed [`CalcTempBus]          temp_m5_10_18_i;
wire signed [`CalcTempBus]          temp_m5_10_19_r;
wire signed [`CalcTempBus]          temp_m5_10_19_i;
wire signed [`CalcTempBus]          temp_m5_10_20_r;
wire signed [`CalcTempBus]          temp_m5_10_20_i;
wire signed [`CalcTempBus]          temp_m5_10_21_r;
wire signed [`CalcTempBus]          temp_m5_10_21_i;
wire signed [`CalcTempBus]          temp_m5_10_22_r;
wire signed [`CalcTempBus]          temp_m5_10_22_i;
wire signed [`CalcTempBus]          temp_m5_10_23_r;
wire signed [`CalcTempBus]          temp_m5_10_23_i;
wire signed [`CalcTempBus]          temp_m5_10_24_r;
wire signed [`CalcTempBus]          temp_m5_10_24_i;
wire signed [`CalcTempBus]          temp_m5_10_25_r;
wire signed [`CalcTempBus]          temp_m5_10_25_i;
wire signed [`CalcTempBus]          temp_m5_10_26_r;
wire signed [`CalcTempBus]          temp_m5_10_26_i;
wire signed [`CalcTempBus]          temp_m5_10_27_r;
wire signed [`CalcTempBus]          temp_m5_10_27_i;
wire signed [`CalcTempBus]          temp_m5_10_28_r;
wire signed [`CalcTempBus]          temp_m5_10_28_i;
wire signed [`CalcTempBus]          temp_m5_10_29_r;
wire signed [`CalcTempBus]          temp_m5_10_29_i;
wire signed [`CalcTempBus]          temp_m5_10_30_r;
wire signed [`CalcTempBus]          temp_m5_10_30_i;
wire signed [`CalcTempBus]          temp_m5_10_31_r;
wire signed [`CalcTempBus]          temp_m5_10_31_i;
wire signed [`CalcTempBus]          temp_m5_10_32_r;
wire signed [`CalcTempBus]          temp_m5_10_32_i;
wire signed [`CalcTempBus]          temp_m5_11_1_r;
wire signed [`CalcTempBus]          temp_m5_11_1_i;
wire signed [`CalcTempBus]          temp_m5_11_2_r;
wire signed [`CalcTempBus]          temp_m5_11_2_i;
wire signed [`CalcTempBus]          temp_m5_11_3_r;
wire signed [`CalcTempBus]          temp_m5_11_3_i;
wire signed [`CalcTempBus]          temp_m5_11_4_r;
wire signed [`CalcTempBus]          temp_m5_11_4_i;
wire signed [`CalcTempBus]          temp_m5_11_5_r;
wire signed [`CalcTempBus]          temp_m5_11_5_i;
wire signed [`CalcTempBus]          temp_m5_11_6_r;
wire signed [`CalcTempBus]          temp_m5_11_6_i;
wire signed [`CalcTempBus]          temp_m5_11_7_r;
wire signed [`CalcTempBus]          temp_m5_11_7_i;
wire signed [`CalcTempBus]          temp_m5_11_8_r;
wire signed [`CalcTempBus]          temp_m5_11_8_i;
wire signed [`CalcTempBus]          temp_m5_11_9_r;
wire signed [`CalcTempBus]          temp_m5_11_9_i;
wire signed [`CalcTempBus]          temp_m5_11_10_r;
wire signed [`CalcTempBus]          temp_m5_11_10_i;
wire signed [`CalcTempBus]          temp_m5_11_11_r;
wire signed [`CalcTempBus]          temp_m5_11_11_i;
wire signed [`CalcTempBus]          temp_m5_11_12_r;
wire signed [`CalcTempBus]          temp_m5_11_12_i;
wire signed [`CalcTempBus]          temp_m5_11_13_r;
wire signed [`CalcTempBus]          temp_m5_11_13_i;
wire signed [`CalcTempBus]          temp_m5_11_14_r;
wire signed [`CalcTempBus]          temp_m5_11_14_i;
wire signed [`CalcTempBus]          temp_m5_11_15_r;
wire signed [`CalcTempBus]          temp_m5_11_15_i;
wire signed [`CalcTempBus]          temp_m5_11_16_r;
wire signed [`CalcTempBus]          temp_m5_11_16_i;
wire signed [`CalcTempBus]          temp_m5_11_17_r;
wire signed [`CalcTempBus]          temp_m5_11_17_i;
wire signed [`CalcTempBus]          temp_m5_11_18_r;
wire signed [`CalcTempBus]          temp_m5_11_18_i;
wire signed [`CalcTempBus]          temp_m5_11_19_r;
wire signed [`CalcTempBus]          temp_m5_11_19_i;
wire signed [`CalcTempBus]          temp_m5_11_20_r;
wire signed [`CalcTempBus]          temp_m5_11_20_i;
wire signed [`CalcTempBus]          temp_m5_11_21_r;
wire signed [`CalcTempBus]          temp_m5_11_21_i;
wire signed [`CalcTempBus]          temp_m5_11_22_r;
wire signed [`CalcTempBus]          temp_m5_11_22_i;
wire signed [`CalcTempBus]          temp_m5_11_23_r;
wire signed [`CalcTempBus]          temp_m5_11_23_i;
wire signed [`CalcTempBus]          temp_m5_11_24_r;
wire signed [`CalcTempBus]          temp_m5_11_24_i;
wire signed [`CalcTempBus]          temp_m5_11_25_r;
wire signed [`CalcTempBus]          temp_m5_11_25_i;
wire signed [`CalcTempBus]          temp_m5_11_26_r;
wire signed [`CalcTempBus]          temp_m5_11_26_i;
wire signed [`CalcTempBus]          temp_m5_11_27_r;
wire signed [`CalcTempBus]          temp_m5_11_27_i;
wire signed [`CalcTempBus]          temp_m5_11_28_r;
wire signed [`CalcTempBus]          temp_m5_11_28_i;
wire signed [`CalcTempBus]          temp_m5_11_29_r;
wire signed [`CalcTempBus]          temp_m5_11_29_i;
wire signed [`CalcTempBus]          temp_m5_11_30_r;
wire signed [`CalcTempBus]          temp_m5_11_30_i;
wire signed [`CalcTempBus]          temp_m5_11_31_r;
wire signed [`CalcTempBus]          temp_m5_11_31_i;
wire signed [`CalcTempBus]          temp_m5_11_32_r;
wire signed [`CalcTempBus]          temp_m5_11_32_i;
wire signed [`CalcTempBus]          temp_m5_12_1_r;
wire signed [`CalcTempBus]          temp_m5_12_1_i;
wire signed [`CalcTempBus]          temp_m5_12_2_r;
wire signed [`CalcTempBus]          temp_m5_12_2_i;
wire signed [`CalcTempBus]          temp_m5_12_3_r;
wire signed [`CalcTempBus]          temp_m5_12_3_i;
wire signed [`CalcTempBus]          temp_m5_12_4_r;
wire signed [`CalcTempBus]          temp_m5_12_4_i;
wire signed [`CalcTempBus]          temp_m5_12_5_r;
wire signed [`CalcTempBus]          temp_m5_12_5_i;
wire signed [`CalcTempBus]          temp_m5_12_6_r;
wire signed [`CalcTempBus]          temp_m5_12_6_i;
wire signed [`CalcTempBus]          temp_m5_12_7_r;
wire signed [`CalcTempBus]          temp_m5_12_7_i;
wire signed [`CalcTempBus]          temp_m5_12_8_r;
wire signed [`CalcTempBus]          temp_m5_12_8_i;
wire signed [`CalcTempBus]          temp_m5_12_9_r;
wire signed [`CalcTempBus]          temp_m5_12_9_i;
wire signed [`CalcTempBus]          temp_m5_12_10_r;
wire signed [`CalcTempBus]          temp_m5_12_10_i;
wire signed [`CalcTempBus]          temp_m5_12_11_r;
wire signed [`CalcTempBus]          temp_m5_12_11_i;
wire signed [`CalcTempBus]          temp_m5_12_12_r;
wire signed [`CalcTempBus]          temp_m5_12_12_i;
wire signed [`CalcTempBus]          temp_m5_12_13_r;
wire signed [`CalcTempBus]          temp_m5_12_13_i;
wire signed [`CalcTempBus]          temp_m5_12_14_r;
wire signed [`CalcTempBus]          temp_m5_12_14_i;
wire signed [`CalcTempBus]          temp_m5_12_15_r;
wire signed [`CalcTempBus]          temp_m5_12_15_i;
wire signed [`CalcTempBus]          temp_m5_12_16_r;
wire signed [`CalcTempBus]          temp_m5_12_16_i;
wire signed [`CalcTempBus]          temp_m5_12_17_r;
wire signed [`CalcTempBus]          temp_m5_12_17_i;
wire signed [`CalcTempBus]          temp_m5_12_18_r;
wire signed [`CalcTempBus]          temp_m5_12_18_i;
wire signed [`CalcTempBus]          temp_m5_12_19_r;
wire signed [`CalcTempBus]          temp_m5_12_19_i;
wire signed [`CalcTempBus]          temp_m5_12_20_r;
wire signed [`CalcTempBus]          temp_m5_12_20_i;
wire signed [`CalcTempBus]          temp_m5_12_21_r;
wire signed [`CalcTempBus]          temp_m5_12_21_i;
wire signed [`CalcTempBus]          temp_m5_12_22_r;
wire signed [`CalcTempBus]          temp_m5_12_22_i;
wire signed [`CalcTempBus]          temp_m5_12_23_r;
wire signed [`CalcTempBus]          temp_m5_12_23_i;
wire signed [`CalcTempBus]          temp_m5_12_24_r;
wire signed [`CalcTempBus]          temp_m5_12_24_i;
wire signed [`CalcTempBus]          temp_m5_12_25_r;
wire signed [`CalcTempBus]          temp_m5_12_25_i;
wire signed [`CalcTempBus]          temp_m5_12_26_r;
wire signed [`CalcTempBus]          temp_m5_12_26_i;
wire signed [`CalcTempBus]          temp_m5_12_27_r;
wire signed [`CalcTempBus]          temp_m5_12_27_i;
wire signed [`CalcTempBus]          temp_m5_12_28_r;
wire signed [`CalcTempBus]          temp_m5_12_28_i;
wire signed [`CalcTempBus]          temp_m5_12_29_r;
wire signed [`CalcTempBus]          temp_m5_12_29_i;
wire signed [`CalcTempBus]          temp_m5_12_30_r;
wire signed [`CalcTempBus]          temp_m5_12_30_i;
wire signed [`CalcTempBus]          temp_m5_12_31_r;
wire signed [`CalcTempBus]          temp_m5_12_31_i;
wire signed [`CalcTempBus]          temp_m5_12_32_r;
wire signed [`CalcTempBus]          temp_m5_12_32_i;
wire signed [`CalcTempBus]          temp_m5_13_1_r;
wire signed [`CalcTempBus]          temp_m5_13_1_i;
wire signed [`CalcTempBus]          temp_m5_13_2_r;
wire signed [`CalcTempBus]          temp_m5_13_2_i;
wire signed [`CalcTempBus]          temp_m5_13_3_r;
wire signed [`CalcTempBus]          temp_m5_13_3_i;
wire signed [`CalcTempBus]          temp_m5_13_4_r;
wire signed [`CalcTempBus]          temp_m5_13_4_i;
wire signed [`CalcTempBus]          temp_m5_13_5_r;
wire signed [`CalcTempBus]          temp_m5_13_5_i;
wire signed [`CalcTempBus]          temp_m5_13_6_r;
wire signed [`CalcTempBus]          temp_m5_13_6_i;
wire signed [`CalcTempBus]          temp_m5_13_7_r;
wire signed [`CalcTempBus]          temp_m5_13_7_i;
wire signed [`CalcTempBus]          temp_m5_13_8_r;
wire signed [`CalcTempBus]          temp_m5_13_8_i;
wire signed [`CalcTempBus]          temp_m5_13_9_r;
wire signed [`CalcTempBus]          temp_m5_13_9_i;
wire signed [`CalcTempBus]          temp_m5_13_10_r;
wire signed [`CalcTempBus]          temp_m5_13_10_i;
wire signed [`CalcTempBus]          temp_m5_13_11_r;
wire signed [`CalcTempBus]          temp_m5_13_11_i;
wire signed [`CalcTempBus]          temp_m5_13_12_r;
wire signed [`CalcTempBus]          temp_m5_13_12_i;
wire signed [`CalcTempBus]          temp_m5_13_13_r;
wire signed [`CalcTempBus]          temp_m5_13_13_i;
wire signed [`CalcTempBus]          temp_m5_13_14_r;
wire signed [`CalcTempBus]          temp_m5_13_14_i;
wire signed [`CalcTempBus]          temp_m5_13_15_r;
wire signed [`CalcTempBus]          temp_m5_13_15_i;
wire signed [`CalcTempBus]          temp_m5_13_16_r;
wire signed [`CalcTempBus]          temp_m5_13_16_i;
wire signed [`CalcTempBus]          temp_m5_13_17_r;
wire signed [`CalcTempBus]          temp_m5_13_17_i;
wire signed [`CalcTempBus]          temp_m5_13_18_r;
wire signed [`CalcTempBus]          temp_m5_13_18_i;
wire signed [`CalcTempBus]          temp_m5_13_19_r;
wire signed [`CalcTempBus]          temp_m5_13_19_i;
wire signed [`CalcTempBus]          temp_m5_13_20_r;
wire signed [`CalcTempBus]          temp_m5_13_20_i;
wire signed [`CalcTempBus]          temp_m5_13_21_r;
wire signed [`CalcTempBus]          temp_m5_13_21_i;
wire signed [`CalcTempBus]          temp_m5_13_22_r;
wire signed [`CalcTempBus]          temp_m5_13_22_i;
wire signed [`CalcTempBus]          temp_m5_13_23_r;
wire signed [`CalcTempBus]          temp_m5_13_23_i;
wire signed [`CalcTempBus]          temp_m5_13_24_r;
wire signed [`CalcTempBus]          temp_m5_13_24_i;
wire signed [`CalcTempBus]          temp_m5_13_25_r;
wire signed [`CalcTempBus]          temp_m5_13_25_i;
wire signed [`CalcTempBus]          temp_m5_13_26_r;
wire signed [`CalcTempBus]          temp_m5_13_26_i;
wire signed [`CalcTempBus]          temp_m5_13_27_r;
wire signed [`CalcTempBus]          temp_m5_13_27_i;
wire signed [`CalcTempBus]          temp_m5_13_28_r;
wire signed [`CalcTempBus]          temp_m5_13_28_i;
wire signed [`CalcTempBus]          temp_m5_13_29_r;
wire signed [`CalcTempBus]          temp_m5_13_29_i;
wire signed [`CalcTempBus]          temp_m5_13_30_r;
wire signed [`CalcTempBus]          temp_m5_13_30_i;
wire signed [`CalcTempBus]          temp_m5_13_31_r;
wire signed [`CalcTempBus]          temp_m5_13_31_i;
wire signed [`CalcTempBus]          temp_m5_13_32_r;
wire signed [`CalcTempBus]          temp_m5_13_32_i;
wire signed [`CalcTempBus]          temp_m5_14_1_r;
wire signed [`CalcTempBus]          temp_m5_14_1_i;
wire signed [`CalcTempBus]          temp_m5_14_2_r;
wire signed [`CalcTempBus]          temp_m5_14_2_i;
wire signed [`CalcTempBus]          temp_m5_14_3_r;
wire signed [`CalcTempBus]          temp_m5_14_3_i;
wire signed [`CalcTempBus]          temp_m5_14_4_r;
wire signed [`CalcTempBus]          temp_m5_14_4_i;
wire signed [`CalcTempBus]          temp_m5_14_5_r;
wire signed [`CalcTempBus]          temp_m5_14_5_i;
wire signed [`CalcTempBus]          temp_m5_14_6_r;
wire signed [`CalcTempBus]          temp_m5_14_6_i;
wire signed [`CalcTempBus]          temp_m5_14_7_r;
wire signed [`CalcTempBus]          temp_m5_14_7_i;
wire signed [`CalcTempBus]          temp_m5_14_8_r;
wire signed [`CalcTempBus]          temp_m5_14_8_i;
wire signed [`CalcTempBus]          temp_m5_14_9_r;
wire signed [`CalcTempBus]          temp_m5_14_9_i;
wire signed [`CalcTempBus]          temp_m5_14_10_r;
wire signed [`CalcTempBus]          temp_m5_14_10_i;
wire signed [`CalcTempBus]          temp_m5_14_11_r;
wire signed [`CalcTempBus]          temp_m5_14_11_i;
wire signed [`CalcTempBus]          temp_m5_14_12_r;
wire signed [`CalcTempBus]          temp_m5_14_12_i;
wire signed [`CalcTempBus]          temp_m5_14_13_r;
wire signed [`CalcTempBus]          temp_m5_14_13_i;
wire signed [`CalcTempBus]          temp_m5_14_14_r;
wire signed [`CalcTempBus]          temp_m5_14_14_i;
wire signed [`CalcTempBus]          temp_m5_14_15_r;
wire signed [`CalcTempBus]          temp_m5_14_15_i;
wire signed [`CalcTempBus]          temp_m5_14_16_r;
wire signed [`CalcTempBus]          temp_m5_14_16_i;
wire signed [`CalcTempBus]          temp_m5_14_17_r;
wire signed [`CalcTempBus]          temp_m5_14_17_i;
wire signed [`CalcTempBus]          temp_m5_14_18_r;
wire signed [`CalcTempBus]          temp_m5_14_18_i;
wire signed [`CalcTempBus]          temp_m5_14_19_r;
wire signed [`CalcTempBus]          temp_m5_14_19_i;
wire signed [`CalcTempBus]          temp_m5_14_20_r;
wire signed [`CalcTempBus]          temp_m5_14_20_i;
wire signed [`CalcTempBus]          temp_m5_14_21_r;
wire signed [`CalcTempBus]          temp_m5_14_21_i;
wire signed [`CalcTempBus]          temp_m5_14_22_r;
wire signed [`CalcTempBus]          temp_m5_14_22_i;
wire signed [`CalcTempBus]          temp_m5_14_23_r;
wire signed [`CalcTempBus]          temp_m5_14_23_i;
wire signed [`CalcTempBus]          temp_m5_14_24_r;
wire signed [`CalcTempBus]          temp_m5_14_24_i;
wire signed [`CalcTempBus]          temp_m5_14_25_r;
wire signed [`CalcTempBus]          temp_m5_14_25_i;
wire signed [`CalcTempBus]          temp_m5_14_26_r;
wire signed [`CalcTempBus]          temp_m5_14_26_i;
wire signed [`CalcTempBus]          temp_m5_14_27_r;
wire signed [`CalcTempBus]          temp_m5_14_27_i;
wire signed [`CalcTempBus]          temp_m5_14_28_r;
wire signed [`CalcTempBus]          temp_m5_14_28_i;
wire signed [`CalcTempBus]          temp_m5_14_29_r;
wire signed [`CalcTempBus]          temp_m5_14_29_i;
wire signed [`CalcTempBus]          temp_m5_14_30_r;
wire signed [`CalcTempBus]          temp_m5_14_30_i;
wire signed [`CalcTempBus]          temp_m5_14_31_r;
wire signed [`CalcTempBus]          temp_m5_14_31_i;
wire signed [`CalcTempBus]          temp_m5_14_32_r;
wire signed [`CalcTempBus]          temp_m5_14_32_i;
wire signed [`CalcTempBus]          temp_m5_15_1_r;
wire signed [`CalcTempBus]          temp_m5_15_1_i;
wire signed [`CalcTempBus]          temp_m5_15_2_r;
wire signed [`CalcTempBus]          temp_m5_15_2_i;
wire signed [`CalcTempBus]          temp_m5_15_3_r;
wire signed [`CalcTempBus]          temp_m5_15_3_i;
wire signed [`CalcTempBus]          temp_m5_15_4_r;
wire signed [`CalcTempBus]          temp_m5_15_4_i;
wire signed [`CalcTempBus]          temp_m5_15_5_r;
wire signed [`CalcTempBus]          temp_m5_15_5_i;
wire signed [`CalcTempBus]          temp_m5_15_6_r;
wire signed [`CalcTempBus]          temp_m5_15_6_i;
wire signed [`CalcTempBus]          temp_m5_15_7_r;
wire signed [`CalcTempBus]          temp_m5_15_7_i;
wire signed [`CalcTempBus]          temp_m5_15_8_r;
wire signed [`CalcTempBus]          temp_m5_15_8_i;
wire signed [`CalcTempBus]          temp_m5_15_9_r;
wire signed [`CalcTempBus]          temp_m5_15_9_i;
wire signed [`CalcTempBus]          temp_m5_15_10_r;
wire signed [`CalcTempBus]          temp_m5_15_10_i;
wire signed [`CalcTempBus]          temp_m5_15_11_r;
wire signed [`CalcTempBus]          temp_m5_15_11_i;
wire signed [`CalcTempBus]          temp_m5_15_12_r;
wire signed [`CalcTempBus]          temp_m5_15_12_i;
wire signed [`CalcTempBus]          temp_m5_15_13_r;
wire signed [`CalcTempBus]          temp_m5_15_13_i;
wire signed [`CalcTempBus]          temp_m5_15_14_r;
wire signed [`CalcTempBus]          temp_m5_15_14_i;
wire signed [`CalcTempBus]          temp_m5_15_15_r;
wire signed [`CalcTempBus]          temp_m5_15_15_i;
wire signed [`CalcTempBus]          temp_m5_15_16_r;
wire signed [`CalcTempBus]          temp_m5_15_16_i;
wire signed [`CalcTempBus]          temp_m5_15_17_r;
wire signed [`CalcTempBus]          temp_m5_15_17_i;
wire signed [`CalcTempBus]          temp_m5_15_18_r;
wire signed [`CalcTempBus]          temp_m5_15_18_i;
wire signed [`CalcTempBus]          temp_m5_15_19_r;
wire signed [`CalcTempBus]          temp_m5_15_19_i;
wire signed [`CalcTempBus]          temp_m5_15_20_r;
wire signed [`CalcTempBus]          temp_m5_15_20_i;
wire signed [`CalcTempBus]          temp_m5_15_21_r;
wire signed [`CalcTempBus]          temp_m5_15_21_i;
wire signed [`CalcTempBus]          temp_m5_15_22_r;
wire signed [`CalcTempBus]          temp_m5_15_22_i;
wire signed [`CalcTempBus]          temp_m5_15_23_r;
wire signed [`CalcTempBus]          temp_m5_15_23_i;
wire signed [`CalcTempBus]          temp_m5_15_24_r;
wire signed [`CalcTempBus]          temp_m5_15_24_i;
wire signed [`CalcTempBus]          temp_m5_15_25_r;
wire signed [`CalcTempBus]          temp_m5_15_25_i;
wire signed [`CalcTempBus]          temp_m5_15_26_r;
wire signed [`CalcTempBus]          temp_m5_15_26_i;
wire signed [`CalcTempBus]          temp_m5_15_27_r;
wire signed [`CalcTempBus]          temp_m5_15_27_i;
wire signed [`CalcTempBus]          temp_m5_15_28_r;
wire signed [`CalcTempBus]          temp_m5_15_28_i;
wire signed [`CalcTempBus]          temp_m5_15_29_r;
wire signed [`CalcTempBus]          temp_m5_15_29_i;
wire signed [`CalcTempBus]          temp_m5_15_30_r;
wire signed [`CalcTempBus]          temp_m5_15_30_i;
wire signed [`CalcTempBus]          temp_m5_15_31_r;
wire signed [`CalcTempBus]          temp_m5_15_31_i;
wire signed [`CalcTempBus]          temp_m5_15_32_r;
wire signed [`CalcTempBus]          temp_m5_15_32_i;
wire signed [`CalcTempBus]          temp_m5_16_1_r;
wire signed [`CalcTempBus]          temp_m5_16_1_i;
wire signed [`CalcTempBus]          temp_m5_16_2_r;
wire signed [`CalcTempBus]          temp_m5_16_2_i;
wire signed [`CalcTempBus]          temp_m5_16_3_r;
wire signed [`CalcTempBus]          temp_m5_16_3_i;
wire signed [`CalcTempBus]          temp_m5_16_4_r;
wire signed [`CalcTempBus]          temp_m5_16_4_i;
wire signed [`CalcTempBus]          temp_m5_16_5_r;
wire signed [`CalcTempBus]          temp_m5_16_5_i;
wire signed [`CalcTempBus]          temp_m5_16_6_r;
wire signed [`CalcTempBus]          temp_m5_16_6_i;
wire signed [`CalcTempBus]          temp_m5_16_7_r;
wire signed [`CalcTempBus]          temp_m5_16_7_i;
wire signed [`CalcTempBus]          temp_m5_16_8_r;
wire signed [`CalcTempBus]          temp_m5_16_8_i;
wire signed [`CalcTempBus]          temp_m5_16_9_r;
wire signed [`CalcTempBus]          temp_m5_16_9_i;
wire signed [`CalcTempBus]          temp_m5_16_10_r;
wire signed [`CalcTempBus]          temp_m5_16_10_i;
wire signed [`CalcTempBus]          temp_m5_16_11_r;
wire signed [`CalcTempBus]          temp_m5_16_11_i;
wire signed [`CalcTempBus]          temp_m5_16_12_r;
wire signed [`CalcTempBus]          temp_m5_16_12_i;
wire signed [`CalcTempBus]          temp_m5_16_13_r;
wire signed [`CalcTempBus]          temp_m5_16_13_i;
wire signed [`CalcTempBus]          temp_m5_16_14_r;
wire signed [`CalcTempBus]          temp_m5_16_14_i;
wire signed [`CalcTempBus]          temp_m5_16_15_r;
wire signed [`CalcTempBus]          temp_m5_16_15_i;
wire signed [`CalcTempBus]          temp_m5_16_16_r;
wire signed [`CalcTempBus]          temp_m5_16_16_i;
wire signed [`CalcTempBus]          temp_m5_16_17_r;
wire signed [`CalcTempBus]          temp_m5_16_17_i;
wire signed [`CalcTempBus]          temp_m5_16_18_r;
wire signed [`CalcTempBus]          temp_m5_16_18_i;
wire signed [`CalcTempBus]          temp_m5_16_19_r;
wire signed [`CalcTempBus]          temp_m5_16_19_i;
wire signed [`CalcTempBus]          temp_m5_16_20_r;
wire signed [`CalcTempBus]          temp_m5_16_20_i;
wire signed [`CalcTempBus]          temp_m5_16_21_r;
wire signed [`CalcTempBus]          temp_m5_16_21_i;
wire signed [`CalcTempBus]          temp_m5_16_22_r;
wire signed [`CalcTempBus]          temp_m5_16_22_i;
wire signed [`CalcTempBus]          temp_m5_16_23_r;
wire signed [`CalcTempBus]          temp_m5_16_23_i;
wire signed [`CalcTempBus]          temp_m5_16_24_r;
wire signed [`CalcTempBus]          temp_m5_16_24_i;
wire signed [`CalcTempBus]          temp_m5_16_25_r;
wire signed [`CalcTempBus]          temp_m5_16_25_i;
wire signed [`CalcTempBus]          temp_m5_16_26_r;
wire signed [`CalcTempBus]          temp_m5_16_26_i;
wire signed [`CalcTempBus]          temp_m5_16_27_r;
wire signed [`CalcTempBus]          temp_m5_16_27_i;
wire signed [`CalcTempBus]          temp_m5_16_28_r;
wire signed [`CalcTempBus]          temp_m5_16_28_i;
wire signed [`CalcTempBus]          temp_m5_16_29_r;
wire signed [`CalcTempBus]          temp_m5_16_29_i;
wire signed [`CalcTempBus]          temp_m5_16_30_r;
wire signed [`CalcTempBus]          temp_m5_16_30_i;
wire signed [`CalcTempBus]          temp_m5_16_31_r;
wire signed [`CalcTempBus]          temp_m5_16_31_i;
wire signed [`CalcTempBus]          temp_m5_16_32_r;
wire signed [`CalcTempBus]          temp_m5_16_32_i;
wire signed [`CalcTempBus]          temp_m5_17_1_r;
wire signed [`CalcTempBus]          temp_m5_17_1_i;
wire signed [`CalcTempBus]          temp_m5_17_2_r;
wire signed [`CalcTempBus]          temp_m5_17_2_i;
wire signed [`CalcTempBus]          temp_m5_17_3_r;
wire signed [`CalcTempBus]          temp_m5_17_3_i;
wire signed [`CalcTempBus]          temp_m5_17_4_r;
wire signed [`CalcTempBus]          temp_m5_17_4_i;
wire signed [`CalcTempBus]          temp_m5_17_5_r;
wire signed [`CalcTempBus]          temp_m5_17_5_i;
wire signed [`CalcTempBus]          temp_m5_17_6_r;
wire signed [`CalcTempBus]          temp_m5_17_6_i;
wire signed [`CalcTempBus]          temp_m5_17_7_r;
wire signed [`CalcTempBus]          temp_m5_17_7_i;
wire signed [`CalcTempBus]          temp_m5_17_8_r;
wire signed [`CalcTempBus]          temp_m5_17_8_i;
wire signed [`CalcTempBus]          temp_m5_17_9_r;
wire signed [`CalcTempBus]          temp_m5_17_9_i;
wire signed [`CalcTempBus]          temp_m5_17_10_r;
wire signed [`CalcTempBus]          temp_m5_17_10_i;
wire signed [`CalcTempBus]          temp_m5_17_11_r;
wire signed [`CalcTempBus]          temp_m5_17_11_i;
wire signed [`CalcTempBus]          temp_m5_17_12_r;
wire signed [`CalcTempBus]          temp_m5_17_12_i;
wire signed [`CalcTempBus]          temp_m5_17_13_r;
wire signed [`CalcTempBus]          temp_m5_17_13_i;
wire signed [`CalcTempBus]          temp_m5_17_14_r;
wire signed [`CalcTempBus]          temp_m5_17_14_i;
wire signed [`CalcTempBus]          temp_m5_17_15_r;
wire signed [`CalcTempBus]          temp_m5_17_15_i;
wire signed [`CalcTempBus]          temp_m5_17_16_r;
wire signed [`CalcTempBus]          temp_m5_17_16_i;
wire signed [`CalcTempBus]          temp_m5_17_17_r;
wire signed [`CalcTempBus]          temp_m5_17_17_i;
wire signed [`CalcTempBus]          temp_m5_17_18_r;
wire signed [`CalcTempBus]          temp_m5_17_18_i;
wire signed [`CalcTempBus]          temp_m5_17_19_r;
wire signed [`CalcTempBus]          temp_m5_17_19_i;
wire signed [`CalcTempBus]          temp_m5_17_20_r;
wire signed [`CalcTempBus]          temp_m5_17_20_i;
wire signed [`CalcTempBus]          temp_m5_17_21_r;
wire signed [`CalcTempBus]          temp_m5_17_21_i;
wire signed [`CalcTempBus]          temp_m5_17_22_r;
wire signed [`CalcTempBus]          temp_m5_17_22_i;
wire signed [`CalcTempBus]          temp_m5_17_23_r;
wire signed [`CalcTempBus]          temp_m5_17_23_i;
wire signed [`CalcTempBus]          temp_m5_17_24_r;
wire signed [`CalcTempBus]          temp_m5_17_24_i;
wire signed [`CalcTempBus]          temp_m5_17_25_r;
wire signed [`CalcTempBus]          temp_m5_17_25_i;
wire signed [`CalcTempBus]          temp_m5_17_26_r;
wire signed [`CalcTempBus]          temp_m5_17_26_i;
wire signed [`CalcTempBus]          temp_m5_17_27_r;
wire signed [`CalcTempBus]          temp_m5_17_27_i;
wire signed [`CalcTempBus]          temp_m5_17_28_r;
wire signed [`CalcTempBus]          temp_m5_17_28_i;
wire signed [`CalcTempBus]          temp_m5_17_29_r;
wire signed [`CalcTempBus]          temp_m5_17_29_i;
wire signed [`CalcTempBus]          temp_m5_17_30_r;
wire signed [`CalcTempBus]          temp_m5_17_30_i;
wire signed [`CalcTempBus]          temp_m5_17_31_r;
wire signed [`CalcTempBus]          temp_m5_17_31_i;
wire signed [`CalcTempBus]          temp_m5_17_32_r;
wire signed [`CalcTempBus]          temp_m5_17_32_i;
wire signed [`CalcTempBus]          temp_m5_18_1_r;
wire signed [`CalcTempBus]          temp_m5_18_1_i;
wire signed [`CalcTempBus]          temp_m5_18_2_r;
wire signed [`CalcTempBus]          temp_m5_18_2_i;
wire signed [`CalcTempBus]          temp_m5_18_3_r;
wire signed [`CalcTempBus]          temp_m5_18_3_i;
wire signed [`CalcTempBus]          temp_m5_18_4_r;
wire signed [`CalcTempBus]          temp_m5_18_4_i;
wire signed [`CalcTempBus]          temp_m5_18_5_r;
wire signed [`CalcTempBus]          temp_m5_18_5_i;
wire signed [`CalcTempBus]          temp_m5_18_6_r;
wire signed [`CalcTempBus]          temp_m5_18_6_i;
wire signed [`CalcTempBus]          temp_m5_18_7_r;
wire signed [`CalcTempBus]          temp_m5_18_7_i;
wire signed [`CalcTempBus]          temp_m5_18_8_r;
wire signed [`CalcTempBus]          temp_m5_18_8_i;
wire signed [`CalcTempBus]          temp_m5_18_9_r;
wire signed [`CalcTempBus]          temp_m5_18_9_i;
wire signed [`CalcTempBus]          temp_m5_18_10_r;
wire signed [`CalcTempBus]          temp_m5_18_10_i;
wire signed [`CalcTempBus]          temp_m5_18_11_r;
wire signed [`CalcTempBus]          temp_m5_18_11_i;
wire signed [`CalcTempBus]          temp_m5_18_12_r;
wire signed [`CalcTempBus]          temp_m5_18_12_i;
wire signed [`CalcTempBus]          temp_m5_18_13_r;
wire signed [`CalcTempBus]          temp_m5_18_13_i;
wire signed [`CalcTempBus]          temp_m5_18_14_r;
wire signed [`CalcTempBus]          temp_m5_18_14_i;
wire signed [`CalcTempBus]          temp_m5_18_15_r;
wire signed [`CalcTempBus]          temp_m5_18_15_i;
wire signed [`CalcTempBus]          temp_m5_18_16_r;
wire signed [`CalcTempBus]          temp_m5_18_16_i;
wire signed [`CalcTempBus]          temp_m5_18_17_r;
wire signed [`CalcTempBus]          temp_m5_18_17_i;
wire signed [`CalcTempBus]          temp_m5_18_18_r;
wire signed [`CalcTempBus]          temp_m5_18_18_i;
wire signed [`CalcTempBus]          temp_m5_18_19_r;
wire signed [`CalcTempBus]          temp_m5_18_19_i;
wire signed [`CalcTempBus]          temp_m5_18_20_r;
wire signed [`CalcTempBus]          temp_m5_18_20_i;
wire signed [`CalcTempBus]          temp_m5_18_21_r;
wire signed [`CalcTempBus]          temp_m5_18_21_i;
wire signed [`CalcTempBus]          temp_m5_18_22_r;
wire signed [`CalcTempBus]          temp_m5_18_22_i;
wire signed [`CalcTempBus]          temp_m5_18_23_r;
wire signed [`CalcTempBus]          temp_m5_18_23_i;
wire signed [`CalcTempBus]          temp_m5_18_24_r;
wire signed [`CalcTempBus]          temp_m5_18_24_i;
wire signed [`CalcTempBus]          temp_m5_18_25_r;
wire signed [`CalcTempBus]          temp_m5_18_25_i;
wire signed [`CalcTempBus]          temp_m5_18_26_r;
wire signed [`CalcTempBus]          temp_m5_18_26_i;
wire signed [`CalcTempBus]          temp_m5_18_27_r;
wire signed [`CalcTempBus]          temp_m5_18_27_i;
wire signed [`CalcTempBus]          temp_m5_18_28_r;
wire signed [`CalcTempBus]          temp_m5_18_28_i;
wire signed [`CalcTempBus]          temp_m5_18_29_r;
wire signed [`CalcTempBus]          temp_m5_18_29_i;
wire signed [`CalcTempBus]          temp_m5_18_30_r;
wire signed [`CalcTempBus]          temp_m5_18_30_i;
wire signed [`CalcTempBus]          temp_m5_18_31_r;
wire signed [`CalcTempBus]          temp_m5_18_31_i;
wire signed [`CalcTempBus]          temp_m5_18_32_r;
wire signed [`CalcTempBus]          temp_m5_18_32_i;
wire signed [`CalcTempBus]          temp_m5_19_1_r;
wire signed [`CalcTempBus]          temp_m5_19_1_i;
wire signed [`CalcTempBus]          temp_m5_19_2_r;
wire signed [`CalcTempBus]          temp_m5_19_2_i;
wire signed [`CalcTempBus]          temp_m5_19_3_r;
wire signed [`CalcTempBus]          temp_m5_19_3_i;
wire signed [`CalcTempBus]          temp_m5_19_4_r;
wire signed [`CalcTempBus]          temp_m5_19_4_i;
wire signed [`CalcTempBus]          temp_m5_19_5_r;
wire signed [`CalcTempBus]          temp_m5_19_5_i;
wire signed [`CalcTempBus]          temp_m5_19_6_r;
wire signed [`CalcTempBus]          temp_m5_19_6_i;
wire signed [`CalcTempBus]          temp_m5_19_7_r;
wire signed [`CalcTempBus]          temp_m5_19_7_i;
wire signed [`CalcTempBus]          temp_m5_19_8_r;
wire signed [`CalcTempBus]          temp_m5_19_8_i;
wire signed [`CalcTempBus]          temp_m5_19_9_r;
wire signed [`CalcTempBus]          temp_m5_19_9_i;
wire signed [`CalcTempBus]          temp_m5_19_10_r;
wire signed [`CalcTempBus]          temp_m5_19_10_i;
wire signed [`CalcTempBus]          temp_m5_19_11_r;
wire signed [`CalcTempBus]          temp_m5_19_11_i;
wire signed [`CalcTempBus]          temp_m5_19_12_r;
wire signed [`CalcTempBus]          temp_m5_19_12_i;
wire signed [`CalcTempBus]          temp_m5_19_13_r;
wire signed [`CalcTempBus]          temp_m5_19_13_i;
wire signed [`CalcTempBus]          temp_m5_19_14_r;
wire signed [`CalcTempBus]          temp_m5_19_14_i;
wire signed [`CalcTempBus]          temp_m5_19_15_r;
wire signed [`CalcTempBus]          temp_m5_19_15_i;
wire signed [`CalcTempBus]          temp_m5_19_16_r;
wire signed [`CalcTempBus]          temp_m5_19_16_i;
wire signed [`CalcTempBus]          temp_m5_19_17_r;
wire signed [`CalcTempBus]          temp_m5_19_17_i;
wire signed [`CalcTempBus]          temp_m5_19_18_r;
wire signed [`CalcTempBus]          temp_m5_19_18_i;
wire signed [`CalcTempBus]          temp_m5_19_19_r;
wire signed [`CalcTempBus]          temp_m5_19_19_i;
wire signed [`CalcTempBus]          temp_m5_19_20_r;
wire signed [`CalcTempBus]          temp_m5_19_20_i;
wire signed [`CalcTempBus]          temp_m5_19_21_r;
wire signed [`CalcTempBus]          temp_m5_19_21_i;
wire signed [`CalcTempBus]          temp_m5_19_22_r;
wire signed [`CalcTempBus]          temp_m5_19_22_i;
wire signed [`CalcTempBus]          temp_m5_19_23_r;
wire signed [`CalcTempBus]          temp_m5_19_23_i;
wire signed [`CalcTempBus]          temp_m5_19_24_r;
wire signed [`CalcTempBus]          temp_m5_19_24_i;
wire signed [`CalcTempBus]          temp_m5_19_25_r;
wire signed [`CalcTempBus]          temp_m5_19_25_i;
wire signed [`CalcTempBus]          temp_m5_19_26_r;
wire signed [`CalcTempBus]          temp_m5_19_26_i;
wire signed [`CalcTempBus]          temp_m5_19_27_r;
wire signed [`CalcTempBus]          temp_m5_19_27_i;
wire signed [`CalcTempBus]          temp_m5_19_28_r;
wire signed [`CalcTempBus]          temp_m5_19_28_i;
wire signed [`CalcTempBus]          temp_m5_19_29_r;
wire signed [`CalcTempBus]          temp_m5_19_29_i;
wire signed [`CalcTempBus]          temp_m5_19_30_r;
wire signed [`CalcTempBus]          temp_m5_19_30_i;
wire signed [`CalcTempBus]          temp_m5_19_31_r;
wire signed [`CalcTempBus]          temp_m5_19_31_i;
wire signed [`CalcTempBus]          temp_m5_19_32_r;
wire signed [`CalcTempBus]          temp_m5_19_32_i;
wire signed [`CalcTempBus]          temp_m5_20_1_r;
wire signed [`CalcTempBus]          temp_m5_20_1_i;
wire signed [`CalcTempBus]          temp_m5_20_2_r;
wire signed [`CalcTempBus]          temp_m5_20_2_i;
wire signed [`CalcTempBus]          temp_m5_20_3_r;
wire signed [`CalcTempBus]          temp_m5_20_3_i;
wire signed [`CalcTempBus]          temp_m5_20_4_r;
wire signed [`CalcTempBus]          temp_m5_20_4_i;
wire signed [`CalcTempBus]          temp_m5_20_5_r;
wire signed [`CalcTempBus]          temp_m5_20_5_i;
wire signed [`CalcTempBus]          temp_m5_20_6_r;
wire signed [`CalcTempBus]          temp_m5_20_6_i;
wire signed [`CalcTempBus]          temp_m5_20_7_r;
wire signed [`CalcTempBus]          temp_m5_20_7_i;
wire signed [`CalcTempBus]          temp_m5_20_8_r;
wire signed [`CalcTempBus]          temp_m5_20_8_i;
wire signed [`CalcTempBus]          temp_m5_20_9_r;
wire signed [`CalcTempBus]          temp_m5_20_9_i;
wire signed [`CalcTempBus]          temp_m5_20_10_r;
wire signed [`CalcTempBus]          temp_m5_20_10_i;
wire signed [`CalcTempBus]          temp_m5_20_11_r;
wire signed [`CalcTempBus]          temp_m5_20_11_i;
wire signed [`CalcTempBus]          temp_m5_20_12_r;
wire signed [`CalcTempBus]          temp_m5_20_12_i;
wire signed [`CalcTempBus]          temp_m5_20_13_r;
wire signed [`CalcTempBus]          temp_m5_20_13_i;
wire signed [`CalcTempBus]          temp_m5_20_14_r;
wire signed [`CalcTempBus]          temp_m5_20_14_i;
wire signed [`CalcTempBus]          temp_m5_20_15_r;
wire signed [`CalcTempBus]          temp_m5_20_15_i;
wire signed [`CalcTempBus]          temp_m5_20_16_r;
wire signed [`CalcTempBus]          temp_m5_20_16_i;
wire signed [`CalcTempBus]          temp_m5_20_17_r;
wire signed [`CalcTempBus]          temp_m5_20_17_i;
wire signed [`CalcTempBus]          temp_m5_20_18_r;
wire signed [`CalcTempBus]          temp_m5_20_18_i;
wire signed [`CalcTempBus]          temp_m5_20_19_r;
wire signed [`CalcTempBus]          temp_m5_20_19_i;
wire signed [`CalcTempBus]          temp_m5_20_20_r;
wire signed [`CalcTempBus]          temp_m5_20_20_i;
wire signed [`CalcTempBus]          temp_m5_20_21_r;
wire signed [`CalcTempBus]          temp_m5_20_21_i;
wire signed [`CalcTempBus]          temp_m5_20_22_r;
wire signed [`CalcTempBus]          temp_m5_20_22_i;
wire signed [`CalcTempBus]          temp_m5_20_23_r;
wire signed [`CalcTempBus]          temp_m5_20_23_i;
wire signed [`CalcTempBus]          temp_m5_20_24_r;
wire signed [`CalcTempBus]          temp_m5_20_24_i;
wire signed [`CalcTempBus]          temp_m5_20_25_r;
wire signed [`CalcTempBus]          temp_m5_20_25_i;
wire signed [`CalcTempBus]          temp_m5_20_26_r;
wire signed [`CalcTempBus]          temp_m5_20_26_i;
wire signed [`CalcTempBus]          temp_m5_20_27_r;
wire signed [`CalcTempBus]          temp_m5_20_27_i;
wire signed [`CalcTempBus]          temp_m5_20_28_r;
wire signed [`CalcTempBus]          temp_m5_20_28_i;
wire signed [`CalcTempBus]          temp_m5_20_29_r;
wire signed [`CalcTempBus]          temp_m5_20_29_i;
wire signed [`CalcTempBus]          temp_m5_20_30_r;
wire signed [`CalcTempBus]          temp_m5_20_30_i;
wire signed [`CalcTempBus]          temp_m5_20_31_r;
wire signed [`CalcTempBus]          temp_m5_20_31_i;
wire signed [`CalcTempBus]          temp_m5_20_32_r;
wire signed [`CalcTempBus]          temp_m5_20_32_i;
wire signed [`CalcTempBus]          temp_m5_21_1_r;
wire signed [`CalcTempBus]          temp_m5_21_1_i;
wire signed [`CalcTempBus]          temp_m5_21_2_r;
wire signed [`CalcTempBus]          temp_m5_21_2_i;
wire signed [`CalcTempBus]          temp_m5_21_3_r;
wire signed [`CalcTempBus]          temp_m5_21_3_i;
wire signed [`CalcTempBus]          temp_m5_21_4_r;
wire signed [`CalcTempBus]          temp_m5_21_4_i;
wire signed [`CalcTempBus]          temp_m5_21_5_r;
wire signed [`CalcTempBus]          temp_m5_21_5_i;
wire signed [`CalcTempBus]          temp_m5_21_6_r;
wire signed [`CalcTempBus]          temp_m5_21_6_i;
wire signed [`CalcTempBus]          temp_m5_21_7_r;
wire signed [`CalcTempBus]          temp_m5_21_7_i;
wire signed [`CalcTempBus]          temp_m5_21_8_r;
wire signed [`CalcTempBus]          temp_m5_21_8_i;
wire signed [`CalcTempBus]          temp_m5_21_9_r;
wire signed [`CalcTempBus]          temp_m5_21_9_i;
wire signed [`CalcTempBus]          temp_m5_21_10_r;
wire signed [`CalcTempBus]          temp_m5_21_10_i;
wire signed [`CalcTempBus]          temp_m5_21_11_r;
wire signed [`CalcTempBus]          temp_m5_21_11_i;
wire signed [`CalcTempBus]          temp_m5_21_12_r;
wire signed [`CalcTempBus]          temp_m5_21_12_i;
wire signed [`CalcTempBus]          temp_m5_21_13_r;
wire signed [`CalcTempBus]          temp_m5_21_13_i;
wire signed [`CalcTempBus]          temp_m5_21_14_r;
wire signed [`CalcTempBus]          temp_m5_21_14_i;
wire signed [`CalcTempBus]          temp_m5_21_15_r;
wire signed [`CalcTempBus]          temp_m5_21_15_i;
wire signed [`CalcTempBus]          temp_m5_21_16_r;
wire signed [`CalcTempBus]          temp_m5_21_16_i;
wire signed [`CalcTempBus]          temp_m5_21_17_r;
wire signed [`CalcTempBus]          temp_m5_21_17_i;
wire signed [`CalcTempBus]          temp_m5_21_18_r;
wire signed [`CalcTempBus]          temp_m5_21_18_i;
wire signed [`CalcTempBus]          temp_m5_21_19_r;
wire signed [`CalcTempBus]          temp_m5_21_19_i;
wire signed [`CalcTempBus]          temp_m5_21_20_r;
wire signed [`CalcTempBus]          temp_m5_21_20_i;
wire signed [`CalcTempBus]          temp_m5_21_21_r;
wire signed [`CalcTempBus]          temp_m5_21_21_i;
wire signed [`CalcTempBus]          temp_m5_21_22_r;
wire signed [`CalcTempBus]          temp_m5_21_22_i;
wire signed [`CalcTempBus]          temp_m5_21_23_r;
wire signed [`CalcTempBus]          temp_m5_21_23_i;
wire signed [`CalcTempBus]          temp_m5_21_24_r;
wire signed [`CalcTempBus]          temp_m5_21_24_i;
wire signed [`CalcTempBus]          temp_m5_21_25_r;
wire signed [`CalcTempBus]          temp_m5_21_25_i;
wire signed [`CalcTempBus]          temp_m5_21_26_r;
wire signed [`CalcTempBus]          temp_m5_21_26_i;
wire signed [`CalcTempBus]          temp_m5_21_27_r;
wire signed [`CalcTempBus]          temp_m5_21_27_i;
wire signed [`CalcTempBus]          temp_m5_21_28_r;
wire signed [`CalcTempBus]          temp_m5_21_28_i;
wire signed [`CalcTempBus]          temp_m5_21_29_r;
wire signed [`CalcTempBus]          temp_m5_21_29_i;
wire signed [`CalcTempBus]          temp_m5_21_30_r;
wire signed [`CalcTempBus]          temp_m5_21_30_i;
wire signed [`CalcTempBus]          temp_m5_21_31_r;
wire signed [`CalcTempBus]          temp_m5_21_31_i;
wire signed [`CalcTempBus]          temp_m5_21_32_r;
wire signed [`CalcTempBus]          temp_m5_21_32_i;
wire signed [`CalcTempBus]          temp_m5_22_1_r;
wire signed [`CalcTempBus]          temp_m5_22_1_i;
wire signed [`CalcTempBus]          temp_m5_22_2_r;
wire signed [`CalcTempBus]          temp_m5_22_2_i;
wire signed [`CalcTempBus]          temp_m5_22_3_r;
wire signed [`CalcTempBus]          temp_m5_22_3_i;
wire signed [`CalcTempBus]          temp_m5_22_4_r;
wire signed [`CalcTempBus]          temp_m5_22_4_i;
wire signed [`CalcTempBus]          temp_m5_22_5_r;
wire signed [`CalcTempBus]          temp_m5_22_5_i;
wire signed [`CalcTempBus]          temp_m5_22_6_r;
wire signed [`CalcTempBus]          temp_m5_22_6_i;
wire signed [`CalcTempBus]          temp_m5_22_7_r;
wire signed [`CalcTempBus]          temp_m5_22_7_i;
wire signed [`CalcTempBus]          temp_m5_22_8_r;
wire signed [`CalcTempBus]          temp_m5_22_8_i;
wire signed [`CalcTempBus]          temp_m5_22_9_r;
wire signed [`CalcTempBus]          temp_m5_22_9_i;
wire signed [`CalcTempBus]          temp_m5_22_10_r;
wire signed [`CalcTempBus]          temp_m5_22_10_i;
wire signed [`CalcTempBus]          temp_m5_22_11_r;
wire signed [`CalcTempBus]          temp_m5_22_11_i;
wire signed [`CalcTempBus]          temp_m5_22_12_r;
wire signed [`CalcTempBus]          temp_m5_22_12_i;
wire signed [`CalcTempBus]          temp_m5_22_13_r;
wire signed [`CalcTempBus]          temp_m5_22_13_i;
wire signed [`CalcTempBus]          temp_m5_22_14_r;
wire signed [`CalcTempBus]          temp_m5_22_14_i;
wire signed [`CalcTempBus]          temp_m5_22_15_r;
wire signed [`CalcTempBus]          temp_m5_22_15_i;
wire signed [`CalcTempBus]          temp_m5_22_16_r;
wire signed [`CalcTempBus]          temp_m5_22_16_i;
wire signed [`CalcTempBus]          temp_m5_22_17_r;
wire signed [`CalcTempBus]          temp_m5_22_17_i;
wire signed [`CalcTempBus]          temp_m5_22_18_r;
wire signed [`CalcTempBus]          temp_m5_22_18_i;
wire signed [`CalcTempBus]          temp_m5_22_19_r;
wire signed [`CalcTempBus]          temp_m5_22_19_i;
wire signed [`CalcTempBus]          temp_m5_22_20_r;
wire signed [`CalcTempBus]          temp_m5_22_20_i;
wire signed [`CalcTempBus]          temp_m5_22_21_r;
wire signed [`CalcTempBus]          temp_m5_22_21_i;
wire signed [`CalcTempBus]          temp_m5_22_22_r;
wire signed [`CalcTempBus]          temp_m5_22_22_i;
wire signed [`CalcTempBus]          temp_m5_22_23_r;
wire signed [`CalcTempBus]          temp_m5_22_23_i;
wire signed [`CalcTempBus]          temp_m5_22_24_r;
wire signed [`CalcTempBus]          temp_m5_22_24_i;
wire signed [`CalcTempBus]          temp_m5_22_25_r;
wire signed [`CalcTempBus]          temp_m5_22_25_i;
wire signed [`CalcTempBus]          temp_m5_22_26_r;
wire signed [`CalcTempBus]          temp_m5_22_26_i;
wire signed [`CalcTempBus]          temp_m5_22_27_r;
wire signed [`CalcTempBus]          temp_m5_22_27_i;
wire signed [`CalcTempBus]          temp_m5_22_28_r;
wire signed [`CalcTempBus]          temp_m5_22_28_i;
wire signed [`CalcTempBus]          temp_m5_22_29_r;
wire signed [`CalcTempBus]          temp_m5_22_29_i;
wire signed [`CalcTempBus]          temp_m5_22_30_r;
wire signed [`CalcTempBus]          temp_m5_22_30_i;
wire signed [`CalcTempBus]          temp_m5_22_31_r;
wire signed [`CalcTempBus]          temp_m5_22_31_i;
wire signed [`CalcTempBus]          temp_m5_22_32_r;
wire signed [`CalcTempBus]          temp_m5_22_32_i;
wire signed [`CalcTempBus]          temp_m5_23_1_r;
wire signed [`CalcTempBus]          temp_m5_23_1_i;
wire signed [`CalcTempBus]          temp_m5_23_2_r;
wire signed [`CalcTempBus]          temp_m5_23_2_i;
wire signed [`CalcTempBus]          temp_m5_23_3_r;
wire signed [`CalcTempBus]          temp_m5_23_3_i;
wire signed [`CalcTempBus]          temp_m5_23_4_r;
wire signed [`CalcTempBus]          temp_m5_23_4_i;
wire signed [`CalcTempBus]          temp_m5_23_5_r;
wire signed [`CalcTempBus]          temp_m5_23_5_i;
wire signed [`CalcTempBus]          temp_m5_23_6_r;
wire signed [`CalcTempBus]          temp_m5_23_6_i;
wire signed [`CalcTempBus]          temp_m5_23_7_r;
wire signed [`CalcTempBus]          temp_m5_23_7_i;
wire signed [`CalcTempBus]          temp_m5_23_8_r;
wire signed [`CalcTempBus]          temp_m5_23_8_i;
wire signed [`CalcTempBus]          temp_m5_23_9_r;
wire signed [`CalcTempBus]          temp_m5_23_9_i;
wire signed [`CalcTempBus]          temp_m5_23_10_r;
wire signed [`CalcTempBus]          temp_m5_23_10_i;
wire signed [`CalcTempBus]          temp_m5_23_11_r;
wire signed [`CalcTempBus]          temp_m5_23_11_i;
wire signed [`CalcTempBus]          temp_m5_23_12_r;
wire signed [`CalcTempBus]          temp_m5_23_12_i;
wire signed [`CalcTempBus]          temp_m5_23_13_r;
wire signed [`CalcTempBus]          temp_m5_23_13_i;
wire signed [`CalcTempBus]          temp_m5_23_14_r;
wire signed [`CalcTempBus]          temp_m5_23_14_i;
wire signed [`CalcTempBus]          temp_m5_23_15_r;
wire signed [`CalcTempBus]          temp_m5_23_15_i;
wire signed [`CalcTempBus]          temp_m5_23_16_r;
wire signed [`CalcTempBus]          temp_m5_23_16_i;
wire signed [`CalcTempBus]          temp_m5_23_17_r;
wire signed [`CalcTempBus]          temp_m5_23_17_i;
wire signed [`CalcTempBus]          temp_m5_23_18_r;
wire signed [`CalcTempBus]          temp_m5_23_18_i;
wire signed [`CalcTempBus]          temp_m5_23_19_r;
wire signed [`CalcTempBus]          temp_m5_23_19_i;
wire signed [`CalcTempBus]          temp_m5_23_20_r;
wire signed [`CalcTempBus]          temp_m5_23_20_i;
wire signed [`CalcTempBus]          temp_m5_23_21_r;
wire signed [`CalcTempBus]          temp_m5_23_21_i;
wire signed [`CalcTempBus]          temp_m5_23_22_r;
wire signed [`CalcTempBus]          temp_m5_23_22_i;
wire signed [`CalcTempBus]          temp_m5_23_23_r;
wire signed [`CalcTempBus]          temp_m5_23_23_i;
wire signed [`CalcTempBus]          temp_m5_23_24_r;
wire signed [`CalcTempBus]          temp_m5_23_24_i;
wire signed [`CalcTempBus]          temp_m5_23_25_r;
wire signed [`CalcTempBus]          temp_m5_23_25_i;
wire signed [`CalcTempBus]          temp_m5_23_26_r;
wire signed [`CalcTempBus]          temp_m5_23_26_i;
wire signed [`CalcTempBus]          temp_m5_23_27_r;
wire signed [`CalcTempBus]          temp_m5_23_27_i;
wire signed [`CalcTempBus]          temp_m5_23_28_r;
wire signed [`CalcTempBus]          temp_m5_23_28_i;
wire signed [`CalcTempBus]          temp_m5_23_29_r;
wire signed [`CalcTempBus]          temp_m5_23_29_i;
wire signed [`CalcTempBus]          temp_m5_23_30_r;
wire signed [`CalcTempBus]          temp_m5_23_30_i;
wire signed [`CalcTempBus]          temp_m5_23_31_r;
wire signed [`CalcTempBus]          temp_m5_23_31_i;
wire signed [`CalcTempBus]          temp_m5_23_32_r;
wire signed [`CalcTempBus]          temp_m5_23_32_i;
wire signed [`CalcTempBus]          temp_m5_24_1_r;
wire signed [`CalcTempBus]          temp_m5_24_1_i;
wire signed [`CalcTempBus]          temp_m5_24_2_r;
wire signed [`CalcTempBus]          temp_m5_24_2_i;
wire signed [`CalcTempBus]          temp_m5_24_3_r;
wire signed [`CalcTempBus]          temp_m5_24_3_i;
wire signed [`CalcTempBus]          temp_m5_24_4_r;
wire signed [`CalcTempBus]          temp_m5_24_4_i;
wire signed [`CalcTempBus]          temp_m5_24_5_r;
wire signed [`CalcTempBus]          temp_m5_24_5_i;
wire signed [`CalcTempBus]          temp_m5_24_6_r;
wire signed [`CalcTempBus]          temp_m5_24_6_i;
wire signed [`CalcTempBus]          temp_m5_24_7_r;
wire signed [`CalcTempBus]          temp_m5_24_7_i;
wire signed [`CalcTempBus]          temp_m5_24_8_r;
wire signed [`CalcTempBus]          temp_m5_24_8_i;
wire signed [`CalcTempBus]          temp_m5_24_9_r;
wire signed [`CalcTempBus]          temp_m5_24_9_i;
wire signed [`CalcTempBus]          temp_m5_24_10_r;
wire signed [`CalcTempBus]          temp_m5_24_10_i;
wire signed [`CalcTempBus]          temp_m5_24_11_r;
wire signed [`CalcTempBus]          temp_m5_24_11_i;
wire signed [`CalcTempBus]          temp_m5_24_12_r;
wire signed [`CalcTempBus]          temp_m5_24_12_i;
wire signed [`CalcTempBus]          temp_m5_24_13_r;
wire signed [`CalcTempBus]          temp_m5_24_13_i;
wire signed [`CalcTempBus]          temp_m5_24_14_r;
wire signed [`CalcTempBus]          temp_m5_24_14_i;
wire signed [`CalcTempBus]          temp_m5_24_15_r;
wire signed [`CalcTempBus]          temp_m5_24_15_i;
wire signed [`CalcTempBus]          temp_m5_24_16_r;
wire signed [`CalcTempBus]          temp_m5_24_16_i;
wire signed [`CalcTempBus]          temp_m5_24_17_r;
wire signed [`CalcTempBus]          temp_m5_24_17_i;
wire signed [`CalcTempBus]          temp_m5_24_18_r;
wire signed [`CalcTempBus]          temp_m5_24_18_i;
wire signed [`CalcTempBus]          temp_m5_24_19_r;
wire signed [`CalcTempBus]          temp_m5_24_19_i;
wire signed [`CalcTempBus]          temp_m5_24_20_r;
wire signed [`CalcTempBus]          temp_m5_24_20_i;
wire signed [`CalcTempBus]          temp_m5_24_21_r;
wire signed [`CalcTempBus]          temp_m5_24_21_i;
wire signed [`CalcTempBus]          temp_m5_24_22_r;
wire signed [`CalcTempBus]          temp_m5_24_22_i;
wire signed [`CalcTempBus]          temp_m5_24_23_r;
wire signed [`CalcTempBus]          temp_m5_24_23_i;
wire signed [`CalcTempBus]          temp_m5_24_24_r;
wire signed [`CalcTempBus]          temp_m5_24_24_i;
wire signed [`CalcTempBus]          temp_m5_24_25_r;
wire signed [`CalcTempBus]          temp_m5_24_25_i;
wire signed [`CalcTempBus]          temp_m5_24_26_r;
wire signed [`CalcTempBus]          temp_m5_24_26_i;
wire signed [`CalcTempBus]          temp_m5_24_27_r;
wire signed [`CalcTempBus]          temp_m5_24_27_i;
wire signed [`CalcTempBus]          temp_m5_24_28_r;
wire signed [`CalcTempBus]          temp_m5_24_28_i;
wire signed [`CalcTempBus]          temp_m5_24_29_r;
wire signed [`CalcTempBus]          temp_m5_24_29_i;
wire signed [`CalcTempBus]          temp_m5_24_30_r;
wire signed [`CalcTempBus]          temp_m5_24_30_i;
wire signed [`CalcTempBus]          temp_m5_24_31_r;
wire signed [`CalcTempBus]          temp_m5_24_31_i;
wire signed [`CalcTempBus]          temp_m5_24_32_r;
wire signed [`CalcTempBus]          temp_m5_24_32_i;
wire signed [`CalcTempBus]          temp_m5_25_1_r;
wire signed [`CalcTempBus]          temp_m5_25_1_i;
wire signed [`CalcTempBus]          temp_m5_25_2_r;
wire signed [`CalcTempBus]          temp_m5_25_2_i;
wire signed [`CalcTempBus]          temp_m5_25_3_r;
wire signed [`CalcTempBus]          temp_m5_25_3_i;
wire signed [`CalcTempBus]          temp_m5_25_4_r;
wire signed [`CalcTempBus]          temp_m5_25_4_i;
wire signed [`CalcTempBus]          temp_m5_25_5_r;
wire signed [`CalcTempBus]          temp_m5_25_5_i;
wire signed [`CalcTempBus]          temp_m5_25_6_r;
wire signed [`CalcTempBus]          temp_m5_25_6_i;
wire signed [`CalcTempBus]          temp_m5_25_7_r;
wire signed [`CalcTempBus]          temp_m5_25_7_i;
wire signed [`CalcTempBus]          temp_m5_25_8_r;
wire signed [`CalcTempBus]          temp_m5_25_8_i;
wire signed [`CalcTempBus]          temp_m5_25_9_r;
wire signed [`CalcTempBus]          temp_m5_25_9_i;
wire signed [`CalcTempBus]          temp_m5_25_10_r;
wire signed [`CalcTempBus]          temp_m5_25_10_i;
wire signed [`CalcTempBus]          temp_m5_25_11_r;
wire signed [`CalcTempBus]          temp_m5_25_11_i;
wire signed [`CalcTempBus]          temp_m5_25_12_r;
wire signed [`CalcTempBus]          temp_m5_25_12_i;
wire signed [`CalcTempBus]          temp_m5_25_13_r;
wire signed [`CalcTempBus]          temp_m5_25_13_i;
wire signed [`CalcTempBus]          temp_m5_25_14_r;
wire signed [`CalcTempBus]          temp_m5_25_14_i;
wire signed [`CalcTempBus]          temp_m5_25_15_r;
wire signed [`CalcTempBus]          temp_m5_25_15_i;
wire signed [`CalcTempBus]          temp_m5_25_16_r;
wire signed [`CalcTempBus]          temp_m5_25_16_i;
wire signed [`CalcTempBus]          temp_m5_25_17_r;
wire signed [`CalcTempBus]          temp_m5_25_17_i;
wire signed [`CalcTempBus]          temp_m5_25_18_r;
wire signed [`CalcTempBus]          temp_m5_25_18_i;
wire signed [`CalcTempBus]          temp_m5_25_19_r;
wire signed [`CalcTempBus]          temp_m5_25_19_i;
wire signed [`CalcTempBus]          temp_m5_25_20_r;
wire signed [`CalcTempBus]          temp_m5_25_20_i;
wire signed [`CalcTempBus]          temp_m5_25_21_r;
wire signed [`CalcTempBus]          temp_m5_25_21_i;
wire signed [`CalcTempBus]          temp_m5_25_22_r;
wire signed [`CalcTempBus]          temp_m5_25_22_i;
wire signed [`CalcTempBus]          temp_m5_25_23_r;
wire signed [`CalcTempBus]          temp_m5_25_23_i;
wire signed [`CalcTempBus]          temp_m5_25_24_r;
wire signed [`CalcTempBus]          temp_m5_25_24_i;
wire signed [`CalcTempBus]          temp_m5_25_25_r;
wire signed [`CalcTempBus]          temp_m5_25_25_i;
wire signed [`CalcTempBus]          temp_m5_25_26_r;
wire signed [`CalcTempBus]          temp_m5_25_26_i;
wire signed [`CalcTempBus]          temp_m5_25_27_r;
wire signed [`CalcTempBus]          temp_m5_25_27_i;
wire signed [`CalcTempBus]          temp_m5_25_28_r;
wire signed [`CalcTempBus]          temp_m5_25_28_i;
wire signed [`CalcTempBus]          temp_m5_25_29_r;
wire signed [`CalcTempBus]          temp_m5_25_29_i;
wire signed [`CalcTempBus]          temp_m5_25_30_r;
wire signed [`CalcTempBus]          temp_m5_25_30_i;
wire signed [`CalcTempBus]          temp_m5_25_31_r;
wire signed [`CalcTempBus]          temp_m5_25_31_i;
wire signed [`CalcTempBus]          temp_m5_25_32_r;
wire signed [`CalcTempBus]          temp_m5_25_32_i;
wire signed [`CalcTempBus]          temp_m5_26_1_r;
wire signed [`CalcTempBus]          temp_m5_26_1_i;
wire signed [`CalcTempBus]          temp_m5_26_2_r;
wire signed [`CalcTempBus]          temp_m5_26_2_i;
wire signed [`CalcTempBus]          temp_m5_26_3_r;
wire signed [`CalcTempBus]          temp_m5_26_3_i;
wire signed [`CalcTempBus]          temp_m5_26_4_r;
wire signed [`CalcTempBus]          temp_m5_26_4_i;
wire signed [`CalcTempBus]          temp_m5_26_5_r;
wire signed [`CalcTempBus]          temp_m5_26_5_i;
wire signed [`CalcTempBus]          temp_m5_26_6_r;
wire signed [`CalcTempBus]          temp_m5_26_6_i;
wire signed [`CalcTempBus]          temp_m5_26_7_r;
wire signed [`CalcTempBus]          temp_m5_26_7_i;
wire signed [`CalcTempBus]          temp_m5_26_8_r;
wire signed [`CalcTempBus]          temp_m5_26_8_i;
wire signed [`CalcTempBus]          temp_m5_26_9_r;
wire signed [`CalcTempBus]          temp_m5_26_9_i;
wire signed [`CalcTempBus]          temp_m5_26_10_r;
wire signed [`CalcTempBus]          temp_m5_26_10_i;
wire signed [`CalcTempBus]          temp_m5_26_11_r;
wire signed [`CalcTempBus]          temp_m5_26_11_i;
wire signed [`CalcTempBus]          temp_m5_26_12_r;
wire signed [`CalcTempBus]          temp_m5_26_12_i;
wire signed [`CalcTempBus]          temp_m5_26_13_r;
wire signed [`CalcTempBus]          temp_m5_26_13_i;
wire signed [`CalcTempBus]          temp_m5_26_14_r;
wire signed [`CalcTempBus]          temp_m5_26_14_i;
wire signed [`CalcTempBus]          temp_m5_26_15_r;
wire signed [`CalcTempBus]          temp_m5_26_15_i;
wire signed [`CalcTempBus]          temp_m5_26_16_r;
wire signed [`CalcTempBus]          temp_m5_26_16_i;
wire signed [`CalcTempBus]          temp_m5_26_17_r;
wire signed [`CalcTempBus]          temp_m5_26_17_i;
wire signed [`CalcTempBus]          temp_m5_26_18_r;
wire signed [`CalcTempBus]          temp_m5_26_18_i;
wire signed [`CalcTempBus]          temp_m5_26_19_r;
wire signed [`CalcTempBus]          temp_m5_26_19_i;
wire signed [`CalcTempBus]          temp_m5_26_20_r;
wire signed [`CalcTempBus]          temp_m5_26_20_i;
wire signed [`CalcTempBus]          temp_m5_26_21_r;
wire signed [`CalcTempBus]          temp_m5_26_21_i;
wire signed [`CalcTempBus]          temp_m5_26_22_r;
wire signed [`CalcTempBus]          temp_m5_26_22_i;
wire signed [`CalcTempBus]          temp_m5_26_23_r;
wire signed [`CalcTempBus]          temp_m5_26_23_i;
wire signed [`CalcTempBus]          temp_m5_26_24_r;
wire signed [`CalcTempBus]          temp_m5_26_24_i;
wire signed [`CalcTempBus]          temp_m5_26_25_r;
wire signed [`CalcTempBus]          temp_m5_26_25_i;
wire signed [`CalcTempBus]          temp_m5_26_26_r;
wire signed [`CalcTempBus]          temp_m5_26_26_i;
wire signed [`CalcTempBus]          temp_m5_26_27_r;
wire signed [`CalcTempBus]          temp_m5_26_27_i;
wire signed [`CalcTempBus]          temp_m5_26_28_r;
wire signed [`CalcTempBus]          temp_m5_26_28_i;
wire signed [`CalcTempBus]          temp_m5_26_29_r;
wire signed [`CalcTempBus]          temp_m5_26_29_i;
wire signed [`CalcTempBus]          temp_m5_26_30_r;
wire signed [`CalcTempBus]          temp_m5_26_30_i;
wire signed [`CalcTempBus]          temp_m5_26_31_r;
wire signed [`CalcTempBus]          temp_m5_26_31_i;
wire signed [`CalcTempBus]          temp_m5_26_32_r;
wire signed [`CalcTempBus]          temp_m5_26_32_i;
wire signed [`CalcTempBus]          temp_m5_27_1_r;
wire signed [`CalcTempBus]          temp_m5_27_1_i;
wire signed [`CalcTempBus]          temp_m5_27_2_r;
wire signed [`CalcTempBus]          temp_m5_27_2_i;
wire signed [`CalcTempBus]          temp_m5_27_3_r;
wire signed [`CalcTempBus]          temp_m5_27_3_i;
wire signed [`CalcTempBus]          temp_m5_27_4_r;
wire signed [`CalcTempBus]          temp_m5_27_4_i;
wire signed [`CalcTempBus]          temp_m5_27_5_r;
wire signed [`CalcTempBus]          temp_m5_27_5_i;
wire signed [`CalcTempBus]          temp_m5_27_6_r;
wire signed [`CalcTempBus]          temp_m5_27_6_i;
wire signed [`CalcTempBus]          temp_m5_27_7_r;
wire signed [`CalcTempBus]          temp_m5_27_7_i;
wire signed [`CalcTempBus]          temp_m5_27_8_r;
wire signed [`CalcTempBus]          temp_m5_27_8_i;
wire signed [`CalcTempBus]          temp_m5_27_9_r;
wire signed [`CalcTempBus]          temp_m5_27_9_i;
wire signed [`CalcTempBus]          temp_m5_27_10_r;
wire signed [`CalcTempBus]          temp_m5_27_10_i;
wire signed [`CalcTempBus]          temp_m5_27_11_r;
wire signed [`CalcTempBus]          temp_m5_27_11_i;
wire signed [`CalcTempBus]          temp_m5_27_12_r;
wire signed [`CalcTempBus]          temp_m5_27_12_i;
wire signed [`CalcTempBus]          temp_m5_27_13_r;
wire signed [`CalcTempBus]          temp_m5_27_13_i;
wire signed [`CalcTempBus]          temp_m5_27_14_r;
wire signed [`CalcTempBus]          temp_m5_27_14_i;
wire signed [`CalcTempBus]          temp_m5_27_15_r;
wire signed [`CalcTempBus]          temp_m5_27_15_i;
wire signed [`CalcTempBus]          temp_m5_27_16_r;
wire signed [`CalcTempBus]          temp_m5_27_16_i;
wire signed [`CalcTempBus]          temp_m5_27_17_r;
wire signed [`CalcTempBus]          temp_m5_27_17_i;
wire signed [`CalcTempBus]          temp_m5_27_18_r;
wire signed [`CalcTempBus]          temp_m5_27_18_i;
wire signed [`CalcTempBus]          temp_m5_27_19_r;
wire signed [`CalcTempBus]          temp_m5_27_19_i;
wire signed [`CalcTempBus]          temp_m5_27_20_r;
wire signed [`CalcTempBus]          temp_m5_27_20_i;
wire signed [`CalcTempBus]          temp_m5_27_21_r;
wire signed [`CalcTempBus]          temp_m5_27_21_i;
wire signed [`CalcTempBus]          temp_m5_27_22_r;
wire signed [`CalcTempBus]          temp_m5_27_22_i;
wire signed [`CalcTempBus]          temp_m5_27_23_r;
wire signed [`CalcTempBus]          temp_m5_27_23_i;
wire signed [`CalcTempBus]          temp_m5_27_24_r;
wire signed [`CalcTempBus]          temp_m5_27_24_i;
wire signed [`CalcTempBus]          temp_m5_27_25_r;
wire signed [`CalcTempBus]          temp_m5_27_25_i;
wire signed [`CalcTempBus]          temp_m5_27_26_r;
wire signed [`CalcTempBus]          temp_m5_27_26_i;
wire signed [`CalcTempBus]          temp_m5_27_27_r;
wire signed [`CalcTempBus]          temp_m5_27_27_i;
wire signed [`CalcTempBus]          temp_m5_27_28_r;
wire signed [`CalcTempBus]          temp_m5_27_28_i;
wire signed [`CalcTempBus]          temp_m5_27_29_r;
wire signed [`CalcTempBus]          temp_m5_27_29_i;
wire signed [`CalcTempBus]          temp_m5_27_30_r;
wire signed [`CalcTempBus]          temp_m5_27_30_i;
wire signed [`CalcTempBus]          temp_m5_27_31_r;
wire signed [`CalcTempBus]          temp_m5_27_31_i;
wire signed [`CalcTempBus]          temp_m5_27_32_r;
wire signed [`CalcTempBus]          temp_m5_27_32_i;
wire signed [`CalcTempBus]          temp_m5_28_1_r;
wire signed [`CalcTempBus]          temp_m5_28_1_i;
wire signed [`CalcTempBus]          temp_m5_28_2_r;
wire signed [`CalcTempBus]          temp_m5_28_2_i;
wire signed [`CalcTempBus]          temp_m5_28_3_r;
wire signed [`CalcTempBus]          temp_m5_28_3_i;
wire signed [`CalcTempBus]          temp_m5_28_4_r;
wire signed [`CalcTempBus]          temp_m5_28_4_i;
wire signed [`CalcTempBus]          temp_m5_28_5_r;
wire signed [`CalcTempBus]          temp_m5_28_5_i;
wire signed [`CalcTempBus]          temp_m5_28_6_r;
wire signed [`CalcTempBus]          temp_m5_28_6_i;
wire signed [`CalcTempBus]          temp_m5_28_7_r;
wire signed [`CalcTempBus]          temp_m5_28_7_i;
wire signed [`CalcTempBus]          temp_m5_28_8_r;
wire signed [`CalcTempBus]          temp_m5_28_8_i;
wire signed [`CalcTempBus]          temp_m5_28_9_r;
wire signed [`CalcTempBus]          temp_m5_28_9_i;
wire signed [`CalcTempBus]          temp_m5_28_10_r;
wire signed [`CalcTempBus]          temp_m5_28_10_i;
wire signed [`CalcTempBus]          temp_m5_28_11_r;
wire signed [`CalcTempBus]          temp_m5_28_11_i;
wire signed [`CalcTempBus]          temp_m5_28_12_r;
wire signed [`CalcTempBus]          temp_m5_28_12_i;
wire signed [`CalcTempBus]          temp_m5_28_13_r;
wire signed [`CalcTempBus]          temp_m5_28_13_i;
wire signed [`CalcTempBus]          temp_m5_28_14_r;
wire signed [`CalcTempBus]          temp_m5_28_14_i;
wire signed [`CalcTempBus]          temp_m5_28_15_r;
wire signed [`CalcTempBus]          temp_m5_28_15_i;
wire signed [`CalcTempBus]          temp_m5_28_16_r;
wire signed [`CalcTempBus]          temp_m5_28_16_i;
wire signed [`CalcTempBus]          temp_m5_28_17_r;
wire signed [`CalcTempBus]          temp_m5_28_17_i;
wire signed [`CalcTempBus]          temp_m5_28_18_r;
wire signed [`CalcTempBus]          temp_m5_28_18_i;
wire signed [`CalcTempBus]          temp_m5_28_19_r;
wire signed [`CalcTempBus]          temp_m5_28_19_i;
wire signed [`CalcTempBus]          temp_m5_28_20_r;
wire signed [`CalcTempBus]          temp_m5_28_20_i;
wire signed [`CalcTempBus]          temp_m5_28_21_r;
wire signed [`CalcTempBus]          temp_m5_28_21_i;
wire signed [`CalcTempBus]          temp_m5_28_22_r;
wire signed [`CalcTempBus]          temp_m5_28_22_i;
wire signed [`CalcTempBus]          temp_m5_28_23_r;
wire signed [`CalcTempBus]          temp_m5_28_23_i;
wire signed [`CalcTempBus]          temp_m5_28_24_r;
wire signed [`CalcTempBus]          temp_m5_28_24_i;
wire signed [`CalcTempBus]          temp_m5_28_25_r;
wire signed [`CalcTempBus]          temp_m5_28_25_i;
wire signed [`CalcTempBus]          temp_m5_28_26_r;
wire signed [`CalcTempBus]          temp_m5_28_26_i;
wire signed [`CalcTempBus]          temp_m5_28_27_r;
wire signed [`CalcTempBus]          temp_m5_28_27_i;
wire signed [`CalcTempBus]          temp_m5_28_28_r;
wire signed [`CalcTempBus]          temp_m5_28_28_i;
wire signed [`CalcTempBus]          temp_m5_28_29_r;
wire signed [`CalcTempBus]          temp_m5_28_29_i;
wire signed [`CalcTempBus]          temp_m5_28_30_r;
wire signed [`CalcTempBus]          temp_m5_28_30_i;
wire signed [`CalcTempBus]          temp_m5_28_31_r;
wire signed [`CalcTempBus]          temp_m5_28_31_i;
wire signed [`CalcTempBus]          temp_m5_28_32_r;
wire signed [`CalcTempBus]          temp_m5_28_32_i;
wire signed [`CalcTempBus]          temp_m5_29_1_r;
wire signed [`CalcTempBus]          temp_m5_29_1_i;
wire signed [`CalcTempBus]          temp_m5_29_2_r;
wire signed [`CalcTempBus]          temp_m5_29_2_i;
wire signed [`CalcTempBus]          temp_m5_29_3_r;
wire signed [`CalcTempBus]          temp_m5_29_3_i;
wire signed [`CalcTempBus]          temp_m5_29_4_r;
wire signed [`CalcTempBus]          temp_m5_29_4_i;
wire signed [`CalcTempBus]          temp_m5_29_5_r;
wire signed [`CalcTempBus]          temp_m5_29_5_i;
wire signed [`CalcTempBus]          temp_m5_29_6_r;
wire signed [`CalcTempBus]          temp_m5_29_6_i;
wire signed [`CalcTempBus]          temp_m5_29_7_r;
wire signed [`CalcTempBus]          temp_m5_29_7_i;
wire signed [`CalcTempBus]          temp_m5_29_8_r;
wire signed [`CalcTempBus]          temp_m5_29_8_i;
wire signed [`CalcTempBus]          temp_m5_29_9_r;
wire signed [`CalcTempBus]          temp_m5_29_9_i;
wire signed [`CalcTempBus]          temp_m5_29_10_r;
wire signed [`CalcTempBus]          temp_m5_29_10_i;
wire signed [`CalcTempBus]          temp_m5_29_11_r;
wire signed [`CalcTempBus]          temp_m5_29_11_i;
wire signed [`CalcTempBus]          temp_m5_29_12_r;
wire signed [`CalcTempBus]          temp_m5_29_12_i;
wire signed [`CalcTempBus]          temp_m5_29_13_r;
wire signed [`CalcTempBus]          temp_m5_29_13_i;
wire signed [`CalcTempBus]          temp_m5_29_14_r;
wire signed [`CalcTempBus]          temp_m5_29_14_i;
wire signed [`CalcTempBus]          temp_m5_29_15_r;
wire signed [`CalcTempBus]          temp_m5_29_15_i;
wire signed [`CalcTempBus]          temp_m5_29_16_r;
wire signed [`CalcTempBus]          temp_m5_29_16_i;
wire signed [`CalcTempBus]          temp_m5_29_17_r;
wire signed [`CalcTempBus]          temp_m5_29_17_i;
wire signed [`CalcTempBus]          temp_m5_29_18_r;
wire signed [`CalcTempBus]          temp_m5_29_18_i;
wire signed [`CalcTempBus]          temp_m5_29_19_r;
wire signed [`CalcTempBus]          temp_m5_29_19_i;
wire signed [`CalcTempBus]          temp_m5_29_20_r;
wire signed [`CalcTempBus]          temp_m5_29_20_i;
wire signed [`CalcTempBus]          temp_m5_29_21_r;
wire signed [`CalcTempBus]          temp_m5_29_21_i;
wire signed [`CalcTempBus]          temp_m5_29_22_r;
wire signed [`CalcTempBus]          temp_m5_29_22_i;
wire signed [`CalcTempBus]          temp_m5_29_23_r;
wire signed [`CalcTempBus]          temp_m5_29_23_i;
wire signed [`CalcTempBus]          temp_m5_29_24_r;
wire signed [`CalcTempBus]          temp_m5_29_24_i;
wire signed [`CalcTempBus]          temp_m5_29_25_r;
wire signed [`CalcTempBus]          temp_m5_29_25_i;
wire signed [`CalcTempBus]          temp_m5_29_26_r;
wire signed [`CalcTempBus]          temp_m5_29_26_i;
wire signed [`CalcTempBus]          temp_m5_29_27_r;
wire signed [`CalcTempBus]          temp_m5_29_27_i;
wire signed [`CalcTempBus]          temp_m5_29_28_r;
wire signed [`CalcTempBus]          temp_m5_29_28_i;
wire signed [`CalcTempBus]          temp_m5_29_29_r;
wire signed [`CalcTempBus]          temp_m5_29_29_i;
wire signed [`CalcTempBus]          temp_m5_29_30_r;
wire signed [`CalcTempBus]          temp_m5_29_30_i;
wire signed [`CalcTempBus]          temp_m5_29_31_r;
wire signed [`CalcTempBus]          temp_m5_29_31_i;
wire signed [`CalcTempBus]          temp_m5_29_32_r;
wire signed [`CalcTempBus]          temp_m5_29_32_i;
wire signed [`CalcTempBus]          temp_m5_30_1_r;
wire signed [`CalcTempBus]          temp_m5_30_1_i;
wire signed [`CalcTempBus]          temp_m5_30_2_r;
wire signed [`CalcTempBus]          temp_m5_30_2_i;
wire signed [`CalcTempBus]          temp_m5_30_3_r;
wire signed [`CalcTempBus]          temp_m5_30_3_i;
wire signed [`CalcTempBus]          temp_m5_30_4_r;
wire signed [`CalcTempBus]          temp_m5_30_4_i;
wire signed [`CalcTempBus]          temp_m5_30_5_r;
wire signed [`CalcTempBus]          temp_m5_30_5_i;
wire signed [`CalcTempBus]          temp_m5_30_6_r;
wire signed [`CalcTempBus]          temp_m5_30_6_i;
wire signed [`CalcTempBus]          temp_m5_30_7_r;
wire signed [`CalcTempBus]          temp_m5_30_7_i;
wire signed [`CalcTempBus]          temp_m5_30_8_r;
wire signed [`CalcTempBus]          temp_m5_30_8_i;
wire signed [`CalcTempBus]          temp_m5_30_9_r;
wire signed [`CalcTempBus]          temp_m5_30_9_i;
wire signed [`CalcTempBus]          temp_m5_30_10_r;
wire signed [`CalcTempBus]          temp_m5_30_10_i;
wire signed [`CalcTempBus]          temp_m5_30_11_r;
wire signed [`CalcTempBus]          temp_m5_30_11_i;
wire signed [`CalcTempBus]          temp_m5_30_12_r;
wire signed [`CalcTempBus]          temp_m5_30_12_i;
wire signed [`CalcTempBus]          temp_m5_30_13_r;
wire signed [`CalcTempBus]          temp_m5_30_13_i;
wire signed [`CalcTempBus]          temp_m5_30_14_r;
wire signed [`CalcTempBus]          temp_m5_30_14_i;
wire signed [`CalcTempBus]          temp_m5_30_15_r;
wire signed [`CalcTempBus]          temp_m5_30_15_i;
wire signed [`CalcTempBus]          temp_m5_30_16_r;
wire signed [`CalcTempBus]          temp_m5_30_16_i;
wire signed [`CalcTempBus]          temp_m5_30_17_r;
wire signed [`CalcTempBus]          temp_m5_30_17_i;
wire signed [`CalcTempBus]          temp_m5_30_18_r;
wire signed [`CalcTempBus]          temp_m5_30_18_i;
wire signed [`CalcTempBus]          temp_m5_30_19_r;
wire signed [`CalcTempBus]          temp_m5_30_19_i;
wire signed [`CalcTempBus]          temp_m5_30_20_r;
wire signed [`CalcTempBus]          temp_m5_30_20_i;
wire signed [`CalcTempBus]          temp_m5_30_21_r;
wire signed [`CalcTempBus]          temp_m5_30_21_i;
wire signed [`CalcTempBus]          temp_m5_30_22_r;
wire signed [`CalcTempBus]          temp_m5_30_22_i;
wire signed [`CalcTempBus]          temp_m5_30_23_r;
wire signed [`CalcTempBus]          temp_m5_30_23_i;
wire signed [`CalcTempBus]          temp_m5_30_24_r;
wire signed [`CalcTempBus]          temp_m5_30_24_i;
wire signed [`CalcTempBus]          temp_m5_30_25_r;
wire signed [`CalcTempBus]          temp_m5_30_25_i;
wire signed [`CalcTempBus]          temp_m5_30_26_r;
wire signed [`CalcTempBus]          temp_m5_30_26_i;
wire signed [`CalcTempBus]          temp_m5_30_27_r;
wire signed [`CalcTempBus]          temp_m5_30_27_i;
wire signed [`CalcTempBus]          temp_m5_30_28_r;
wire signed [`CalcTempBus]          temp_m5_30_28_i;
wire signed [`CalcTempBus]          temp_m5_30_29_r;
wire signed [`CalcTempBus]          temp_m5_30_29_i;
wire signed [`CalcTempBus]          temp_m5_30_30_r;
wire signed [`CalcTempBus]          temp_m5_30_30_i;
wire signed [`CalcTempBus]          temp_m5_30_31_r;
wire signed [`CalcTempBus]          temp_m5_30_31_i;
wire signed [`CalcTempBus]          temp_m5_30_32_r;
wire signed [`CalcTempBus]          temp_m5_30_32_i;
wire signed [`CalcTempBus]          temp_m5_31_1_r;
wire signed [`CalcTempBus]          temp_m5_31_1_i;
wire signed [`CalcTempBus]          temp_m5_31_2_r;
wire signed [`CalcTempBus]          temp_m5_31_2_i;
wire signed [`CalcTempBus]          temp_m5_31_3_r;
wire signed [`CalcTempBus]          temp_m5_31_3_i;
wire signed [`CalcTempBus]          temp_m5_31_4_r;
wire signed [`CalcTempBus]          temp_m5_31_4_i;
wire signed [`CalcTempBus]          temp_m5_31_5_r;
wire signed [`CalcTempBus]          temp_m5_31_5_i;
wire signed [`CalcTempBus]          temp_m5_31_6_r;
wire signed [`CalcTempBus]          temp_m5_31_6_i;
wire signed [`CalcTempBus]          temp_m5_31_7_r;
wire signed [`CalcTempBus]          temp_m5_31_7_i;
wire signed [`CalcTempBus]          temp_m5_31_8_r;
wire signed [`CalcTempBus]          temp_m5_31_8_i;
wire signed [`CalcTempBus]          temp_m5_31_9_r;
wire signed [`CalcTempBus]          temp_m5_31_9_i;
wire signed [`CalcTempBus]          temp_m5_31_10_r;
wire signed [`CalcTempBus]          temp_m5_31_10_i;
wire signed [`CalcTempBus]          temp_m5_31_11_r;
wire signed [`CalcTempBus]          temp_m5_31_11_i;
wire signed [`CalcTempBus]          temp_m5_31_12_r;
wire signed [`CalcTempBus]          temp_m5_31_12_i;
wire signed [`CalcTempBus]          temp_m5_31_13_r;
wire signed [`CalcTempBus]          temp_m5_31_13_i;
wire signed [`CalcTempBus]          temp_m5_31_14_r;
wire signed [`CalcTempBus]          temp_m5_31_14_i;
wire signed [`CalcTempBus]          temp_m5_31_15_r;
wire signed [`CalcTempBus]          temp_m5_31_15_i;
wire signed [`CalcTempBus]          temp_m5_31_16_r;
wire signed [`CalcTempBus]          temp_m5_31_16_i;
wire signed [`CalcTempBus]          temp_m5_31_17_r;
wire signed [`CalcTempBus]          temp_m5_31_17_i;
wire signed [`CalcTempBus]          temp_m5_31_18_r;
wire signed [`CalcTempBus]          temp_m5_31_18_i;
wire signed [`CalcTempBus]          temp_m5_31_19_r;
wire signed [`CalcTempBus]          temp_m5_31_19_i;
wire signed [`CalcTempBus]          temp_m5_31_20_r;
wire signed [`CalcTempBus]          temp_m5_31_20_i;
wire signed [`CalcTempBus]          temp_m5_31_21_r;
wire signed [`CalcTempBus]          temp_m5_31_21_i;
wire signed [`CalcTempBus]          temp_m5_31_22_r;
wire signed [`CalcTempBus]          temp_m5_31_22_i;
wire signed [`CalcTempBus]          temp_m5_31_23_r;
wire signed [`CalcTempBus]          temp_m5_31_23_i;
wire signed [`CalcTempBus]          temp_m5_31_24_r;
wire signed [`CalcTempBus]          temp_m5_31_24_i;
wire signed [`CalcTempBus]          temp_m5_31_25_r;
wire signed [`CalcTempBus]          temp_m5_31_25_i;
wire signed [`CalcTempBus]          temp_m5_31_26_r;
wire signed [`CalcTempBus]          temp_m5_31_26_i;
wire signed [`CalcTempBus]          temp_m5_31_27_r;
wire signed [`CalcTempBus]          temp_m5_31_27_i;
wire signed [`CalcTempBus]          temp_m5_31_28_r;
wire signed [`CalcTempBus]          temp_m5_31_28_i;
wire signed [`CalcTempBus]          temp_m5_31_29_r;
wire signed [`CalcTempBus]          temp_m5_31_29_i;
wire signed [`CalcTempBus]          temp_m5_31_30_r;
wire signed [`CalcTempBus]          temp_m5_31_30_i;
wire signed [`CalcTempBus]          temp_m5_31_31_r;
wire signed [`CalcTempBus]          temp_m5_31_31_i;
wire signed [`CalcTempBus]          temp_m5_31_32_r;
wire signed [`CalcTempBus]          temp_m5_31_32_i;
wire signed [`CalcTempBus]          temp_m5_32_1_r;
wire signed [`CalcTempBus]          temp_m5_32_1_i;
wire signed [`CalcTempBus]          temp_m5_32_2_r;
wire signed [`CalcTempBus]          temp_m5_32_2_i;
wire signed [`CalcTempBus]          temp_m5_32_3_r;
wire signed [`CalcTempBus]          temp_m5_32_3_i;
wire signed [`CalcTempBus]          temp_m5_32_4_r;
wire signed [`CalcTempBus]          temp_m5_32_4_i;
wire signed [`CalcTempBus]          temp_m5_32_5_r;
wire signed [`CalcTempBus]          temp_m5_32_5_i;
wire signed [`CalcTempBus]          temp_m5_32_6_r;
wire signed [`CalcTempBus]          temp_m5_32_6_i;
wire signed [`CalcTempBus]          temp_m5_32_7_r;
wire signed [`CalcTempBus]          temp_m5_32_7_i;
wire signed [`CalcTempBus]          temp_m5_32_8_r;
wire signed [`CalcTempBus]          temp_m5_32_8_i;
wire signed [`CalcTempBus]          temp_m5_32_9_r;
wire signed [`CalcTempBus]          temp_m5_32_9_i;
wire signed [`CalcTempBus]          temp_m5_32_10_r;
wire signed [`CalcTempBus]          temp_m5_32_10_i;
wire signed [`CalcTempBus]          temp_m5_32_11_r;
wire signed [`CalcTempBus]          temp_m5_32_11_i;
wire signed [`CalcTempBus]          temp_m5_32_12_r;
wire signed [`CalcTempBus]          temp_m5_32_12_i;
wire signed [`CalcTempBus]          temp_m5_32_13_r;
wire signed [`CalcTempBus]          temp_m5_32_13_i;
wire signed [`CalcTempBus]          temp_m5_32_14_r;
wire signed [`CalcTempBus]          temp_m5_32_14_i;
wire signed [`CalcTempBus]          temp_m5_32_15_r;
wire signed [`CalcTempBus]          temp_m5_32_15_i;
wire signed [`CalcTempBus]          temp_m5_32_16_r;
wire signed [`CalcTempBus]          temp_m5_32_16_i;
wire signed [`CalcTempBus]          temp_m5_32_17_r;
wire signed [`CalcTempBus]          temp_m5_32_17_i;
wire signed [`CalcTempBus]          temp_m5_32_18_r;
wire signed [`CalcTempBus]          temp_m5_32_18_i;
wire signed [`CalcTempBus]          temp_m5_32_19_r;
wire signed [`CalcTempBus]          temp_m5_32_19_i;
wire signed [`CalcTempBus]          temp_m5_32_20_r;
wire signed [`CalcTempBus]          temp_m5_32_20_i;
wire signed [`CalcTempBus]          temp_m5_32_21_r;
wire signed [`CalcTempBus]          temp_m5_32_21_i;
wire signed [`CalcTempBus]          temp_m5_32_22_r;
wire signed [`CalcTempBus]          temp_m5_32_22_i;
wire signed [`CalcTempBus]          temp_m5_32_23_r;
wire signed [`CalcTempBus]          temp_m5_32_23_i;
wire signed [`CalcTempBus]          temp_m5_32_24_r;
wire signed [`CalcTempBus]          temp_m5_32_24_i;
wire signed [`CalcTempBus]          temp_m5_32_25_r;
wire signed [`CalcTempBus]          temp_m5_32_25_i;
wire signed [`CalcTempBus]          temp_m5_32_26_r;
wire signed [`CalcTempBus]          temp_m5_32_26_i;
wire signed [`CalcTempBus]          temp_m5_32_27_r;
wire signed [`CalcTempBus]          temp_m5_32_27_i;
wire signed [`CalcTempBus]          temp_m5_32_28_r;
wire signed [`CalcTempBus]          temp_m5_32_28_i;
wire signed [`CalcTempBus]          temp_m5_32_29_r;
wire signed [`CalcTempBus]          temp_m5_32_29_i;
wire signed [`CalcTempBus]          temp_m5_32_30_r;
wire signed [`CalcTempBus]          temp_m5_32_30_i;
wire signed [`CalcTempBus]          temp_m5_32_31_r;
wire signed [`CalcTempBus]          temp_m5_32_31_i;
wire signed [`CalcTempBus]          temp_m5_32_32_r;
wire signed [`CalcTempBus]          temp_m5_32_32_i;

wire signed [`CalcTempBus]          temp_b1_1_1_r;
wire signed [`CalcTempBus]          temp_b1_1_1_i;
wire signed [`CalcTempBus]          temp_b1_1_2_r;
wire signed [`CalcTempBus]          temp_b1_1_2_i;
wire signed [`CalcTempBus]          temp_b1_1_3_r;
wire signed [`CalcTempBus]          temp_b1_1_3_i;
wire signed [`CalcTempBus]          temp_b1_1_4_r;
wire signed [`CalcTempBus]          temp_b1_1_4_i;
wire signed [`CalcTempBus]          temp_b1_1_5_r;
wire signed [`CalcTempBus]          temp_b1_1_5_i;
wire signed [`CalcTempBus]          temp_b1_1_6_r;
wire signed [`CalcTempBus]          temp_b1_1_6_i;
wire signed [`CalcTempBus]          temp_b1_1_7_r;
wire signed [`CalcTempBus]          temp_b1_1_7_i;
wire signed [`CalcTempBus]          temp_b1_1_8_r;
wire signed [`CalcTempBus]          temp_b1_1_8_i;
wire signed [`CalcTempBus]          temp_b1_1_9_r;
wire signed [`CalcTempBus]          temp_b1_1_9_i;
wire signed [`CalcTempBus]          temp_b1_1_10_r;
wire signed [`CalcTempBus]          temp_b1_1_10_i;
wire signed [`CalcTempBus]          temp_b1_1_11_r;
wire signed [`CalcTempBus]          temp_b1_1_11_i;
wire signed [`CalcTempBus]          temp_b1_1_12_r;
wire signed [`CalcTempBus]          temp_b1_1_12_i;
wire signed [`CalcTempBus]          temp_b1_1_13_r;
wire signed [`CalcTempBus]          temp_b1_1_13_i;
wire signed [`CalcTempBus]          temp_b1_1_14_r;
wire signed [`CalcTempBus]          temp_b1_1_14_i;
wire signed [`CalcTempBus]          temp_b1_1_15_r;
wire signed [`CalcTempBus]          temp_b1_1_15_i;
wire signed [`CalcTempBus]          temp_b1_1_16_r;
wire signed [`CalcTempBus]          temp_b1_1_16_i;
wire signed [`CalcTempBus]          temp_b1_1_17_r;
wire signed [`CalcTempBus]          temp_b1_1_17_i;
wire signed [`CalcTempBus]          temp_b1_1_18_r;
wire signed [`CalcTempBus]          temp_b1_1_18_i;
wire signed [`CalcTempBus]          temp_b1_1_19_r;
wire signed [`CalcTempBus]          temp_b1_1_19_i;
wire signed [`CalcTempBus]          temp_b1_1_20_r;
wire signed [`CalcTempBus]          temp_b1_1_20_i;
wire signed [`CalcTempBus]          temp_b1_1_21_r;
wire signed [`CalcTempBus]          temp_b1_1_21_i;
wire signed [`CalcTempBus]          temp_b1_1_22_r;
wire signed [`CalcTempBus]          temp_b1_1_22_i;
wire signed [`CalcTempBus]          temp_b1_1_23_r;
wire signed [`CalcTempBus]          temp_b1_1_23_i;
wire signed [`CalcTempBus]          temp_b1_1_24_r;
wire signed [`CalcTempBus]          temp_b1_1_24_i;
wire signed [`CalcTempBus]          temp_b1_1_25_r;
wire signed [`CalcTempBus]          temp_b1_1_25_i;
wire signed [`CalcTempBus]          temp_b1_1_26_r;
wire signed [`CalcTempBus]          temp_b1_1_26_i;
wire signed [`CalcTempBus]          temp_b1_1_27_r;
wire signed [`CalcTempBus]          temp_b1_1_27_i;
wire signed [`CalcTempBus]          temp_b1_1_28_r;
wire signed [`CalcTempBus]          temp_b1_1_28_i;
wire signed [`CalcTempBus]          temp_b1_1_29_r;
wire signed [`CalcTempBus]          temp_b1_1_29_i;
wire signed [`CalcTempBus]          temp_b1_1_30_r;
wire signed [`CalcTempBus]          temp_b1_1_30_i;
wire signed [`CalcTempBus]          temp_b1_1_31_r;
wire signed [`CalcTempBus]          temp_b1_1_31_i;
wire signed [`CalcTempBus]          temp_b1_1_32_r;
wire signed [`CalcTempBus]          temp_b1_1_32_i;
wire signed [`CalcTempBus]          temp_b1_2_1_r;
wire signed [`CalcTempBus]          temp_b1_2_1_i;
wire signed [`CalcTempBus]          temp_b1_2_2_r;
wire signed [`CalcTempBus]          temp_b1_2_2_i;
wire signed [`CalcTempBus]          temp_b1_2_3_r;
wire signed [`CalcTempBus]          temp_b1_2_3_i;
wire signed [`CalcTempBus]          temp_b1_2_4_r;
wire signed [`CalcTempBus]          temp_b1_2_4_i;
wire signed [`CalcTempBus]          temp_b1_2_5_r;
wire signed [`CalcTempBus]          temp_b1_2_5_i;
wire signed [`CalcTempBus]          temp_b1_2_6_r;
wire signed [`CalcTempBus]          temp_b1_2_6_i;
wire signed [`CalcTempBus]          temp_b1_2_7_r;
wire signed [`CalcTempBus]          temp_b1_2_7_i;
wire signed [`CalcTempBus]          temp_b1_2_8_r;
wire signed [`CalcTempBus]          temp_b1_2_8_i;
wire signed [`CalcTempBus]          temp_b1_2_9_r;
wire signed [`CalcTempBus]          temp_b1_2_9_i;
wire signed [`CalcTempBus]          temp_b1_2_10_r;
wire signed [`CalcTempBus]          temp_b1_2_10_i;
wire signed [`CalcTempBus]          temp_b1_2_11_r;
wire signed [`CalcTempBus]          temp_b1_2_11_i;
wire signed [`CalcTempBus]          temp_b1_2_12_r;
wire signed [`CalcTempBus]          temp_b1_2_12_i;
wire signed [`CalcTempBus]          temp_b1_2_13_r;
wire signed [`CalcTempBus]          temp_b1_2_13_i;
wire signed [`CalcTempBus]          temp_b1_2_14_r;
wire signed [`CalcTempBus]          temp_b1_2_14_i;
wire signed [`CalcTempBus]          temp_b1_2_15_r;
wire signed [`CalcTempBus]          temp_b1_2_15_i;
wire signed [`CalcTempBus]          temp_b1_2_16_r;
wire signed [`CalcTempBus]          temp_b1_2_16_i;
wire signed [`CalcTempBus]          temp_b1_2_17_r;
wire signed [`CalcTempBus]          temp_b1_2_17_i;
wire signed [`CalcTempBus]          temp_b1_2_18_r;
wire signed [`CalcTempBus]          temp_b1_2_18_i;
wire signed [`CalcTempBus]          temp_b1_2_19_r;
wire signed [`CalcTempBus]          temp_b1_2_19_i;
wire signed [`CalcTempBus]          temp_b1_2_20_r;
wire signed [`CalcTempBus]          temp_b1_2_20_i;
wire signed [`CalcTempBus]          temp_b1_2_21_r;
wire signed [`CalcTempBus]          temp_b1_2_21_i;
wire signed [`CalcTempBus]          temp_b1_2_22_r;
wire signed [`CalcTempBus]          temp_b1_2_22_i;
wire signed [`CalcTempBus]          temp_b1_2_23_r;
wire signed [`CalcTempBus]          temp_b1_2_23_i;
wire signed [`CalcTempBus]          temp_b1_2_24_r;
wire signed [`CalcTempBus]          temp_b1_2_24_i;
wire signed [`CalcTempBus]          temp_b1_2_25_r;
wire signed [`CalcTempBus]          temp_b1_2_25_i;
wire signed [`CalcTempBus]          temp_b1_2_26_r;
wire signed [`CalcTempBus]          temp_b1_2_26_i;
wire signed [`CalcTempBus]          temp_b1_2_27_r;
wire signed [`CalcTempBus]          temp_b1_2_27_i;
wire signed [`CalcTempBus]          temp_b1_2_28_r;
wire signed [`CalcTempBus]          temp_b1_2_28_i;
wire signed [`CalcTempBus]          temp_b1_2_29_r;
wire signed [`CalcTempBus]          temp_b1_2_29_i;
wire signed [`CalcTempBus]          temp_b1_2_30_r;
wire signed [`CalcTempBus]          temp_b1_2_30_i;
wire signed [`CalcTempBus]          temp_b1_2_31_r;
wire signed [`CalcTempBus]          temp_b1_2_31_i;
wire signed [`CalcTempBus]          temp_b1_2_32_r;
wire signed [`CalcTempBus]          temp_b1_2_32_i;
wire signed [`CalcTempBus]          temp_b1_3_1_r;
wire signed [`CalcTempBus]          temp_b1_3_1_i;
wire signed [`CalcTempBus]          temp_b1_3_2_r;
wire signed [`CalcTempBus]          temp_b1_3_2_i;
wire signed [`CalcTempBus]          temp_b1_3_3_r;
wire signed [`CalcTempBus]          temp_b1_3_3_i;
wire signed [`CalcTempBus]          temp_b1_3_4_r;
wire signed [`CalcTempBus]          temp_b1_3_4_i;
wire signed [`CalcTempBus]          temp_b1_3_5_r;
wire signed [`CalcTempBus]          temp_b1_3_5_i;
wire signed [`CalcTempBus]          temp_b1_3_6_r;
wire signed [`CalcTempBus]          temp_b1_3_6_i;
wire signed [`CalcTempBus]          temp_b1_3_7_r;
wire signed [`CalcTempBus]          temp_b1_3_7_i;
wire signed [`CalcTempBus]          temp_b1_3_8_r;
wire signed [`CalcTempBus]          temp_b1_3_8_i;
wire signed [`CalcTempBus]          temp_b1_3_9_r;
wire signed [`CalcTempBus]          temp_b1_3_9_i;
wire signed [`CalcTempBus]          temp_b1_3_10_r;
wire signed [`CalcTempBus]          temp_b1_3_10_i;
wire signed [`CalcTempBus]          temp_b1_3_11_r;
wire signed [`CalcTempBus]          temp_b1_3_11_i;
wire signed [`CalcTempBus]          temp_b1_3_12_r;
wire signed [`CalcTempBus]          temp_b1_3_12_i;
wire signed [`CalcTempBus]          temp_b1_3_13_r;
wire signed [`CalcTempBus]          temp_b1_3_13_i;
wire signed [`CalcTempBus]          temp_b1_3_14_r;
wire signed [`CalcTempBus]          temp_b1_3_14_i;
wire signed [`CalcTempBus]          temp_b1_3_15_r;
wire signed [`CalcTempBus]          temp_b1_3_15_i;
wire signed [`CalcTempBus]          temp_b1_3_16_r;
wire signed [`CalcTempBus]          temp_b1_3_16_i;
wire signed [`CalcTempBus]          temp_b1_3_17_r;
wire signed [`CalcTempBus]          temp_b1_3_17_i;
wire signed [`CalcTempBus]          temp_b1_3_18_r;
wire signed [`CalcTempBus]          temp_b1_3_18_i;
wire signed [`CalcTempBus]          temp_b1_3_19_r;
wire signed [`CalcTempBus]          temp_b1_3_19_i;
wire signed [`CalcTempBus]          temp_b1_3_20_r;
wire signed [`CalcTempBus]          temp_b1_3_20_i;
wire signed [`CalcTempBus]          temp_b1_3_21_r;
wire signed [`CalcTempBus]          temp_b1_3_21_i;
wire signed [`CalcTempBus]          temp_b1_3_22_r;
wire signed [`CalcTempBus]          temp_b1_3_22_i;
wire signed [`CalcTempBus]          temp_b1_3_23_r;
wire signed [`CalcTempBus]          temp_b1_3_23_i;
wire signed [`CalcTempBus]          temp_b1_3_24_r;
wire signed [`CalcTempBus]          temp_b1_3_24_i;
wire signed [`CalcTempBus]          temp_b1_3_25_r;
wire signed [`CalcTempBus]          temp_b1_3_25_i;
wire signed [`CalcTempBus]          temp_b1_3_26_r;
wire signed [`CalcTempBus]          temp_b1_3_26_i;
wire signed [`CalcTempBus]          temp_b1_3_27_r;
wire signed [`CalcTempBus]          temp_b1_3_27_i;
wire signed [`CalcTempBus]          temp_b1_3_28_r;
wire signed [`CalcTempBus]          temp_b1_3_28_i;
wire signed [`CalcTempBus]          temp_b1_3_29_r;
wire signed [`CalcTempBus]          temp_b1_3_29_i;
wire signed [`CalcTempBus]          temp_b1_3_30_r;
wire signed [`CalcTempBus]          temp_b1_3_30_i;
wire signed [`CalcTempBus]          temp_b1_3_31_r;
wire signed [`CalcTempBus]          temp_b1_3_31_i;
wire signed [`CalcTempBus]          temp_b1_3_32_r;
wire signed [`CalcTempBus]          temp_b1_3_32_i;
wire signed [`CalcTempBus]          temp_b1_4_1_r;
wire signed [`CalcTempBus]          temp_b1_4_1_i;
wire signed [`CalcTempBus]          temp_b1_4_2_r;
wire signed [`CalcTempBus]          temp_b1_4_2_i;
wire signed [`CalcTempBus]          temp_b1_4_3_r;
wire signed [`CalcTempBus]          temp_b1_4_3_i;
wire signed [`CalcTempBus]          temp_b1_4_4_r;
wire signed [`CalcTempBus]          temp_b1_4_4_i;
wire signed [`CalcTempBus]          temp_b1_4_5_r;
wire signed [`CalcTempBus]          temp_b1_4_5_i;
wire signed [`CalcTempBus]          temp_b1_4_6_r;
wire signed [`CalcTempBus]          temp_b1_4_6_i;
wire signed [`CalcTempBus]          temp_b1_4_7_r;
wire signed [`CalcTempBus]          temp_b1_4_7_i;
wire signed [`CalcTempBus]          temp_b1_4_8_r;
wire signed [`CalcTempBus]          temp_b1_4_8_i;
wire signed [`CalcTempBus]          temp_b1_4_9_r;
wire signed [`CalcTempBus]          temp_b1_4_9_i;
wire signed [`CalcTempBus]          temp_b1_4_10_r;
wire signed [`CalcTempBus]          temp_b1_4_10_i;
wire signed [`CalcTempBus]          temp_b1_4_11_r;
wire signed [`CalcTempBus]          temp_b1_4_11_i;
wire signed [`CalcTempBus]          temp_b1_4_12_r;
wire signed [`CalcTempBus]          temp_b1_4_12_i;
wire signed [`CalcTempBus]          temp_b1_4_13_r;
wire signed [`CalcTempBus]          temp_b1_4_13_i;
wire signed [`CalcTempBus]          temp_b1_4_14_r;
wire signed [`CalcTempBus]          temp_b1_4_14_i;
wire signed [`CalcTempBus]          temp_b1_4_15_r;
wire signed [`CalcTempBus]          temp_b1_4_15_i;
wire signed [`CalcTempBus]          temp_b1_4_16_r;
wire signed [`CalcTempBus]          temp_b1_4_16_i;
wire signed [`CalcTempBus]          temp_b1_4_17_r;
wire signed [`CalcTempBus]          temp_b1_4_17_i;
wire signed [`CalcTempBus]          temp_b1_4_18_r;
wire signed [`CalcTempBus]          temp_b1_4_18_i;
wire signed [`CalcTempBus]          temp_b1_4_19_r;
wire signed [`CalcTempBus]          temp_b1_4_19_i;
wire signed [`CalcTempBus]          temp_b1_4_20_r;
wire signed [`CalcTempBus]          temp_b1_4_20_i;
wire signed [`CalcTempBus]          temp_b1_4_21_r;
wire signed [`CalcTempBus]          temp_b1_4_21_i;
wire signed [`CalcTempBus]          temp_b1_4_22_r;
wire signed [`CalcTempBus]          temp_b1_4_22_i;
wire signed [`CalcTempBus]          temp_b1_4_23_r;
wire signed [`CalcTempBus]          temp_b1_4_23_i;
wire signed [`CalcTempBus]          temp_b1_4_24_r;
wire signed [`CalcTempBus]          temp_b1_4_24_i;
wire signed [`CalcTempBus]          temp_b1_4_25_r;
wire signed [`CalcTempBus]          temp_b1_4_25_i;
wire signed [`CalcTempBus]          temp_b1_4_26_r;
wire signed [`CalcTempBus]          temp_b1_4_26_i;
wire signed [`CalcTempBus]          temp_b1_4_27_r;
wire signed [`CalcTempBus]          temp_b1_4_27_i;
wire signed [`CalcTempBus]          temp_b1_4_28_r;
wire signed [`CalcTempBus]          temp_b1_4_28_i;
wire signed [`CalcTempBus]          temp_b1_4_29_r;
wire signed [`CalcTempBus]          temp_b1_4_29_i;
wire signed [`CalcTempBus]          temp_b1_4_30_r;
wire signed [`CalcTempBus]          temp_b1_4_30_i;
wire signed [`CalcTempBus]          temp_b1_4_31_r;
wire signed [`CalcTempBus]          temp_b1_4_31_i;
wire signed [`CalcTempBus]          temp_b1_4_32_r;
wire signed [`CalcTempBus]          temp_b1_4_32_i;
wire signed [`CalcTempBus]          temp_b1_5_1_r;
wire signed [`CalcTempBus]          temp_b1_5_1_i;
wire signed [`CalcTempBus]          temp_b1_5_2_r;
wire signed [`CalcTempBus]          temp_b1_5_2_i;
wire signed [`CalcTempBus]          temp_b1_5_3_r;
wire signed [`CalcTempBus]          temp_b1_5_3_i;
wire signed [`CalcTempBus]          temp_b1_5_4_r;
wire signed [`CalcTempBus]          temp_b1_5_4_i;
wire signed [`CalcTempBus]          temp_b1_5_5_r;
wire signed [`CalcTempBus]          temp_b1_5_5_i;
wire signed [`CalcTempBus]          temp_b1_5_6_r;
wire signed [`CalcTempBus]          temp_b1_5_6_i;
wire signed [`CalcTempBus]          temp_b1_5_7_r;
wire signed [`CalcTempBus]          temp_b1_5_7_i;
wire signed [`CalcTempBus]          temp_b1_5_8_r;
wire signed [`CalcTempBus]          temp_b1_5_8_i;
wire signed [`CalcTempBus]          temp_b1_5_9_r;
wire signed [`CalcTempBus]          temp_b1_5_9_i;
wire signed [`CalcTempBus]          temp_b1_5_10_r;
wire signed [`CalcTempBus]          temp_b1_5_10_i;
wire signed [`CalcTempBus]          temp_b1_5_11_r;
wire signed [`CalcTempBus]          temp_b1_5_11_i;
wire signed [`CalcTempBus]          temp_b1_5_12_r;
wire signed [`CalcTempBus]          temp_b1_5_12_i;
wire signed [`CalcTempBus]          temp_b1_5_13_r;
wire signed [`CalcTempBus]          temp_b1_5_13_i;
wire signed [`CalcTempBus]          temp_b1_5_14_r;
wire signed [`CalcTempBus]          temp_b1_5_14_i;
wire signed [`CalcTempBus]          temp_b1_5_15_r;
wire signed [`CalcTempBus]          temp_b1_5_15_i;
wire signed [`CalcTempBus]          temp_b1_5_16_r;
wire signed [`CalcTempBus]          temp_b1_5_16_i;
wire signed [`CalcTempBus]          temp_b1_5_17_r;
wire signed [`CalcTempBus]          temp_b1_5_17_i;
wire signed [`CalcTempBus]          temp_b1_5_18_r;
wire signed [`CalcTempBus]          temp_b1_5_18_i;
wire signed [`CalcTempBus]          temp_b1_5_19_r;
wire signed [`CalcTempBus]          temp_b1_5_19_i;
wire signed [`CalcTempBus]          temp_b1_5_20_r;
wire signed [`CalcTempBus]          temp_b1_5_20_i;
wire signed [`CalcTempBus]          temp_b1_5_21_r;
wire signed [`CalcTempBus]          temp_b1_5_21_i;
wire signed [`CalcTempBus]          temp_b1_5_22_r;
wire signed [`CalcTempBus]          temp_b1_5_22_i;
wire signed [`CalcTempBus]          temp_b1_5_23_r;
wire signed [`CalcTempBus]          temp_b1_5_23_i;
wire signed [`CalcTempBus]          temp_b1_5_24_r;
wire signed [`CalcTempBus]          temp_b1_5_24_i;
wire signed [`CalcTempBus]          temp_b1_5_25_r;
wire signed [`CalcTempBus]          temp_b1_5_25_i;
wire signed [`CalcTempBus]          temp_b1_5_26_r;
wire signed [`CalcTempBus]          temp_b1_5_26_i;
wire signed [`CalcTempBus]          temp_b1_5_27_r;
wire signed [`CalcTempBus]          temp_b1_5_27_i;
wire signed [`CalcTempBus]          temp_b1_5_28_r;
wire signed [`CalcTempBus]          temp_b1_5_28_i;
wire signed [`CalcTempBus]          temp_b1_5_29_r;
wire signed [`CalcTempBus]          temp_b1_5_29_i;
wire signed [`CalcTempBus]          temp_b1_5_30_r;
wire signed [`CalcTempBus]          temp_b1_5_30_i;
wire signed [`CalcTempBus]          temp_b1_5_31_r;
wire signed [`CalcTempBus]          temp_b1_5_31_i;
wire signed [`CalcTempBus]          temp_b1_5_32_r;
wire signed [`CalcTempBus]          temp_b1_5_32_i;
wire signed [`CalcTempBus]          temp_b1_6_1_r;
wire signed [`CalcTempBus]          temp_b1_6_1_i;
wire signed [`CalcTempBus]          temp_b1_6_2_r;
wire signed [`CalcTempBus]          temp_b1_6_2_i;
wire signed [`CalcTempBus]          temp_b1_6_3_r;
wire signed [`CalcTempBus]          temp_b1_6_3_i;
wire signed [`CalcTempBus]          temp_b1_6_4_r;
wire signed [`CalcTempBus]          temp_b1_6_4_i;
wire signed [`CalcTempBus]          temp_b1_6_5_r;
wire signed [`CalcTempBus]          temp_b1_6_5_i;
wire signed [`CalcTempBus]          temp_b1_6_6_r;
wire signed [`CalcTempBus]          temp_b1_6_6_i;
wire signed [`CalcTempBus]          temp_b1_6_7_r;
wire signed [`CalcTempBus]          temp_b1_6_7_i;
wire signed [`CalcTempBus]          temp_b1_6_8_r;
wire signed [`CalcTempBus]          temp_b1_6_8_i;
wire signed [`CalcTempBus]          temp_b1_6_9_r;
wire signed [`CalcTempBus]          temp_b1_6_9_i;
wire signed [`CalcTempBus]          temp_b1_6_10_r;
wire signed [`CalcTempBus]          temp_b1_6_10_i;
wire signed [`CalcTempBus]          temp_b1_6_11_r;
wire signed [`CalcTempBus]          temp_b1_6_11_i;
wire signed [`CalcTempBus]          temp_b1_6_12_r;
wire signed [`CalcTempBus]          temp_b1_6_12_i;
wire signed [`CalcTempBus]          temp_b1_6_13_r;
wire signed [`CalcTempBus]          temp_b1_6_13_i;
wire signed [`CalcTempBus]          temp_b1_6_14_r;
wire signed [`CalcTempBus]          temp_b1_6_14_i;
wire signed [`CalcTempBus]          temp_b1_6_15_r;
wire signed [`CalcTempBus]          temp_b1_6_15_i;
wire signed [`CalcTempBus]          temp_b1_6_16_r;
wire signed [`CalcTempBus]          temp_b1_6_16_i;
wire signed [`CalcTempBus]          temp_b1_6_17_r;
wire signed [`CalcTempBus]          temp_b1_6_17_i;
wire signed [`CalcTempBus]          temp_b1_6_18_r;
wire signed [`CalcTempBus]          temp_b1_6_18_i;
wire signed [`CalcTempBus]          temp_b1_6_19_r;
wire signed [`CalcTempBus]          temp_b1_6_19_i;
wire signed [`CalcTempBus]          temp_b1_6_20_r;
wire signed [`CalcTempBus]          temp_b1_6_20_i;
wire signed [`CalcTempBus]          temp_b1_6_21_r;
wire signed [`CalcTempBus]          temp_b1_6_21_i;
wire signed [`CalcTempBus]          temp_b1_6_22_r;
wire signed [`CalcTempBus]          temp_b1_6_22_i;
wire signed [`CalcTempBus]          temp_b1_6_23_r;
wire signed [`CalcTempBus]          temp_b1_6_23_i;
wire signed [`CalcTempBus]          temp_b1_6_24_r;
wire signed [`CalcTempBus]          temp_b1_6_24_i;
wire signed [`CalcTempBus]          temp_b1_6_25_r;
wire signed [`CalcTempBus]          temp_b1_6_25_i;
wire signed [`CalcTempBus]          temp_b1_6_26_r;
wire signed [`CalcTempBus]          temp_b1_6_26_i;
wire signed [`CalcTempBus]          temp_b1_6_27_r;
wire signed [`CalcTempBus]          temp_b1_6_27_i;
wire signed [`CalcTempBus]          temp_b1_6_28_r;
wire signed [`CalcTempBus]          temp_b1_6_28_i;
wire signed [`CalcTempBus]          temp_b1_6_29_r;
wire signed [`CalcTempBus]          temp_b1_6_29_i;
wire signed [`CalcTempBus]          temp_b1_6_30_r;
wire signed [`CalcTempBus]          temp_b1_6_30_i;
wire signed [`CalcTempBus]          temp_b1_6_31_r;
wire signed [`CalcTempBus]          temp_b1_6_31_i;
wire signed [`CalcTempBus]          temp_b1_6_32_r;
wire signed [`CalcTempBus]          temp_b1_6_32_i;
wire signed [`CalcTempBus]          temp_b1_7_1_r;
wire signed [`CalcTempBus]          temp_b1_7_1_i;
wire signed [`CalcTempBus]          temp_b1_7_2_r;
wire signed [`CalcTempBus]          temp_b1_7_2_i;
wire signed [`CalcTempBus]          temp_b1_7_3_r;
wire signed [`CalcTempBus]          temp_b1_7_3_i;
wire signed [`CalcTempBus]          temp_b1_7_4_r;
wire signed [`CalcTempBus]          temp_b1_7_4_i;
wire signed [`CalcTempBus]          temp_b1_7_5_r;
wire signed [`CalcTempBus]          temp_b1_7_5_i;
wire signed [`CalcTempBus]          temp_b1_7_6_r;
wire signed [`CalcTempBus]          temp_b1_7_6_i;
wire signed [`CalcTempBus]          temp_b1_7_7_r;
wire signed [`CalcTempBus]          temp_b1_7_7_i;
wire signed [`CalcTempBus]          temp_b1_7_8_r;
wire signed [`CalcTempBus]          temp_b1_7_8_i;
wire signed [`CalcTempBus]          temp_b1_7_9_r;
wire signed [`CalcTempBus]          temp_b1_7_9_i;
wire signed [`CalcTempBus]          temp_b1_7_10_r;
wire signed [`CalcTempBus]          temp_b1_7_10_i;
wire signed [`CalcTempBus]          temp_b1_7_11_r;
wire signed [`CalcTempBus]          temp_b1_7_11_i;
wire signed [`CalcTempBus]          temp_b1_7_12_r;
wire signed [`CalcTempBus]          temp_b1_7_12_i;
wire signed [`CalcTempBus]          temp_b1_7_13_r;
wire signed [`CalcTempBus]          temp_b1_7_13_i;
wire signed [`CalcTempBus]          temp_b1_7_14_r;
wire signed [`CalcTempBus]          temp_b1_7_14_i;
wire signed [`CalcTempBus]          temp_b1_7_15_r;
wire signed [`CalcTempBus]          temp_b1_7_15_i;
wire signed [`CalcTempBus]          temp_b1_7_16_r;
wire signed [`CalcTempBus]          temp_b1_7_16_i;
wire signed [`CalcTempBus]          temp_b1_7_17_r;
wire signed [`CalcTempBus]          temp_b1_7_17_i;
wire signed [`CalcTempBus]          temp_b1_7_18_r;
wire signed [`CalcTempBus]          temp_b1_7_18_i;
wire signed [`CalcTempBus]          temp_b1_7_19_r;
wire signed [`CalcTempBus]          temp_b1_7_19_i;
wire signed [`CalcTempBus]          temp_b1_7_20_r;
wire signed [`CalcTempBus]          temp_b1_7_20_i;
wire signed [`CalcTempBus]          temp_b1_7_21_r;
wire signed [`CalcTempBus]          temp_b1_7_21_i;
wire signed [`CalcTempBus]          temp_b1_7_22_r;
wire signed [`CalcTempBus]          temp_b1_7_22_i;
wire signed [`CalcTempBus]          temp_b1_7_23_r;
wire signed [`CalcTempBus]          temp_b1_7_23_i;
wire signed [`CalcTempBus]          temp_b1_7_24_r;
wire signed [`CalcTempBus]          temp_b1_7_24_i;
wire signed [`CalcTempBus]          temp_b1_7_25_r;
wire signed [`CalcTempBus]          temp_b1_7_25_i;
wire signed [`CalcTempBus]          temp_b1_7_26_r;
wire signed [`CalcTempBus]          temp_b1_7_26_i;
wire signed [`CalcTempBus]          temp_b1_7_27_r;
wire signed [`CalcTempBus]          temp_b1_7_27_i;
wire signed [`CalcTempBus]          temp_b1_7_28_r;
wire signed [`CalcTempBus]          temp_b1_7_28_i;
wire signed [`CalcTempBus]          temp_b1_7_29_r;
wire signed [`CalcTempBus]          temp_b1_7_29_i;
wire signed [`CalcTempBus]          temp_b1_7_30_r;
wire signed [`CalcTempBus]          temp_b1_7_30_i;
wire signed [`CalcTempBus]          temp_b1_7_31_r;
wire signed [`CalcTempBus]          temp_b1_7_31_i;
wire signed [`CalcTempBus]          temp_b1_7_32_r;
wire signed [`CalcTempBus]          temp_b1_7_32_i;
wire signed [`CalcTempBus]          temp_b1_8_1_r;
wire signed [`CalcTempBus]          temp_b1_8_1_i;
wire signed [`CalcTempBus]          temp_b1_8_2_r;
wire signed [`CalcTempBus]          temp_b1_8_2_i;
wire signed [`CalcTempBus]          temp_b1_8_3_r;
wire signed [`CalcTempBus]          temp_b1_8_3_i;
wire signed [`CalcTempBus]          temp_b1_8_4_r;
wire signed [`CalcTempBus]          temp_b1_8_4_i;
wire signed [`CalcTempBus]          temp_b1_8_5_r;
wire signed [`CalcTempBus]          temp_b1_8_5_i;
wire signed [`CalcTempBus]          temp_b1_8_6_r;
wire signed [`CalcTempBus]          temp_b1_8_6_i;
wire signed [`CalcTempBus]          temp_b1_8_7_r;
wire signed [`CalcTempBus]          temp_b1_8_7_i;
wire signed [`CalcTempBus]          temp_b1_8_8_r;
wire signed [`CalcTempBus]          temp_b1_8_8_i;
wire signed [`CalcTempBus]          temp_b1_8_9_r;
wire signed [`CalcTempBus]          temp_b1_8_9_i;
wire signed [`CalcTempBus]          temp_b1_8_10_r;
wire signed [`CalcTempBus]          temp_b1_8_10_i;
wire signed [`CalcTempBus]          temp_b1_8_11_r;
wire signed [`CalcTempBus]          temp_b1_8_11_i;
wire signed [`CalcTempBus]          temp_b1_8_12_r;
wire signed [`CalcTempBus]          temp_b1_8_12_i;
wire signed [`CalcTempBus]          temp_b1_8_13_r;
wire signed [`CalcTempBus]          temp_b1_8_13_i;
wire signed [`CalcTempBus]          temp_b1_8_14_r;
wire signed [`CalcTempBus]          temp_b1_8_14_i;
wire signed [`CalcTempBus]          temp_b1_8_15_r;
wire signed [`CalcTempBus]          temp_b1_8_15_i;
wire signed [`CalcTempBus]          temp_b1_8_16_r;
wire signed [`CalcTempBus]          temp_b1_8_16_i;
wire signed [`CalcTempBus]          temp_b1_8_17_r;
wire signed [`CalcTempBus]          temp_b1_8_17_i;
wire signed [`CalcTempBus]          temp_b1_8_18_r;
wire signed [`CalcTempBus]          temp_b1_8_18_i;
wire signed [`CalcTempBus]          temp_b1_8_19_r;
wire signed [`CalcTempBus]          temp_b1_8_19_i;
wire signed [`CalcTempBus]          temp_b1_8_20_r;
wire signed [`CalcTempBus]          temp_b1_8_20_i;
wire signed [`CalcTempBus]          temp_b1_8_21_r;
wire signed [`CalcTempBus]          temp_b1_8_21_i;
wire signed [`CalcTempBus]          temp_b1_8_22_r;
wire signed [`CalcTempBus]          temp_b1_8_22_i;
wire signed [`CalcTempBus]          temp_b1_8_23_r;
wire signed [`CalcTempBus]          temp_b1_8_23_i;
wire signed [`CalcTempBus]          temp_b1_8_24_r;
wire signed [`CalcTempBus]          temp_b1_8_24_i;
wire signed [`CalcTempBus]          temp_b1_8_25_r;
wire signed [`CalcTempBus]          temp_b1_8_25_i;
wire signed [`CalcTempBus]          temp_b1_8_26_r;
wire signed [`CalcTempBus]          temp_b1_8_26_i;
wire signed [`CalcTempBus]          temp_b1_8_27_r;
wire signed [`CalcTempBus]          temp_b1_8_27_i;
wire signed [`CalcTempBus]          temp_b1_8_28_r;
wire signed [`CalcTempBus]          temp_b1_8_28_i;
wire signed [`CalcTempBus]          temp_b1_8_29_r;
wire signed [`CalcTempBus]          temp_b1_8_29_i;
wire signed [`CalcTempBus]          temp_b1_8_30_r;
wire signed [`CalcTempBus]          temp_b1_8_30_i;
wire signed [`CalcTempBus]          temp_b1_8_31_r;
wire signed [`CalcTempBus]          temp_b1_8_31_i;
wire signed [`CalcTempBus]          temp_b1_8_32_r;
wire signed [`CalcTempBus]          temp_b1_8_32_i;
wire signed [`CalcTempBus]          temp_b1_9_1_r;
wire signed [`CalcTempBus]          temp_b1_9_1_i;
wire signed [`CalcTempBus]          temp_b1_9_2_r;
wire signed [`CalcTempBus]          temp_b1_9_2_i;
wire signed [`CalcTempBus]          temp_b1_9_3_r;
wire signed [`CalcTempBus]          temp_b1_9_3_i;
wire signed [`CalcTempBus]          temp_b1_9_4_r;
wire signed [`CalcTempBus]          temp_b1_9_4_i;
wire signed [`CalcTempBus]          temp_b1_9_5_r;
wire signed [`CalcTempBus]          temp_b1_9_5_i;
wire signed [`CalcTempBus]          temp_b1_9_6_r;
wire signed [`CalcTempBus]          temp_b1_9_6_i;
wire signed [`CalcTempBus]          temp_b1_9_7_r;
wire signed [`CalcTempBus]          temp_b1_9_7_i;
wire signed [`CalcTempBus]          temp_b1_9_8_r;
wire signed [`CalcTempBus]          temp_b1_9_8_i;
wire signed [`CalcTempBus]          temp_b1_9_9_r;
wire signed [`CalcTempBus]          temp_b1_9_9_i;
wire signed [`CalcTempBus]          temp_b1_9_10_r;
wire signed [`CalcTempBus]          temp_b1_9_10_i;
wire signed [`CalcTempBus]          temp_b1_9_11_r;
wire signed [`CalcTempBus]          temp_b1_9_11_i;
wire signed [`CalcTempBus]          temp_b1_9_12_r;
wire signed [`CalcTempBus]          temp_b1_9_12_i;
wire signed [`CalcTempBus]          temp_b1_9_13_r;
wire signed [`CalcTempBus]          temp_b1_9_13_i;
wire signed [`CalcTempBus]          temp_b1_9_14_r;
wire signed [`CalcTempBus]          temp_b1_9_14_i;
wire signed [`CalcTempBus]          temp_b1_9_15_r;
wire signed [`CalcTempBus]          temp_b1_9_15_i;
wire signed [`CalcTempBus]          temp_b1_9_16_r;
wire signed [`CalcTempBus]          temp_b1_9_16_i;
wire signed [`CalcTempBus]          temp_b1_9_17_r;
wire signed [`CalcTempBus]          temp_b1_9_17_i;
wire signed [`CalcTempBus]          temp_b1_9_18_r;
wire signed [`CalcTempBus]          temp_b1_9_18_i;
wire signed [`CalcTempBus]          temp_b1_9_19_r;
wire signed [`CalcTempBus]          temp_b1_9_19_i;
wire signed [`CalcTempBus]          temp_b1_9_20_r;
wire signed [`CalcTempBus]          temp_b1_9_20_i;
wire signed [`CalcTempBus]          temp_b1_9_21_r;
wire signed [`CalcTempBus]          temp_b1_9_21_i;
wire signed [`CalcTempBus]          temp_b1_9_22_r;
wire signed [`CalcTempBus]          temp_b1_9_22_i;
wire signed [`CalcTempBus]          temp_b1_9_23_r;
wire signed [`CalcTempBus]          temp_b1_9_23_i;
wire signed [`CalcTempBus]          temp_b1_9_24_r;
wire signed [`CalcTempBus]          temp_b1_9_24_i;
wire signed [`CalcTempBus]          temp_b1_9_25_r;
wire signed [`CalcTempBus]          temp_b1_9_25_i;
wire signed [`CalcTempBus]          temp_b1_9_26_r;
wire signed [`CalcTempBus]          temp_b1_9_26_i;
wire signed [`CalcTempBus]          temp_b1_9_27_r;
wire signed [`CalcTempBus]          temp_b1_9_27_i;
wire signed [`CalcTempBus]          temp_b1_9_28_r;
wire signed [`CalcTempBus]          temp_b1_9_28_i;
wire signed [`CalcTempBus]          temp_b1_9_29_r;
wire signed [`CalcTempBus]          temp_b1_9_29_i;
wire signed [`CalcTempBus]          temp_b1_9_30_r;
wire signed [`CalcTempBus]          temp_b1_9_30_i;
wire signed [`CalcTempBus]          temp_b1_9_31_r;
wire signed [`CalcTempBus]          temp_b1_9_31_i;
wire signed [`CalcTempBus]          temp_b1_9_32_r;
wire signed [`CalcTempBus]          temp_b1_9_32_i;
wire signed [`CalcTempBus]          temp_b1_10_1_r;
wire signed [`CalcTempBus]          temp_b1_10_1_i;
wire signed [`CalcTempBus]          temp_b1_10_2_r;
wire signed [`CalcTempBus]          temp_b1_10_2_i;
wire signed [`CalcTempBus]          temp_b1_10_3_r;
wire signed [`CalcTempBus]          temp_b1_10_3_i;
wire signed [`CalcTempBus]          temp_b1_10_4_r;
wire signed [`CalcTempBus]          temp_b1_10_4_i;
wire signed [`CalcTempBus]          temp_b1_10_5_r;
wire signed [`CalcTempBus]          temp_b1_10_5_i;
wire signed [`CalcTempBus]          temp_b1_10_6_r;
wire signed [`CalcTempBus]          temp_b1_10_6_i;
wire signed [`CalcTempBus]          temp_b1_10_7_r;
wire signed [`CalcTempBus]          temp_b1_10_7_i;
wire signed [`CalcTempBus]          temp_b1_10_8_r;
wire signed [`CalcTempBus]          temp_b1_10_8_i;
wire signed [`CalcTempBus]          temp_b1_10_9_r;
wire signed [`CalcTempBus]          temp_b1_10_9_i;
wire signed [`CalcTempBus]          temp_b1_10_10_r;
wire signed [`CalcTempBus]          temp_b1_10_10_i;
wire signed [`CalcTempBus]          temp_b1_10_11_r;
wire signed [`CalcTempBus]          temp_b1_10_11_i;
wire signed [`CalcTempBus]          temp_b1_10_12_r;
wire signed [`CalcTempBus]          temp_b1_10_12_i;
wire signed [`CalcTempBus]          temp_b1_10_13_r;
wire signed [`CalcTempBus]          temp_b1_10_13_i;
wire signed [`CalcTempBus]          temp_b1_10_14_r;
wire signed [`CalcTempBus]          temp_b1_10_14_i;
wire signed [`CalcTempBus]          temp_b1_10_15_r;
wire signed [`CalcTempBus]          temp_b1_10_15_i;
wire signed [`CalcTempBus]          temp_b1_10_16_r;
wire signed [`CalcTempBus]          temp_b1_10_16_i;
wire signed [`CalcTempBus]          temp_b1_10_17_r;
wire signed [`CalcTempBus]          temp_b1_10_17_i;
wire signed [`CalcTempBus]          temp_b1_10_18_r;
wire signed [`CalcTempBus]          temp_b1_10_18_i;
wire signed [`CalcTempBus]          temp_b1_10_19_r;
wire signed [`CalcTempBus]          temp_b1_10_19_i;
wire signed [`CalcTempBus]          temp_b1_10_20_r;
wire signed [`CalcTempBus]          temp_b1_10_20_i;
wire signed [`CalcTempBus]          temp_b1_10_21_r;
wire signed [`CalcTempBus]          temp_b1_10_21_i;
wire signed [`CalcTempBus]          temp_b1_10_22_r;
wire signed [`CalcTempBus]          temp_b1_10_22_i;
wire signed [`CalcTempBus]          temp_b1_10_23_r;
wire signed [`CalcTempBus]          temp_b1_10_23_i;
wire signed [`CalcTempBus]          temp_b1_10_24_r;
wire signed [`CalcTempBus]          temp_b1_10_24_i;
wire signed [`CalcTempBus]          temp_b1_10_25_r;
wire signed [`CalcTempBus]          temp_b1_10_25_i;
wire signed [`CalcTempBus]          temp_b1_10_26_r;
wire signed [`CalcTempBus]          temp_b1_10_26_i;
wire signed [`CalcTempBus]          temp_b1_10_27_r;
wire signed [`CalcTempBus]          temp_b1_10_27_i;
wire signed [`CalcTempBus]          temp_b1_10_28_r;
wire signed [`CalcTempBus]          temp_b1_10_28_i;
wire signed [`CalcTempBus]          temp_b1_10_29_r;
wire signed [`CalcTempBus]          temp_b1_10_29_i;
wire signed [`CalcTempBus]          temp_b1_10_30_r;
wire signed [`CalcTempBus]          temp_b1_10_30_i;
wire signed [`CalcTempBus]          temp_b1_10_31_r;
wire signed [`CalcTempBus]          temp_b1_10_31_i;
wire signed [`CalcTempBus]          temp_b1_10_32_r;
wire signed [`CalcTempBus]          temp_b1_10_32_i;
wire signed [`CalcTempBus]          temp_b1_11_1_r;
wire signed [`CalcTempBus]          temp_b1_11_1_i;
wire signed [`CalcTempBus]          temp_b1_11_2_r;
wire signed [`CalcTempBus]          temp_b1_11_2_i;
wire signed [`CalcTempBus]          temp_b1_11_3_r;
wire signed [`CalcTempBus]          temp_b1_11_3_i;
wire signed [`CalcTempBus]          temp_b1_11_4_r;
wire signed [`CalcTempBus]          temp_b1_11_4_i;
wire signed [`CalcTempBus]          temp_b1_11_5_r;
wire signed [`CalcTempBus]          temp_b1_11_5_i;
wire signed [`CalcTempBus]          temp_b1_11_6_r;
wire signed [`CalcTempBus]          temp_b1_11_6_i;
wire signed [`CalcTempBus]          temp_b1_11_7_r;
wire signed [`CalcTempBus]          temp_b1_11_7_i;
wire signed [`CalcTempBus]          temp_b1_11_8_r;
wire signed [`CalcTempBus]          temp_b1_11_8_i;
wire signed [`CalcTempBus]          temp_b1_11_9_r;
wire signed [`CalcTempBus]          temp_b1_11_9_i;
wire signed [`CalcTempBus]          temp_b1_11_10_r;
wire signed [`CalcTempBus]          temp_b1_11_10_i;
wire signed [`CalcTempBus]          temp_b1_11_11_r;
wire signed [`CalcTempBus]          temp_b1_11_11_i;
wire signed [`CalcTempBus]          temp_b1_11_12_r;
wire signed [`CalcTempBus]          temp_b1_11_12_i;
wire signed [`CalcTempBus]          temp_b1_11_13_r;
wire signed [`CalcTempBus]          temp_b1_11_13_i;
wire signed [`CalcTempBus]          temp_b1_11_14_r;
wire signed [`CalcTempBus]          temp_b1_11_14_i;
wire signed [`CalcTempBus]          temp_b1_11_15_r;
wire signed [`CalcTempBus]          temp_b1_11_15_i;
wire signed [`CalcTempBus]          temp_b1_11_16_r;
wire signed [`CalcTempBus]          temp_b1_11_16_i;
wire signed [`CalcTempBus]          temp_b1_11_17_r;
wire signed [`CalcTempBus]          temp_b1_11_17_i;
wire signed [`CalcTempBus]          temp_b1_11_18_r;
wire signed [`CalcTempBus]          temp_b1_11_18_i;
wire signed [`CalcTempBus]          temp_b1_11_19_r;
wire signed [`CalcTempBus]          temp_b1_11_19_i;
wire signed [`CalcTempBus]          temp_b1_11_20_r;
wire signed [`CalcTempBus]          temp_b1_11_20_i;
wire signed [`CalcTempBus]          temp_b1_11_21_r;
wire signed [`CalcTempBus]          temp_b1_11_21_i;
wire signed [`CalcTempBus]          temp_b1_11_22_r;
wire signed [`CalcTempBus]          temp_b1_11_22_i;
wire signed [`CalcTempBus]          temp_b1_11_23_r;
wire signed [`CalcTempBus]          temp_b1_11_23_i;
wire signed [`CalcTempBus]          temp_b1_11_24_r;
wire signed [`CalcTempBus]          temp_b1_11_24_i;
wire signed [`CalcTempBus]          temp_b1_11_25_r;
wire signed [`CalcTempBus]          temp_b1_11_25_i;
wire signed [`CalcTempBus]          temp_b1_11_26_r;
wire signed [`CalcTempBus]          temp_b1_11_26_i;
wire signed [`CalcTempBus]          temp_b1_11_27_r;
wire signed [`CalcTempBus]          temp_b1_11_27_i;
wire signed [`CalcTempBus]          temp_b1_11_28_r;
wire signed [`CalcTempBus]          temp_b1_11_28_i;
wire signed [`CalcTempBus]          temp_b1_11_29_r;
wire signed [`CalcTempBus]          temp_b1_11_29_i;
wire signed [`CalcTempBus]          temp_b1_11_30_r;
wire signed [`CalcTempBus]          temp_b1_11_30_i;
wire signed [`CalcTempBus]          temp_b1_11_31_r;
wire signed [`CalcTempBus]          temp_b1_11_31_i;
wire signed [`CalcTempBus]          temp_b1_11_32_r;
wire signed [`CalcTempBus]          temp_b1_11_32_i;
wire signed [`CalcTempBus]          temp_b1_12_1_r;
wire signed [`CalcTempBus]          temp_b1_12_1_i;
wire signed [`CalcTempBus]          temp_b1_12_2_r;
wire signed [`CalcTempBus]          temp_b1_12_2_i;
wire signed [`CalcTempBus]          temp_b1_12_3_r;
wire signed [`CalcTempBus]          temp_b1_12_3_i;
wire signed [`CalcTempBus]          temp_b1_12_4_r;
wire signed [`CalcTempBus]          temp_b1_12_4_i;
wire signed [`CalcTempBus]          temp_b1_12_5_r;
wire signed [`CalcTempBus]          temp_b1_12_5_i;
wire signed [`CalcTempBus]          temp_b1_12_6_r;
wire signed [`CalcTempBus]          temp_b1_12_6_i;
wire signed [`CalcTempBus]          temp_b1_12_7_r;
wire signed [`CalcTempBus]          temp_b1_12_7_i;
wire signed [`CalcTempBus]          temp_b1_12_8_r;
wire signed [`CalcTempBus]          temp_b1_12_8_i;
wire signed [`CalcTempBus]          temp_b1_12_9_r;
wire signed [`CalcTempBus]          temp_b1_12_9_i;
wire signed [`CalcTempBus]          temp_b1_12_10_r;
wire signed [`CalcTempBus]          temp_b1_12_10_i;
wire signed [`CalcTempBus]          temp_b1_12_11_r;
wire signed [`CalcTempBus]          temp_b1_12_11_i;
wire signed [`CalcTempBus]          temp_b1_12_12_r;
wire signed [`CalcTempBus]          temp_b1_12_12_i;
wire signed [`CalcTempBus]          temp_b1_12_13_r;
wire signed [`CalcTempBus]          temp_b1_12_13_i;
wire signed [`CalcTempBus]          temp_b1_12_14_r;
wire signed [`CalcTempBus]          temp_b1_12_14_i;
wire signed [`CalcTempBus]          temp_b1_12_15_r;
wire signed [`CalcTempBus]          temp_b1_12_15_i;
wire signed [`CalcTempBus]          temp_b1_12_16_r;
wire signed [`CalcTempBus]          temp_b1_12_16_i;
wire signed [`CalcTempBus]          temp_b1_12_17_r;
wire signed [`CalcTempBus]          temp_b1_12_17_i;
wire signed [`CalcTempBus]          temp_b1_12_18_r;
wire signed [`CalcTempBus]          temp_b1_12_18_i;
wire signed [`CalcTempBus]          temp_b1_12_19_r;
wire signed [`CalcTempBus]          temp_b1_12_19_i;
wire signed [`CalcTempBus]          temp_b1_12_20_r;
wire signed [`CalcTempBus]          temp_b1_12_20_i;
wire signed [`CalcTempBus]          temp_b1_12_21_r;
wire signed [`CalcTempBus]          temp_b1_12_21_i;
wire signed [`CalcTempBus]          temp_b1_12_22_r;
wire signed [`CalcTempBus]          temp_b1_12_22_i;
wire signed [`CalcTempBus]          temp_b1_12_23_r;
wire signed [`CalcTempBus]          temp_b1_12_23_i;
wire signed [`CalcTempBus]          temp_b1_12_24_r;
wire signed [`CalcTempBus]          temp_b1_12_24_i;
wire signed [`CalcTempBus]          temp_b1_12_25_r;
wire signed [`CalcTempBus]          temp_b1_12_25_i;
wire signed [`CalcTempBus]          temp_b1_12_26_r;
wire signed [`CalcTempBus]          temp_b1_12_26_i;
wire signed [`CalcTempBus]          temp_b1_12_27_r;
wire signed [`CalcTempBus]          temp_b1_12_27_i;
wire signed [`CalcTempBus]          temp_b1_12_28_r;
wire signed [`CalcTempBus]          temp_b1_12_28_i;
wire signed [`CalcTempBus]          temp_b1_12_29_r;
wire signed [`CalcTempBus]          temp_b1_12_29_i;
wire signed [`CalcTempBus]          temp_b1_12_30_r;
wire signed [`CalcTempBus]          temp_b1_12_30_i;
wire signed [`CalcTempBus]          temp_b1_12_31_r;
wire signed [`CalcTempBus]          temp_b1_12_31_i;
wire signed [`CalcTempBus]          temp_b1_12_32_r;
wire signed [`CalcTempBus]          temp_b1_12_32_i;
wire signed [`CalcTempBus]          temp_b1_13_1_r;
wire signed [`CalcTempBus]          temp_b1_13_1_i;
wire signed [`CalcTempBus]          temp_b1_13_2_r;
wire signed [`CalcTempBus]          temp_b1_13_2_i;
wire signed [`CalcTempBus]          temp_b1_13_3_r;
wire signed [`CalcTempBus]          temp_b1_13_3_i;
wire signed [`CalcTempBus]          temp_b1_13_4_r;
wire signed [`CalcTempBus]          temp_b1_13_4_i;
wire signed [`CalcTempBus]          temp_b1_13_5_r;
wire signed [`CalcTempBus]          temp_b1_13_5_i;
wire signed [`CalcTempBus]          temp_b1_13_6_r;
wire signed [`CalcTempBus]          temp_b1_13_6_i;
wire signed [`CalcTempBus]          temp_b1_13_7_r;
wire signed [`CalcTempBus]          temp_b1_13_7_i;
wire signed [`CalcTempBus]          temp_b1_13_8_r;
wire signed [`CalcTempBus]          temp_b1_13_8_i;
wire signed [`CalcTempBus]          temp_b1_13_9_r;
wire signed [`CalcTempBus]          temp_b1_13_9_i;
wire signed [`CalcTempBus]          temp_b1_13_10_r;
wire signed [`CalcTempBus]          temp_b1_13_10_i;
wire signed [`CalcTempBus]          temp_b1_13_11_r;
wire signed [`CalcTempBus]          temp_b1_13_11_i;
wire signed [`CalcTempBus]          temp_b1_13_12_r;
wire signed [`CalcTempBus]          temp_b1_13_12_i;
wire signed [`CalcTempBus]          temp_b1_13_13_r;
wire signed [`CalcTempBus]          temp_b1_13_13_i;
wire signed [`CalcTempBus]          temp_b1_13_14_r;
wire signed [`CalcTempBus]          temp_b1_13_14_i;
wire signed [`CalcTempBus]          temp_b1_13_15_r;
wire signed [`CalcTempBus]          temp_b1_13_15_i;
wire signed [`CalcTempBus]          temp_b1_13_16_r;
wire signed [`CalcTempBus]          temp_b1_13_16_i;
wire signed [`CalcTempBus]          temp_b1_13_17_r;
wire signed [`CalcTempBus]          temp_b1_13_17_i;
wire signed [`CalcTempBus]          temp_b1_13_18_r;
wire signed [`CalcTempBus]          temp_b1_13_18_i;
wire signed [`CalcTempBus]          temp_b1_13_19_r;
wire signed [`CalcTempBus]          temp_b1_13_19_i;
wire signed [`CalcTempBus]          temp_b1_13_20_r;
wire signed [`CalcTempBus]          temp_b1_13_20_i;
wire signed [`CalcTempBus]          temp_b1_13_21_r;
wire signed [`CalcTempBus]          temp_b1_13_21_i;
wire signed [`CalcTempBus]          temp_b1_13_22_r;
wire signed [`CalcTempBus]          temp_b1_13_22_i;
wire signed [`CalcTempBus]          temp_b1_13_23_r;
wire signed [`CalcTempBus]          temp_b1_13_23_i;
wire signed [`CalcTempBus]          temp_b1_13_24_r;
wire signed [`CalcTempBus]          temp_b1_13_24_i;
wire signed [`CalcTempBus]          temp_b1_13_25_r;
wire signed [`CalcTempBus]          temp_b1_13_25_i;
wire signed [`CalcTempBus]          temp_b1_13_26_r;
wire signed [`CalcTempBus]          temp_b1_13_26_i;
wire signed [`CalcTempBus]          temp_b1_13_27_r;
wire signed [`CalcTempBus]          temp_b1_13_27_i;
wire signed [`CalcTempBus]          temp_b1_13_28_r;
wire signed [`CalcTempBus]          temp_b1_13_28_i;
wire signed [`CalcTempBus]          temp_b1_13_29_r;
wire signed [`CalcTempBus]          temp_b1_13_29_i;
wire signed [`CalcTempBus]          temp_b1_13_30_r;
wire signed [`CalcTempBus]          temp_b1_13_30_i;
wire signed [`CalcTempBus]          temp_b1_13_31_r;
wire signed [`CalcTempBus]          temp_b1_13_31_i;
wire signed [`CalcTempBus]          temp_b1_13_32_r;
wire signed [`CalcTempBus]          temp_b1_13_32_i;
wire signed [`CalcTempBus]          temp_b1_14_1_r;
wire signed [`CalcTempBus]          temp_b1_14_1_i;
wire signed [`CalcTempBus]          temp_b1_14_2_r;
wire signed [`CalcTempBus]          temp_b1_14_2_i;
wire signed [`CalcTempBus]          temp_b1_14_3_r;
wire signed [`CalcTempBus]          temp_b1_14_3_i;
wire signed [`CalcTempBus]          temp_b1_14_4_r;
wire signed [`CalcTempBus]          temp_b1_14_4_i;
wire signed [`CalcTempBus]          temp_b1_14_5_r;
wire signed [`CalcTempBus]          temp_b1_14_5_i;
wire signed [`CalcTempBus]          temp_b1_14_6_r;
wire signed [`CalcTempBus]          temp_b1_14_6_i;
wire signed [`CalcTempBus]          temp_b1_14_7_r;
wire signed [`CalcTempBus]          temp_b1_14_7_i;
wire signed [`CalcTempBus]          temp_b1_14_8_r;
wire signed [`CalcTempBus]          temp_b1_14_8_i;
wire signed [`CalcTempBus]          temp_b1_14_9_r;
wire signed [`CalcTempBus]          temp_b1_14_9_i;
wire signed [`CalcTempBus]          temp_b1_14_10_r;
wire signed [`CalcTempBus]          temp_b1_14_10_i;
wire signed [`CalcTempBus]          temp_b1_14_11_r;
wire signed [`CalcTempBus]          temp_b1_14_11_i;
wire signed [`CalcTempBus]          temp_b1_14_12_r;
wire signed [`CalcTempBus]          temp_b1_14_12_i;
wire signed [`CalcTempBus]          temp_b1_14_13_r;
wire signed [`CalcTempBus]          temp_b1_14_13_i;
wire signed [`CalcTempBus]          temp_b1_14_14_r;
wire signed [`CalcTempBus]          temp_b1_14_14_i;
wire signed [`CalcTempBus]          temp_b1_14_15_r;
wire signed [`CalcTempBus]          temp_b1_14_15_i;
wire signed [`CalcTempBus]          temp_b1_14_16_r;
wire signed [`CalcTempBus]          temp_b1_14_16_i;
wire signed [`CalcTempBus]          temp_b1_14_17_r;
wire signed [`CalcTempBus]          temp_b1_14_17_i;
wire signed [`CalcTempBus]          temp_b1_14_18_r;
wire signed [`CalcTempBus]          temp_b1_14_18_i;
wire signed [`CalcTempBus]          temp_b1_14_19_r;
wire signed [`CalcTempBus]          temp_b1_14_19_i;
wire signed [`CalcTempBus]          temp_b1_14_20_r;
wire signed [`CalcTempBus]          temp_b1_14_20_i;
wire signed [`CalcTempBus]          temp_b1_14_21_r;
wire signed [`CalcTempBus]          temp_b1_14_21_i;
wire signed [`CalcTempBus]          temp_b1_14_22_r;
wire signed [`CalcTempBus]          temp_b1_14_22_i;
wire signed [`CalcTempBus]          temp_b1_14_23_r;
wire signed [`CalcTempBus]          temp_b1_14_23_i;
wire signed [`CalcTempBus]          temp_b1_14_24_r;
wire signed [`CalcTempBus]          temp_b1_14_24_i;
wire signed [`CalcTempBus]          temp_b1_14_25_r;
wire signed [`CalcTempBus]          temp_b1_14_25_i;
wire signed [`CalcTempBus]          temp_b1_14_26_r;
wire signed [`CalcTempBus]          temp_b1_14_26_i;
wire signed [`CalcTempBus]          temp_b1_14_27_r;
wire signed [`CalcTempBus]          temp_b1_14_27_i;
wire signed [`CalcTempBus]          temp_b1_14_28_r;
wire signed [`CalcTempBus]          temp_b1_14_28_i;
wire signed [`CalcTempBus]          temp_b1_14_29_r;
wire signed [`CalcTempBus]          temp_b1_14_29_i;
wire signed [`CalcTempBus]          temp_b1_14_30_r;
wire signed [`CalcTempBus]          temp_b1_14_30_i;
wire signed [`CalcTempBus]          temp_b1_14_31_r;
wire signed [`CalcTempBus]          temp_b1_14_31_i;
wire signed [`CalcTempBus]          temp_b1_14_32_r;
wire signed [`CalcTempBus]          temp_b1_14_32_i;
wire signed [`CalcTempBus]          temp_b1_15_1_r;
wire signed [`CalcTempBus]          temp_b1_15_1_i;
wire signed [`CalcTempBus]          temp_b1_15_2_r;
wire signed [`CalcTempBus]          temp_b1_15_2_i;
wire signed [`CalcTempBus]          temp_b1_15_3_r;
wire signed [`CalcTempBus]          temp_b1_15_3_i;
wire signed [`CalcTempBus]          temp_b1_15_4_r;
wire signed [`CalcTempBus]          temp_b1_15_4_i;
wire signed [`CalcTempBus]          temp_b1_15_5_r;
wire signed [`CalcTempBus]          temp_b1_15_5_i;
wire signed [`CalcTempBus]          temp_b1_15_6_r;
wire signed [`CalcTempBus]          temp_b1_15_6_i;
wire signed [`CalcTempBus]          temp_b1_15_7_r;
wire signed [`CalcTempBus]          temp_b1_15_7_i;
wire signed [`CalcTempBus]          temp_b1_15_8_r;
wire signed [`CalcTempBus]          temp_b1_15_8_i;
wire signed [`CalcTempBus]          temp_b1_15_9_r;
wire signed [`CalcTempBus]          temp_b1_15_9_i;
wire signed [`CalcTempBus]          temp_b1_15_10_r;
wire signed [`CalcTempBus]          temp_b1_15_10_i;
wire signed [`CalcTempBus]          temp_b1_15_11_r;
wire signed [`CalcTempBus]          temp_b1_15_11_i;
wire signed [`CalcTempBus]          temp_b1_15_12_r;
wire signed [`CalcTempBus]          temp_b1_15_12_i;
wire signed [`CalcTempBus]          temp_b1_15_13_r;
wire signed [`CalcTempBus]          temp_b1_15_13_i;
wire signed [`CalcTempBus]          temp_b1_15_14_r;
wire signed [`CalcTempBus]          temp_b1_15_14_i;
wire signed [`CalcTempBus]          temp_b1_15_15_r;
wire signed [`CalcTempBus]          temp_b1_15_15_i;
wire signed [`CalcTempBus]          temp_b1_15_16_r;
wire signed [`CalcTempBus]          temp_b1_15_16_i;
wire signed [`CalcTempBus]          temp_b1_15_17_r;
wire signed [`CalcTempBus]          temp_b1_15_17_i;
wire signed [`CalcTempBus]          temp_b1_15_18_r;
wire signed [`CalcTempBus]          temp_b1_15_18_i;
wire signed [`CalcTempBus]          temp_b1_15_19_r;
wire signed [`CalcTempBus]          temp_b1_15_19_i;
wire signed [`CalcTempBus]          temp_b1_15_20_r;
wire signed [`CalcTempBus]          temp_b1_15_20_i;
wire signed [`CalcTempBus]          temp_b1_15_21_r;
wire signed [`CalcTempBus]          temp_b1_15_21_i;
wire signed [`CalcTempBus]          temp_b1_15_22_r;
wire signed [`CalcTempBus]          temp_b1_15_22_i;
wire signed [`CalcTempBus]          temp_b1_15_23_r;
wire signed [`CalcTempBus]          temp_b1_15_23_i;
wire signed [`CalcTempBus]          temp_b1_15_24_r;
wire signed [`CalcTempBus]          temp_b1_15_24_i;
wire signed [`CalcTempBus]          temp_b1_15_25_r;
wire signed [`CalcTempBus]          temp_b1_15_25_i;
wire signed [`CalcTempBus]          temp_b1_15_26_r;
wire signed [`CalcTempBus]          temp_b1_15_26_i;
wire signed [`CalcTempBus]          temp_b1_15_27_r;
wire signed [`CalcTempBus]          temp_b1_15_27_i;
wire signed [`CalcTempBus]          temp_b1_15_28_r;
wire signed [`CalcTempBus]          temp_b1_15_28_i;
wire signed [`CalcTempBus]          temp_b1_15_29_r;
wire signed [`CalcTempBus]          temp_b1_15_29_i;
wire signed [`CalcTempBus]          temp_b1_15_30_r;
wire signed [`CalcTempBus]          temp_b1_15_30_i;
wire signed [`CalcTempBus]          temp_b1_15_31_r;
wire signed [`CalcTempBus]          temp_b1_15_31_i;
wire signed [`CalcTempBus]          temp_b1_15_32_r;
wire signed [`CalcTempBus]          temp_b1_15_32_i;
wire signed [`CalcTempBus]          temp_b1_16_1_r;
wire signed [`CalcTempBus]          temp_b1_16_1_i;
wire signed [`CalcTempBus]          temp_b1_16_2_r;
wire signed [`CalcTempBus]          temp_b1_16_2_i;
wire signed [`CalcTempBus]          temp_b1_16_3_r;
wire signed [`CalcTempBus]          temp_b1_16_3_i;
wire signed [`CalcTempBus]          temp_b1_16_4_r;
wire signed [`CalcTempBus]          temp_b1_16_4_i;
wire signed [`CalcTempBus]          temp_b1_16_5_r;
wire signed [`CalcTempBus]          temp_b1_16_5_i;
wire signed [`CalcTempBus]          temp_b1_16_6_r;
wire signed [`CalcTempBus]          temp_b1_16_6_i;
wire signed [`CalcTempBus]          temp_b1_16_7_r;
wire signed [`CalcTempBus]          temp_b1_16_7_i;
wire signed [`CalcTempBus]          temp_b1_16_8_r;
wire signed [`CalcTempBus]          temp_b1_16_8_i;
wire signed [`CalcTempBus]          temp_b1_16_9_r;
wire signed [`CalcTempBus]          temp_b1_16_9_i;
wire signed [`CalcTempBus]          temp_b1_16_10_r;
wire signed [`CalcTempBus]          temp_b1_16_10_i;
wire signed [`CalcTempBus]          temp_b1_16_11_r;
wire signed [`CalcTempBus]          temp_b1_16_11_i;
wire signed [`CalcTempBus]          temp_b1_16_12_r;
wire signed [`CalcTempBus]          temp_b1_16_12_i;
wire signed [`CalcTempBus]          temp_b1_16_13_r;
wire signed [`CalcTempBus]          temp_b1_16_13_i;
wire signed [`CalcTempBus]          temp_b1_16_14_r;
wire signed [`CalcTempBus]          temp_b1_16_14_i;
wire signed [`CalcTempBus]          temp_b1_16_15_r;
wire signed [`CalcTempBus]          temp_b1_16_15_i;
wire signed [`CalcTempBus]          temp_b1_16_16_r;
wire signed [`CalcTempBus]          temp_b1_16_16_i;
wire signed [`CalcTempBus]          temp_b1_16_17_r;
wire signed [`CalcTempBus]          temp_b1_16_17_i;
wire signed [`CalcTempBus]          temp_b1_16_18_r;
wire signed [`CalcTempBus]          temp_b1_16_18_i;
wire signed [`CalcTempBus]          temp_b1_16_19_r;
wire signed [`CalcTempBus]          temp_b1_16_19_i;
wire signed [`CalcTempBus]          temp_b1_16_20_r;
wire signed [`CalcTempBus]          temp_b1_16_20_i;
wire signed [`CalcTempBus]          temp_b1_16_21_r;
wire signed [`CalcTempBus]          temp_b1_16_21_i;
wire signed [`CalcTempBus]          temp_b1_16_22_r;
wire signed [`CalcTempBus]          temp_b1_16_22_i;
wire signed [`CalcTempBus]          temp_b1_16_23_r;
wire signed [`CalcTempBus]          temp_b1_16_23_i;
wire signed [`CalcTempBus]          temp_b1_16_24_r;
wire signed [`CalcTempBus]          temp_b1_16_24_i;
wire signed [`CalcTempBus]          temp_b1_16_25_r;
wire signed [`CalcTempBus]          temp_b1_16_25_i;
wire signed [`CalcTempBus]          temp_b1_16_26_r;
wire signed [`CalcTempBus]          temp_b1_16_26_i;
wire signed [`CalcTempBus]          temp_b1_16_27_r;
wire signed [`CalcTempBus]          temp_b1_16_27_i;
wire signed [`CalcTempBus]          temp_b1_16_28_r;
wire signed [`CalcTempBus]          temp_b1_16_28_i;
wire signed [`CalcTempBus]          temp_b1_16_29_r;
wire signed [`CalcTempBus]          temp_b1_16_29_i;
wire signed [`CalcTempBus]          temp_b1_16_30_r;
wire signed [`CalcTempBus]          temp_b1_16_30_i;
wire signed [`CalcTempBus]          temp_b1_16_31_r;
wire signed [`CalcTempBus]          temp_b1_16_31_i;
wire signed [`CalcTempBus]          temp_b1_16_32_r;
wire signed [`CalcTempBus]          temp_b1_16_32_i;
wire signed [`CalcTempBus]          temp_b1_17_1_r;
wire signed [`CalcTempBus]          temp_b1_17_1_i;
wire signed [`CalcTempBus]          temp_b1_17_2_r;
wire signed [`CalcTempBus]          temp_b1_17_2_i;
wire signed [`CalcTempBus]          temp_b1_17_3_r;
wire signed [`CalcTempBus]          temp_b1_17_3_i;
wire signed [`CalcTempBus]          temp_b1_17_4_r;
wire signed [`CalcTempBus]          temp_b1_17_4_i;
wire signed [`CalcTempBus]          temp_b1_17_5_r;
wire signed [`CalcTempBus]          temp_b1_17_5_i;
wire signed [`CalcTempBus]          temp_b1_17_6_r;
wire signed [`CalcTempBus]          temp_b1_17_6_i;
wire signed [`CalcTempBus]          temp_b1_17_7_r;
wire signed [`CalcTempBus]          temp_b1_17_7_i;
wire signed [`CalcTempBus]          temp_b1_17_8_r;
wire signed [`CalcTempBus]          temp_b1_17_8_i;
wire signed [`CalcTempBus]          temp_b1_17_9_r;
wire signed [`CalcTempBus]          temp_b1_17_9_i;
wire signed [`CalcTempBus]          temp_b1_17_10_r;
wire signed [`CalcTempBus]          temp_b1_17_10_i;
wire signed [`CalcTempBus]          temp_b1_17_11_r;
wire signed [`CalcTempBus]          temp_b1_17_11_i;
wire signed [`CalcTempBus]          temp_b1_17_12_r;
wire signed [`CalcTempBus]          temp_b1_17_12_i;
wire signed [`CalcTempBus]          temp_b1_17_13_r;
wire signed [`CalcTempBus]          temp_b1_17_13_i;
wire signed [`CalcTempBus]          temp_b1_17_14_r;
wire signed [`CalcTempBus]          temp_b1_17_14_i;
wire signed [`CalcTempBus]          temp_b1_17_15_r;
wire signed [`CalcTempBus]          temp_b1_17_15_i;
wire signed [`CalcTempBus]          temp_b1_17_16_r;
wire signed [`CalcTempBus]          temp_b1_17_16_i;
wire signed [`CalcTempBus]          temp_b1_17_17_r;
wire signed [`CalcTempBus]          temp_b1_17_17_i;
wire signed [`CalcTempBus]          temp_b1_17_18_r;
wire signed [`CalcTempBus]          temp_b1_17_18_i;
wire signed [`CalcTempBus]          temp_b1_17_19_r;
wire signed [`CalcTempBus]          temp_b1_17_19_i;
wire signed [`CalcTempBus]          temp_b1_17_20_r;
wire signed [`CalcTempBus]          temp_b1_17_20_i;
wire signed [`CalcTempBus]          temp_b1_17_21_r;
wire signed [`CalcTempBus]          temp_b1_17_21_i;
wire signed [`CalcTempBus]          temp_b1_17_22_r;
wire signed [`CalcTempBus]          temp_b1_17_22_i;
wire signed [`CalcTempBus]          temp_b1_17_23_r;
wire signed [`CalcTempBus]          temp_b1_17_23_i;
wire signed [`CalcTempBus]          temp_b1_17_24_r;
wire signed [`CalcTempBus]          temp_b1_17_24_i;
wire signed [`CalcTempBus]          temp_b1_17_25_r;
wire signed [`CalcTempBus]          temp_b1_17_25_i;
wire signed [`CalcTempBus]          temp_b1_17_26_r;
wire signed [`CalcTempBus]          temp_b1_17_26_i;
wire signed [`CalcTempBus]          temp_b1_17_27_r;
wire signed [`CalcTempBus]          temp_b1_17_27_i;
wire signed [`CalcTempBus]          temp_b1_17_28_r;
wire signed [`CalcTempBus]          temp_b1_17_28_i;
wire signed [`CalcTempBus]          temp_b1_17_29_r;
wire signed [`CalcTempBus]          temp_b1_17_29_i;
wire signed [`CalcTempBus]          temp_b1_17_30_r;
wire signed [`CalcTempBus]          temp_b1_17_30_i;
wire signed [`CalcTempBus]          temp_b1_17_31_r;
wire signed [`CalcTempBus]          temp_b1_17_31_i;
wire signed [`CalcTempBus]          temp_b1_17_32_r;
wire signed [`CalcTempBus]          temp_b1_17_32_i;
wire signed [`CalcTempBus]          temp_b1_18_1_r;
wire signed [`CalcTempBus]          temp_b1_18_1_i;
wire signed [`CalcTempBus]          temp_b1_18_2_r;
wire signed [`CalcTempBus]          temp_b1_18_2_i;
wire signed [`CalcTempBus]          temp_b1_18_3_r;
wire signed [`CalcTempBus]          temp_b1_18_3_i;
wire signed [`CalcTempBus]          temp_b1_18_4_r;
wire signed [`CalcTempBus]          temp_b1_18_4_i;
wire signed [`CalcTempBus]          temp_b1_18_5_r;
wire signed [`CalcTempBus]          temp_b1_18_5_i;
wire signed [`CalcTempBus]          temp_b1_18_6_r;
wire signed [`CalcTempBus]          temp_b1_18_6_i;
wire signed [`CalcTempBus]          temp_b1_18_7_r;
wire signed [`CalcTempBus]          temp_b1_18_7_i;
wire signed [`CalcTempBus]          temp_b1_18_8_r;
wire signed [`CalcTempBus]          temp_b1_18_8_i;
wire signed [`CalcTempBus]          temp_b1_18_9_r;
wire signed [`CalcTempBus]          temp_b1_18_9_i;
wire signed [`CalcTempBus]          temp_b1_18_10_r;
wire signed [`CalcTempBus]          temp_b1_18_10_i;
wire signed [`CalcTempBus]          temp_b1_18_11_r;
wire signed [`CalcTempBus]          temp_b1_18_11_i;
wire signed [`CalcTempBus]          temp_b1_18_12_r;
wire signed [`CalcTempBus]          temp_b1_18_12_i;
wire signed [`CalcTempBus]          temp_b1_18_13_r;
wire signed [`CalcTempBus]          temp_b1_18_13_i;
wire signed [`CalcTempBus]          temp_b1_18_14_r;
wire signed [`CalcTempBus]          temp_b1_18_14_i;
wire signed [`CalcTempBus]          temp_b1_18_15_r;
wire signed [`CalcTempBus]          temp_b1_18_15_i;
wire signed [`CalcTempBus]          temp_b1_18_16_r;
wire signed [`CalcTempBus]          temp_b1_18_16_i;
wire signed [`CalcTempBus]          temp_b1_18_17_r;
wire signed [`CalcTempBus]          temp_b1_18_17_i;
wire signed [`CalcTempBus]          temp_b1_18_18_r;
wire signed [`CalcTempBus]          temp_b1_18_18_i;
wire signed [`CalcTempBus]          temp_b1_18_19_r;
wire signed [`CalcTempBus]          temp_b1_18_19_i;
wire signed [`CalcTempBus]          temp_b1_18_20_r;
wire signed [`CalcTempBus]          temp_b1_18_20_i;
wire signed [`CalcTempBus]          temp_b1_18_21_r;
wire signed [`CalcTempBus]          temp_b1_18_21_i;
wire signed [`CalcTempBus]          temp_b1_18_22_r;
wire signed [`CalcTempBus]          temp_b1_18_22_i;
wire signed [`CalcTempBus]          temp_b1_18_23_r;
wire signed [`CalcTempBus]          temp_b1_18_23_i;
wire signed [`CalcTempBus]          temp_b1_18_24_r;
wire signed [`CalcTempBus]          temp_b1_18_24_i;
wire signed [`CalcTempBus]          temp_b1_18_25_r;
wire signed [`CalcTempBus]          temp_b1_18_25_i;
wire signed [`CalcTempBus]          temp_b1_18_26_r;
wire signed [`CalcTempBus]          temp_b1_18_26_i;
wire signed [`CalcTempBus]          temp_b1_18_27_r;
wire signed [`CalcTempBus]          temp_b1_18_27_i;
wire signed [`CalcTempBus]          temp_b1_18_28_r;
wire signed [`CalcTempBus]          temp_b1_18_28_i;
wire signed [`CalcTempBus]          temp_b1_18_29_r;
wire signed [`CalcTempBus]          temp_b1_18_29_i;
wire signed [`CalcTempBus]          temp_b1_18_30_r;
wire signed [`CalcTempBus]          temp_b1_18_30_i;
wire signed [`CalcTempBus]          temp_b1_18_31_r;
wire signed [`CalcTempBus]          temp_b1_18_31_i;
wire signed [`CalcTempBus]          temp_b1_18_32_r;
wire signed [`CalcTempBus]          temp_b1_18_32_i;
wire signed [`CalcTempBus]          temp_b1_19_1_r;
wire signed [`CalcTempBus]          temp_b1_19_1_i;
wire signed [`CalcTempBus]          temp_b1_19_2_r;
wire signed [`CalcTempBus]          temp_b1_19_2_i;
wire signed [`CalcTempBus]          temp_b1_19_3_r;
wire signed [`CalcTempBus]          temp_b1_19_3_i;
wire signed [`CalcTempBus]          temp_b1_19_4_r;
wire signed [`CalcTempBus]          temp_b1_19_4_i;
wire signed [`CalcTempBus]          temp_b1_19_5_r;
wire signed [`CalcTempBus]          temp_b1_19_5_i;
wire signed [`CalcTempBus]          temp_b1_19_6_r;
wire signed [`CalcTempBus]          temp_b1_19_6_i;
wire signed [`CalcTempBus]          temp_b1_19_7_r;
wire signed [`CalcTempBus]          temp_b1_19_7_i;
wire signed [`CalcTempBus]          temp_b1_19_8_r;
wire signed [`CalcTempBus]          temp_b1_19_8_i;
wire signed [`CalcTempBus]          temp_b1_19_9_r;
wire signed [`CalcTempBus]          temp_b1_19_9_i;
wire signed [`CalcTempBus]          temp_b1_19_10_r;
wire signed [`CalcTempBus]          temp_b1_19_10_i;
wire signed [`CalcTempBus]          temp_b1_19_11_r;
wire signed [`CalcTempBus]          temp_b1_19_11_i;
wire signed [`CalcTempBus]          temp_b1_19_12_r;
wire signed [`CalcTempBus]          temp_b1_19_12_i;
wire signed [`CalcTempBus]          temp_b1_19_13_r;
wire signed [`CalcTempBus]          temp_b1_19_13_i;
wire signed [`CalcTempBus]          temp_b1_19_14_r;
wire signed [`CalcTempBus]          temp_b1_19_14_i;
wire signed [`CalcTempBus]          temp_b1_19_15_r;
wire signed [`CalcTempBus]          temp_b1_19_15_i;
wire signed [`CalcTempBus]          temp_b1_19_16_r;
wire signed [`CalcTempBus]          temp_b1_19_16_i;
wire signed [`CalcTempBus]          temp_b1_19_17_r;
wire signed [`CalcTempBus]          temp_b1_19_17_i;
wire signed [`CalcTempBus]          temp_b1_19_18_r;
wire signed [`CalcTempBus]          temp_b1_19_18_i;
wire signed [`CalcTempBus]          temp_b1_19_19_r;
wire signed [`CalcTempBus]          temp_b1_19_19_i;
wire signed [`CalcTempBus]          temp_b1_19_20_r;
wire signed [`CalcTempBus]          temp_b1_19_20_i;
wire signed [`CalcTempBus]          temp_b1_19_21_r;
wire signed [`CalcTempBus]          temp_b1_19_21_i;
wire signed [`CalcTempBus]          temp_b1_19_22_r;
wire signed [`CalcTempBus]          temp_b1_19_22_i;
wire signed [`CalcTempBus]          temp_b1_19_23_r;
wire signed [`CalcTempBus]          temp_b1_19_23_i;
wire signed [`CalcTempBus]          temp_b1_19_24_r;
wire signed [`CalcTempBus]          temp_b1_19_24_i;
wire signed [`CalcTempBus]          temp_b1_19_25_r;
wire signed [`CalcTempBus]          temp_b1_19_25_i;
wire signed [`CalcTempBus]          temp_b1_19_26_r;
wire signed [`CalcTempBus]          temp_b1_19_26_i;
wire signed [`CalcTempBus]          temp_b1_19_27_r;
wire signed [`CalcTempBus]          temp_b1_19_27_i;
wire signed [`CalcTempBus]          temp_b1_19_28_r;
wire signed [`CalcTempBus]          temp_b1_19_28_i;
wire signed [`CalcTempBus]          temp_b1_19_29_r;
wire signed [`CalcTempBus]          temp_b1_19_29_i;
wire signed [`CalcTempBus]          temp_b1_19_30_r;
wire signed [`CalcTempBus]          temp_b1_19_30_i;
wire signed [`CalcTempBus]          temp_b1_19_31_r;
wire signed [`CalcTempBus]          temp_b1_19_31_i;
wire signed [`CalcTempBus]          temp_b1_19_32_r;
wire signed [`CalcTempBus]          temp_b1_19_32_i;
wire signed [`CalcTempBus]          temp_b1_20_1_r;
wire signed [`CalcTempBus]          temp_b1_20_1_i;
wire signed [`CalcTempBus]          temp_b1_20_2_r;
wire signed [`CalcTempBus]          temp_b1_20_2_i;
wire signed [`CalcTempBus]          temp_b1_20_3_r;
wire signed [`CalcTempBus]          temp_b1_20_3_i;
wire signed [`CalcTempBus]          temp_b1_20_4_r;
wire signed [`CalcTempBus]          temp_b1_20_4_i;
wire signed [`CalcTempBus]          temp_b1_20_5_r;
wire signed [`CalcTempBus]          temp_b1_20_5_i;
wire signed [`CalcTempBus]          temp_b1_20_6_r;
wire signed [`CalcTempBus]          temp_b1_20_6_i;
wire signed [`CalcTempBus]          temp_b1_20_7_r;
wire signed [`CalcTempBus]          temp_b1_20_7_i;
wire signed [`CalcTempBus]          temp_b1_20_8_r;
wire signed [`CalcTempBus]          temp_b1_20_8_i;
wire signed [`CalcTempBus]          temp_b1_20_9_r;
wire signed [`CalcTempBus]          temp_b1_20_9_i;
wire signed [`CalcTempBus]          temp_b1_20_10_r;
wire signed [`CalcTempBus]          temp_b1_20_10_i;
wire signed [`CalcTempBus]          temp_b1_20_11_r;
wire signed [`CalcTempBus]          temp_b1_20_11_i;
wire signed [`CalcTempBus]          temp_b1_20_12_r;
wire signed [`CalcTempBus]          temp_b1_20_12_i;
wire signed [`CalcTempBus]          temp_b1_20_13_r;
wire signed [`CalcTempBus]          temp_b1_20_13_i;
wire signed [`CalcTempBus]          temp_b1_20_14_r;
wire signed [`CalcTempBus]          temp_b1_20_14_i;
wire signed [`CalcTempBus]          temp_b1_20_15_r;
wire signed [`CalcTempBus]          temp_b1_20_15_i;
wire signed [`CalcTempBus]          temp_b1_20_16_r;
wire signed [`CalcTempBus]          temp_b1_20_16_i;
wire signed [`CalcTempBus]          temp_b1_20_17_r;
wire signed [`CalcTempBus]          temp_b1_20_17_i;
wire signed [`CalcTempBus]          temp_b1_20_18_r;
wire signed [`CalcTempBus]          temp_b1_20_18_i;
wire signed [`CalcTempBus]          temp_b1_20_19_r;
wire signed [`CalcTempBus]          temp_b1_20_19_i;
wire signed [`CalcTempBus]          temp_b1_20_20_r;
wire signed [`CalcTempBus]          temp_b1_20_20_i;
wire signed [`CalcTempBus]          temp_b1_20_21_r;
wire signed [`CalcTempBus]          temp_b1_20_21_i;
wire signed [`CalcTempBus]          temp_b1_20_22_r;
wire signed [`CalcTempBus]          temp_b1_20_22_i;
wire signed [`CalcTempBus]          temp_b1_20_23_r;
wire signed [`CalcTempBus]          temp_b1_20_23_i;
wire signed [`CalcTempBus]          temp_b1_20_24_r;
wire signed [`CalcTempBus]          temp_b1_20_24_i;
wire signed [`CalcTempBus]          temp_b1_20_25_r;
wire signed [`CalcTempBus]          temp_b1_20_25_i;
wire signed [`CalcTempBus]          temp_b1_20_26_r;
wire signed [`CalcTempBus]          temp_b1_20_26_i;
wire signed [`CalcTempBus]          temp_b1_20_27_r;
wire signed [`CalcTempBus]          temp_b1_20_27_i;
wire signed [`CalcTempBus]          temp_b1_20_28_r;
wire signed [`CalcTempBus]          temp_b1_20_28_i;
wire signed [`CalcTempBus]          temp_b1_20_29_r;
wire signed [`CalcTempBus]          temp_b1_20_29_i;
wire signed [`CalcTempBus]          temp_b1_20_30_r;
wire signed [`CalcTempBus]          temp_b1_20_30_i;
wire signed [`CalcTempBus]          temp_b1_20_31_r;
wire signed [`CalcTempBus]          temp_b1_20_31_i;
wire signed [`CalcTempBus]          temp_b1_20_32_r;
wire signed [`CalcTempBus]          temp_b1_20_32_i;
wire signed [`CalcTempBus]          temp_b1_21_1_r;
wire signed [`CalcTempBus]          temp_b1_21_1_i;
wire signed [`CalcTempBus]          temp_b1_21_2_r;
wire signed [`CalcTempBus]          temp_b1_21_2_i;
wire signed [`CalcTempBus]          temp_b1_21_3_r;
wire signed [`CalcTempBus]          temp_b1_21_3_i;
wire signed [`CalcTempBus]          temp_b1_21_4_r;
wire signed [`CalcTempBus]          temp_b1_21_4_i;
wire signed [`CalcTempBus]          temp_b1_21_5_r;
wire signed [`CalcTempBus]          temp_b1_21_5_i;
wire signed [`CalcTempBus]          temp_b1_21_6_r;
wire signed [`CalcTempBus]          temp_b1_21_6_i;
wire signed [`CalcTempBus]          temp_b1_21_7_r;
wire signed [`CalcTempBus]          temp_b1_21_7_i;
wire signed [`CalcTempBus]          temp_b1_21_8_r;
wire signed [`CalcTempBus]          temp_b1_21_8_i;
wire signed [`CalcTempBus]          temp_b1_21_9_r;
wire signed [`CalcTempBus]          temp_b1_21_9_i;
wire signed [`CalcTempBus]          temp_b1_21_10_r;
wire signed [`CalcTempBus]          temp_b1_21_10_i;
wire signed [`CalcTempBus]          temp_b1_21_11_r;
wire signed [`CalcTempBus]          temp_b1_21_11_i;
wire signed [`CalcTempBus]          temp_b1_21_12_r;
wire signed [`CalcTempBus]          temp_b1_21_12_i;
wire signed [`CalcTempBus]          temp_b1_21_13_r;
wire signed [`CalcTempBus]          temp_b1_21_13_i;
wire signed [`CalcTempBus]          temp_b1_21_14_r;
wire signed [`CalcTempBus]          temp_b1_21_14_i;
wire signed [`CalcTempBus]          temp_b1_21_15_r;
wire signed [`CalcTempBus]          temp_b1_21_15_i;
wire signed [`CalcTempBus]          temp_b1_21_16_r;
wire signed [`CalcTempBus]          temp_b1_21_16_i;
wire signed [`CalcTempBus]          temp_b1_21_17_r;
wire signed [`CalcTempBus]          temp_b1_21_17_i;
wire signed [`CalcTempBus]          temp_b1_21_18_r;
wire signed [`CalcTempBus]          temp_b1_21_18_i;
wire signed [`CalcTempBus]          temp_b1_21_19_r;
wire signed [`CalcTempBus]          temp_b1_21_19_i;
wire signed [`CalcTempBus]          temp_b1_21_20_r;
wire signed [`CalcTempBus]          temp_b1_21_20_i;
wire signed [`CalcTempBus]          temp_b1_21_21_r;
wire signed [`CalcTempBus]          temp_b1_21_21_i;
wire signed [`CalcTempBus]          temp_b1_21_22_r;
wire signed [`CalcTempBus]          temp_b1_21_22_i;
wire signed [`CalcTempBus]          temp_b1_21_23_r;
wire signed [`CalcTempBus]          temp_b1_21_23_i;
wire signed [`CalcTempBus]          temp_b1_21_24_r;
wire signed [`CalcTempBus]          temp_b1_21_24_i;
wire signed [`CalcTempBus]          temp_b1_21_25_r;
wire signed [`CalcTempBus]          temp_b1_21_25_i;
wire signed [`CalcTempBus]          temp_b1_21_26_r;
wire signed [`CalcTempBus]          temp_b1_21_26_i;
wire signed [`CalcTempBus]          temp_b1_21_27_r;
wire signed [`CalcTempBus]          temp_b1_21_27_i;
wire signed [`CalcTempBus]          temp_b1_21_28_r;
wire signed [`CalcTempBus]          temp_b1_21_28_i;
wire signed [`CalcTempBus]          temp_b1_21_29_r;
wire signed [`CalcTempBus]          temp_b1_21_29_i;
wire signed [`CalcTempBus]          temp_b1_21_30_r;
wire signed [`CalcTempBus]          temp_b1_21_30_i;
wire signed [`CalcTempBus]          temp_b1_21_31_r;
wire signed [`CalcTempBus]          temp_b1_21_31_i;
wire signed [`CalcTempBus]          temp_b1_21_32_r;
wire signed [`CalcTempBus]          temp_b1_21_32_i;
wire signed [`CalcTempBus]          temp_b1_22_1_r;
wire signed [`CalcTempBus]          temp_b1_22_1_i;
wire signed [`CalcTempBus]          temp_b1_22_2_r;
wire signed [`CalcTempBus]          temp_b1_22_2_i;
wire signed [`CalcTempBus]          temp_b1_22_3_r;
wire signed [`CalcTempBus]          temp_b1_22_3_i;
wire signed [`CalcTempBus]          temp_b1_22_4_r;
wire signed [`CalcTempBus]          temp_b1_22_4_i;
wire signed [`CalcTempBus]          temp_b1_22_5_r;
wire signed [`CalcTempBus]          temp_b1_22_5_i;
wire signed [`CalcTempBus]          temp_b1_22_6_r;
wire signed [`CalcTempBus]          temp_b1_22_6_i;
wire signed [`CalcTempBus]          temp_b1_22_7_r;
wire signed [`CalcTempBus]          temp_b1_22_7_i;
wire signed [`CalcTempBus]          temp_b1_22_8_r;
wire signed [`CalcTempBus]          temp_b1_22_8_i;
wire signed [`CalcTempBus]          temp_b1_22_9_r;
wire signed [`CalcTempBus]          temp_b1_22_9_i;
wire signed [`CalcTempBus]          temp_b1_22_10_r;
wire signed [`CalcTempBus]          temp_b1_22_10_i;
wire signed [`CalcTempBus]          temp_b1_22_11_r;
wire signed [`CalcTempBus]          temp_b1_22_11_i;
wire signed [`CalcTempBus]          temp_b1_22_12_r;
wire signed [`CalcTempBus]          temp_b1_22_12_i;
wire signed [`CalcTempBus]          temp_b1_22_13_r;
wire signed [`CalcTempBus]          temp_b1_22_13_i;
wire signed [`CalcTempBus]          temp_b1_22_14_r;
wire signed [`CalcTempBus]          temp_b1_22_14_i;
wire signed [`CalcTempBus]          temp_b1_22_15_r;
wire signed [`CalcTempBus]          temp_b1_22_15_i;
wire signed [`CalcTempBus]          temp_b1_22_16_r;
wire signed [`CalcTempBus]          temp_b1_22_16_i;
wire signed [`CalcTempBus]          temp_b1_22_17_r;
wire signed [`CalcTempBus]          temp_b1_22_17_i;
wire signed [`CalcTempBus]          temp_b1_22_18_r;
wire signed [`CalcTempBus]          temp_b1_22_18_i;
wire signed [`CalcTempBus]          temp_b1_22_19_r;
wire signed [`CalcTempBus]          temp_b1_22_19_i;
wire signed [`CalcTempBus]          temp_b1_22_20_r;
wire signed [`CalcTempBus]          temp_b1_22_20_i;
wire signed [`CalcTempBus]          temp_b1_22_21_r;
wire signed [`CalcTempBus]          temp_b1_22_21_i;
wire signed [`CalcTempBus]          temp_b1_22_22_r;
wire signed [`CalcTempBus]          temp_b1_22_22_i;
wire signed [`CalcTempBus]          temp_b1_22_23_r;
wire signed [`CalcTempBus]          temp_b1_22_23_i;
wire signed [`CalcTempBus]          temp_b1_22_24_r;
wire signed [`CalcTempBus]          temp_b1_22_24_i;
wire signed [`CalcTempBus]          temp_b1_22_25_r;
wire signed [`CalcTempBus]          temp_b1_22_25_i;
wire signed [`CalcTempBus]          temp_b1_22_26_r;
wire signed [`CalcTempBus]          temp_b1_22_26_i;
wire signed [`CalcTempBus]          temp_b1_22_27_r;
wire signed [`CalcTempBus]          temp_b1_22_27_i;
wire signed [`CalcTempBus]          temp_b1_22_28_r;
wire signed [`CalcTempBus]          temp_b1_22_28_i;
wire signed [`CalcTempBus]          temp_b1_22_29_r;
wire signed [`CalcTempBus]          temp_b1_22_29_i;
wire signed [`CalcTempBus]          temp_b1_22_30_r;
wire signed [`CalcTempBus]          temp_b1_22_30_i;
wire signed [`CalcTempBus]          temp_b1_22_31_r;
wire signed [`CalcTempBus]          temp_b1_22_31_i;
wire signed [`CalcTempBus]          temp_b1_22_32_r;
wire signed [`CalcTempBus]          temp_b1_22_32_i;
wire signed [`CalcTempBus]          temp_b1_23_1_r;
wire signed [`CalcTempBus]          temp_b1_23_1_i;
wire signed [`CalcTempBus]          temp_b1_23_2_r;
wire signed [`CalcTempBus]          temp_b1_23_2_i;
wire signed [`CalcTempBus]          temp_b1_23_3_r;
wire signed [`CalcTempBus]          temp_b1_23_3_i;
wire signed [`CalcTempBus]          temp_b1_23_4_r;
wire signed [`CalcTempBus]          temp_b1_23_4_i;
wire signed [`CalcTempBus]          temp_b1_23_5_r;
wire signed [`CalcTempBus]          temp_b1_23_5_i;
wire signed [`CalcTempBus]          temp_b1_23_6_r;
wire signed [`CalcTempBus]          temp_b1_23_6_i;
wire signed [`CalcTempBus]          temp_b1_23_7_r;
wire signed [`CalcTempBus]          temp_b1_23_7_i;
wire signed [`CalcTempBus]          temp_b1_23_8_r;
wire signed [`CalcTempBus]          temp_b1_23_8_i;
wire signed [`CalcTempBus]          temp_b1_23_9_r;
wire signed [`CalcTempBus]          temp_b1_23_9_i;
wire signed [`CalcTempBus]          temp_b1_23_10_r;
wire signed [`CalcTempBus]          temp_b1_23_10_i;
wire signed [`CalcTempBus]          temp_b1_23_11_r;
wire signed [`CalcTempBus]          temp_b1_23_11_i;
wire signed [`CalcTempBus]          temp_b1_23_12_r;
wire signed [`CalcTempBus]          temp_b1_23_12_i;
wire signed [`CalcTempBus]          temp_b1_23_13_r;
wire signed [`CalcTempBus]          temp_b1_23_13_i;
wire signed [`CalcTempBus]          temp_b1_23_14_r;
wire signed [`CalcTempBus]          temp_b1_23_14_i;
wire signed [`CalcTempBus]          temp_b1_23_15_r;
wire signed [`CalcTempBus]          temp_b1_23_15_i;
wire signed [`CalcTempBus]          temp_b1_23_16_r;
wire signed [`CalcTempBus]          temp_b1_23_16_i;
wire signed [`CalcTempBus]          temp_b1_23_17_r;
wire signed [`CalcTempBus]          temp_b1_23_17_i;
wire signed [`CalcTempBus]          temp_b1_23_18_r;
wire signed [`CalcTempBus]          temp_b1_23_18_i;
wire signed [`CalcTempBus]          temp_b1_23_19_r;
wire signed [`CalcTempBus]          temp_b1_23_19_i;
wire signed [`CalcTempBus]          temp_b1_23_20_r;
wire signed [`CalcTempBus]          temp_b1_23_20_i;
wire signed [`CalcTempBus]          temp_b1_23_21_r;
wire signed [`CalcTempBus]          temp_b1_23_21_i;
wire signed [`CalcTempBus]          temp_b1_23_22_r;
wire signed [`CalcTempBus]          temp_b1_23_22_i;
wire signed [`CalcTempBus]          temp_b1_23_23_r;
wire signed [`CalcTempBus]          temp_b1_23_23_i;
wire signed [`CalcTempBus]          temp_b1_23_24_r;
wire signed [`CalcTempBus]          temp_b1_23_24_i;
wire signed [`CalcTempBus]          temp_b1_23_25_r;
wire signed [`CalcTempBus]          temp_b1_23_25_i;
wire signed [`CalcTempBus]          temp_b1_23_26_r;
wire signed [`CalcTempBus]          temp_b1_23_26_i;
wire signed [`CalcTempBus]          temp_b1_23_27_r;
wire signed [`CalcTempBus]          temp_b1_23_27_i;
wire signed [`CalcTempBus]          temp_b1_23_28_r;
wire signed [`CalcTempBus]          temp_b1_23_28_i;
wire signed [`CalcTempBus]          temp_b1_23_29_r;
wire signed [`CalcTempBus]          temp_b1_23_29_i;
wire signed [`CalcTempBus]          temp_b1_23_30_r;
wire signed [`CalcTempBus]          temp_b1_23_30_i;
wire signed [`CalcTempBus]          temp_b1_23_31_r;
wire signed [`CalcTempBus]          temp_b1_23_31_i;
wire signed [`CalcTempBus]          temp_b1_23_32_r;
wire signed [`CalcTempBus]          temp_b1_23_32_i;
wire signed [`CalcTempBus]          temp_b1_24_1_r;
wire signed [`CalcTempBus]          temp_b1_24_1_i;
wire signed [`CalcTempBus]          temp_b1_24_2_r;
wire signed [`CalcTempBus]          temp_b1_24_2_i;
wire signed [`CalcTempBus]          temp_b1_24_3_r;
wire signed [`CalcTempBus]          temp_b1_24_3_i;
wire signed [`CalcTempBus]          temp_b1_24_4_r;
wire signed [`CalcTempBus]          temp_b1_24_4_i;
wire signed [`CalcTempBus]          temp_b1_24_5_r;
wire signed [`CalcTempBus]          temp_b1_24_5_i;
wire signed [`CalcTempBus]          temp_b1_24_6_r;
wire signed [`CalcTempBus]          temp_b1_24_6_i;
wire signed [`CalcTempBus]          temp_b1_24_7_r;
wire signed [`CalcTempBus]          temp_b1_24_7_i;
wire signed [`CalcTempBus]          temp_b1_24_8_r;
wire signed [`CalcTempBus]          temp_b1_24_8_i;
wire signed [`CalcTempBus]          temp_b1_24_9_r;
wire signed [`CalcTempBus]          temp_b1_24_9_i;
wire signed [`CalcTempBus]          temp_b1_24_10_r;
wire signed [`CalcTempBus]          temp_b1_24_10_i;
wire signed [`CalcTempBus]          temp_b1_24_11_r;
wire signed [`CalcTempBus]          temp_b1_24_11_i;
wire signed [`CalcTempBus]          temp_b1_24_12_r;
wire signed [`CalcTempBus]          temp_b1_24_12_i;
wire signed [`CalcTempBus]          temp_b1_24_13_r;
wire signed [`CalcTempBus]          temp_b1_24_13_i;
wire signed [`CalcTempBus]          temp_b1_24_14_r;
wire signed [`CalcTempBus]          temp_b1_24_14_i;
wire signed [`CalcTempBus]          temp_b1_24_15_r;
wire signed [`CalcTempBus]          temp_b1_24_15_i;
wire signed [`CalcTempBus]          temp_b1_24_16_r;
wire signed [`CalcTempBus]          temp_b1_24_16_i;
wire signed [`CalcTempBus]          temp_b1_24_17_r;
wire signed [`CalcTempBus]          temp_b1_24_17_i;
wire signed [`CalcTempBus]          temp_b1_24_18_r;
wire signed [`CalcTempBus]          temp_b1_24_18_i;
wire signed [`CalcTempBus]          temp_b1_24_19_r;
wire signed [`CalcTempBus]          temp_b1_24_19_i;
wire signed [`CalcTempBus]          temp_b1_24_20_r;
wire signed [`CalcTempBus]          temp_b1_24_20_i;
wire signed [`CalcTempBus]          temp_b1_24_21_r;
wire signed [`CalcTempBus]          temp_b1_24_21_i;
wire signed [`CalcTempBus]          temp_b1_24_22_r;
wire signed [`CalcTempBus]          temp_b1_24_22_i;
wire signed [`CalcTempBus]          temp_b1_24_23_r;
wire signed [`CalcTempBus]          temp_b1_24_23_i;
wire signed [`CalcTempBus]          temp_b1_24_24_r;
wire signed [`CalcTempBus]          temp_b1_24_24_i;
wire signed [`CalcTempBus]          temp_b1_24_25_r;
wire signed [`CalcTempBus]          temp_b1_24_25_i;
wire signed [`CalcTempBus]          temp_b1_24_26_r;
wire signed [`CalcTempBus]          temp_b1_24_26_i;
wire signed [`CalcTempBus]          temp_b1_24_27_r;
wire signed [`CalcTempBus]          temp_b1_24_27_i;
wire signed [`CalcTempBus]          temp_b1_24_28_r;
wire signed [`CalcTempBus]          temp_b1_24_28_i;
wire signed [`CalcTempBus]          temp_b1_24_29_r;
wire signed [`CalcTempBus]          temp_b1_24_29_i;
wire signed [`CalcTempBus]          temp_b1_24_30_r;
wire signed [`CalcTempBus]          temp_b1_24_30_i;
wire signed [`CalcTempBus]          temp_b1_24_31_r;
wire signed [`CalcTempBus]          temp_b1_24_31_i;
wire signed [`CalcTempBus]          temp_b1_24_32_r;
wire signed [`CalcTempBus]          temp_b1_24_32_i;
wire signed [`CalcTempBus]          temp_b1_25_1_r;
wire signed [`CalcTempBus]          temp_b1_25_1_i;
wire signed [`CalcTempBus]          temp_b1_25_2_r;
wire signed [`CalcTempBus]          temp_b1_25_2_i;
wire signed [`CalcTempBus]          temp_b1_25_3_r;
wire signed [`CalcTempBus]          temp_b1_25_3_i;
wire signed [`CalcTempBus]          temp_b1_25_4_r;
wire signed [`CalcTempBus]          temp_b1_25_4_i;
wire signed [`CalcTempBus]          temp_b1_25_5_r;
wire signed [`CalcTempBus]          temp_b1_25_5_i;
wire signed [`CalcTempBus]          temp_b1_25_6_r;
wire signed [`CalcTempBus]          temp_b1_25_6_i;
wire signed [`CalcTempBus]          temp_b1_25_7_r;
wire signed [`CalcTempBus]          temp_b1_25_7_i;
wire signed [`CalcTempBus]          temp_b1_25_8_r;
wire signed [`CalcTempBus]          temp_b1_25_8_i;
wire signed [`CalcTempBus]          temp_b1_25_9_r;
wire signed [`CalcTempBus]          temp_b1_25_9_i;
wire signed [`CalcTempBus]          temp_b1_25_10_r;
wire signed [`CalcTempBus]          temp_b1_25_10_i;
wire signed [`CalcTempBus]          temp_b1_25_11_r;
wire signed [`CalcTempBus]          temp_b1_25_11_i;
wire signed [`CalcTempBus]          temp_b1_25_12_r;
wire signed [`CalcTempBus]          temp_b1_25_12_i;
wire signed [`CalcTempBus]          temp_b1_25_13_r;
wire signed [`CalcTempBus]          temp_b1_25_13_i;
wire signed [`CalcTempBus]          temp_b1_25_14_r;
wire signed [`CalcTempBus]          temp_b1_25_14_i;
wire signed [`CalcTempBus]          temp_b1_25_15_r;
wire signed [`CalcTempBus]          temp_b1_25_15_i;
wire signed [`CalcTempBus]          temp_b1_25_16_r;
wire signed [`CalcTempBus]          temp_b1_25_16_i;
wire signed [`CalcTempBus]          temp_b1_25_17_r;
wire signed [`CalcTempBus]          temp_b1_25_17_i;
wire signed [`CalcTempBus]          temp_b1_25_18_r;
wire signed [`CalcTempBus]          temp_b1_25_18_i;
wire signed [`CalcTempBus]          temp_b1_25_19_r;
wire signed [`CalcTempBus]          temp_b1_25_19_i;
wire signed [`CalcTempBus]          temp_b1_25_20_r;
wire signed [`CalcTempBus]          temp_b1_25_20_i;
wire signed [`CalcTempBus]          temp_b1_25_21_r;
wire signed [`CalcTempBus]          temp_b1_25_21_i;
wire signed [`CalcTempBus]          temp_b1_25_22_r;
wire signed [`CalcTempBus]          temp_b1_25_22_i;
wire signed [`CalcTempBus]          temp_b1_25_23_r;
wire signed [`CalcTempBus]          temp_b1_25_23_i;
wire signed [`CalcTempBus]          temp_b1_25_24_r;
wire signed [`CalcTempBus]          temp_b1_25_24_i;
wire signed [`CalcTempBus]          temp_b1_25_25_r;
wire signed [`CalcTempBus]          temp_b1_25_25_i;
wire signed [`CalcTempBus]          temp_b1_25_26_r;
wire signed [`CalcTempBus]          temp_b1_25_26_i;
wire signed [`CalcTempBus]          temp_b1_25_27_r;
wire signed [`CalcTempBus]          temp_b1_25_27_i;
wire signed [`CalcTempBus]          temp_b1_25_28_r;
wire signed [`CalcTempBus]          temp_b1_25_28_i;
wire signed [`CalcTempBus]          temp_b1_25_29_r;
wire signed [`CalcTempBus]          temp_b1_25_29_i;
wire signed [`CalcTempBus]          temp_b1_25_30_r;
wire signed [`CalcTempBus]          temp_b1_25_30_i;
wire signed [`CalcTempBus]          temp_b1_25_31_r;
wire signed [`CalcTempBus]          temp_b1_25_31_i;
wire signed [`CalcTempBus]          temp_b1_25_32_r;
wire signed [`CalcTempBus]          temp_b1_25_32_i;
wire signed [`CalcTempBus]          temp_b1_26_1_r;
wire signed [`CalcTempBus]          temp_b1_26_1_i;
wire signed [`CalcTempBus]          temp_b1_26_2_r;
wire signed [`CalcTempBus]          temp_b1_26_2_i;
wire signed [`CalcTempBus]          temp_b1_26_3_r;
wire signed [`CalcTempBus]          temp_b1_26_3_i;
wire signed [`CalcTempBus]          temp_b1_26_4_r;
wire signed [`CalcTempBus]          temp_b1_26_4_i;
wire signed [`CalcTempBus]          temp_b1_26_5_r;
wire signed [`CalcTempBus]          temp_b1_26_5_i;
wire signed [`CalcTempBus]          temp_b1_26_6_r;
wire signed [`CalcTempBus]          temp_b1_26_6_i;
wire signed [`CalcTempBus]          temp_b1_26_7_r;
wire signed [`CalcTempBus]          temp_b1_26_7_i;
wire signed [`CalcTempBus]          temp_b1_26_8_r;
wire signed [`CalcTempBus]          temp_b1_26_8_i;
wire signed [`CalcTempBus]          temp_b1_26_9_r;
wire signed [`CalcTempBus]          temp_b1_26_9_i;
wire signed [`CalcTempBus]          temp_b1_26_10_r;
wire signed [`CalcTempBus]          temp_b1_26_10_i;
wire signed [`CalcTempBus]          temp_b1_26_11_r;
wire signed [`CalcTempBus]          temp_b1_26_11_i;
wire signed [`CalcTempBus]          temp_b1_26_12_r;
wire signed [`CalcTempBus]          temp_b1_26_12_i;
wire signed [`CalcTempBus]          temp_b1_26_13_r;
wire signed [`CalcTempBus]          temp_b1_26_13_i;
wire signed [`CalcTempBus]          temp_b1_26_14_r;
wire signed [`CalcTempBus]          temp_b1_26_14_i;
wire signed [`CalcTempBus]          temp_b1_26_15_r;
wire signed [`CalcTempBus]          temp_b1_26_15_i;
wire signed [`CalcTempBus]          temp_b1_26_16_r;
wire signed [`CalcTempBus]          temp_b1_26_16_i;
wire signed [`CalcTempBus]          temp_b1_26_17_r;
wire signed [`CalcTempBus]          temp_b1_26_17_i;
wire signed [`CalcTempBus]          temp_b1_26_18_r;
wire signed [`CalcTempBus]          temp_b1_26_18_i;
wire signed [`CalcTempBus]          temp_b1_26_19_r;
wire signed [`CalcTempBus]          temp_b1_26_19_i;
wire signed [`CalcTempBus]          temp_b1_26_20_r;
wire signed [`CalcTempBus]          temp_b1_26_20_i;
wire signed [`CalcTempBus]          temp_b1_26_21_r;
wire signed [`CalcTempBus]          temp_b1_26_21_i;
wire signed [`CalcTempBus]          temp_b1_26_22_r;
wire signed [`CalcTempBus]          temp_b1_26_22_i;
wire signed [`CalcTempBus]          temp_b1_26_23_r;
wire signed [`CalcTempBus]          temp_b1_26_23_i;
wire signed [`CalcTempBus]          temp_b1_26_24_r;
wire signed [`CalcTempBus]          temp_b1_26_24_i;
wire signed [`CalcTempBus]          temp_b1_26_25_r;
wire signed [`CalcTempBus]          temp_b1_26_25_i;
wire signed [`CalcTempBus]          temp_b1_26_26_r;
wire signed [`CalcTempBus]          temp_b1_26_26_i;
wire signed [`CalcTempBus]          temp_b1_26_27_r;
wire signed [`CalcTempBus]          temp_b1_26_27_i;
wire signed [`CalcTempBus]          temp_b1_26_28_r;
wire signed [`CalcTempBus]          temp_b1_26_28_i;
wire signed [`CalcTempBus]          temp_b1_26_29_r;
wire signed [`CalcTempBus]          temp_b1_26_29_i;
wire signed [`CalcTempBus]          temp_b1_26_30_r;
wire signed [`CalcTempBus]          temp_b1_26_30_i;
wire signed [`CalcTempBus]          temp_b1_26_31_r;
wire signed [`CalcTempBus]          temp_b1_26_31_i;
wire signed [`CalcTempBus]          temp_b1_26_32_r;
wire signed [`CalcTempBus]          temp_b1_26_32_i;
wire signed [`CalcTempBus]          temp_b1_27_1_r;
wire signed [`CalcTempBus]          temp_b1_27_1_i;
wire signed [`CalcTempBus]          temp_b1_27_2_r;
wire signed [`CalcTempBus]          temp_b1_27_2_i;
wire signed [`CalcTempBus]          temp_b1_27_3_r;
wire signed [`CalcTempBus]          temp_b1_27_3_i;
wire signed [`CalcTempBus]          temp_b1_27_4_r;
wire signed [`CalcTempBus]          temp_b1_27_4_i;
wire signed [`CalcTempBus]          temp_b1_27_5_r;
wire signed [`CalcTempBus]          temp_b1_27_5_i;
wire signed [`CalcTempBus]          temp_b1_27_6_r;
wire signed [`CalcTempBus]          temp_b1_27_6_i;
wire signed [`CalcTempBus]          temp_b1_27_7_r;
wire signed [`CalcTempBus]          temp_b1_27_7_i;
wire signed [`CalcTempBus]          temp_b1_27_8_r;
wire signed [`CalcTempBus]          temp_b1_27_8_i;
wire signed [`CalcTempBus]          temp_b1_27_9_r;
wire signed [`CalcTempBus]          temp_b1_27_9_i;
wire signed [`CalcTempBus]          temp_b1_27_10_r;
wire signed [`CalcTempBus]          temp_b1_27_10_i;
wire signed [`CalcTempBus]          temp_b1_27_11_r;
wire signed [`CalcTempBus]          temp_b1_27_11_i;
wire signed [`CalcTempBus]          temp_b1_27_12_r;
wire signed [`CalcTempBus]          temp_b1_27_12_i;
wire signed [`CalcTempBus]          temp_b1_27_13_r;
wire signed [`CalcTempBus]          temp_b1_27_13_i;
wire signed [`CalcTempBus]          temp_b1_27_14_r;
wire signed [`CalcTempBus]          temp_b1_27_14_i;
wire signed [`CalcTempBus]          temp_b1_27_15_r;
wire signed [`CalcTempBus]          temp_b1_27_15_i;
wire signed [`CalcTempBus]          temp_b1_27_16_r;
wire signed [`CalcTempBus]          temp_b1_27_16_i;
wire signed [`CalcTempBus]          temp_b1_27_17_r;
wire signed [`CalcTempBus]          temp_b1_27_17_i;
wire signed [`CalcTempBus]          temp_b1_27_18_r;
wire signed [`CalcTempBus]          temp_b1_27_18_i;
wire signed [`CalcTempBus]          temp_b1_27_19_r;
wire signed [`CalcTempBus]          temp_b1_27_19_i;
wire signed [`CalcTempBus]          temp_b1_27_20_r;
wire signed [`CalcTempBus]          temp_b1_27_20_i;
wire signed [`CalcTempBus]          temp_b1_27_21_r;
wire signed [`CalcTempBus]          temp_b1_27_21_i;
wire signed [`CalcTempBus]          temp_b1_27_22_r;
wire signed [`CalcTempBus]          temp_b1_27_22_i;
wire signed [`CalcTempBus]          temp_b1_27_23_r;
wire signed [`CalcTempBus]          temp_b1_27_23_i;
wire signed [`CalcTempBus]          temp_b1_27_24_r;
wire signed [`CalcTempBus]          temp_b1_27_24_i;
wire signed [`CalcTempBus]          temp_b1_27_25_r;
wire signed [`CalcTempBus]          temp_b1_27_25_i;
wire signed [`CalcTempBus]          temp_b1_27_26_r;
wire signed [`CalcTempBus]          temp_b1_27_26_i;
wire signed [`CalcTempBus]          temp_b1_27_27_r;
wire signed [`CalcTempBus]          temp_b1_27_27_i;
wire signed [`CalcTempBus]          temp_b1_27_28_r;
wire signed [`CalcTempBus]          temp_b1_27_28_i;
wire signed [`CalcTempBus]          temp_b1_27_29_r;
wire signed [`CalcTempBus]          temp_b1_27_29_i;
wire signed [`CalcTempBus]          temp_b1_27_30_r;
wire signed [`CalcTempBus]          temp_b1_27_30_i;
wire signed [`CalcTempBus]          temp_b1_27_31_r;
wire signed [`CalcTempBus]          temp_b1_27_31_i;
wire signed [`CalcTempBus]          temp_b1_27_32_r;
wire signed [`CalcTempBus]          temp_b1_27_32_i;
wire signed [`CalcTempBus]          temp_b1_28_1_r;
wire signed [`CalcTempBus]          temp_b1_28_1_i;
wire signed [`CalcTempBus]          temp_b1_28_2_r;
wire signed [`CalcTempBus]          temp_b1_28_2_i;
wire signed [`CalcTempBus]          temp_b1_28_3_r;
wire signed [`CalcTempBus]          temp_b1_28_3_i;
wire signed [`CalcTempBus]          temp_b1_28_4_r;
wire signed [`CalcTempBus]          temp_b1_28_4_i;
wire signed [`CalcTempBus]          temp_b1_28_5_r;
wire signed [`CalcTempBus]          temp_b1_28_5_i;
wire signed [`CalcTempBus]          temp_b1_28_6_r;
wire signed [`CalcTempBus]          temp_b1_28_6_i;
wire signed [`CalcTempBus]          temp_b1_28_7_r;
wire signed [`CalcTempBus]          temp_b1_28_7_i;
wire signed [`CalcTempBus]          temp_b1_28_8_r;
wire signed [`CalcTempBus]          temp_b1_28_8_i;
wire signed [`CalcTempBus]          temp_b1_28_9_r;
wire signed [`CalcTempBus]          temp_b1_28_9_i;
wire signed [`CalcTempBus]          temp_b1_28_10_r;
wire signed [`CalcTempBus]          temp_b1_28_10_i;
wire signed [`CalcTempBus]          temp_b1_28_11_r;
wire signed [`CalcTempBus]          temp_b1_28_11_i;
wire signed [`CalcTempBus]          temp_b1_28_12_r;
wire signed [`CalcTempBus]          temp_b1_28_12_i;
wire signed [`CalcTempBus]          temp_b1_28_13_r;
wire signed [`CalcTempBus]          temp_b1_28_13_i;
wire signed [`CalcTempBus]          temp_b1_28_14_r;
wire signed [`CalcTempBus]          temp_b1_28_14_i;
wire signed [`CalcTempBus]          temp_b1_28_15_r;
wire signed [`CalcTempBus]          temp_b1_28_15_i;
wire signed [`CalcTempBus]          temp_b1_28_16_r;
wire signed [`CalcTempBus]          temp_b1_28_16_i;
wire signed [`CalcTempBus]          temp_b1_28_17_r;
wire signed [`CalcTempBus]          temp_b1_28_17_i;
wire signed [`CalcTempBus]          temp_b1_28_18_r;
wire signed [`CalcTempBus]          temp_b1_28_18_i;
wire signed [`CalcTempBus]          temp_b1_28_19_r;
wire signed [`CalcTempBus]          temp_b1_28_19_i;
wire signed [`CalcTempBus]          temp_b1_28_20_r;
wire signed [`CalcTempBus]          temp_b1_28_20_i;
wire signed [`CalcTempBus]          temp_b1_28_21_r;
wire signed [`CalcTempBus]          temp_b1_28_21_i;
wire signed [`CalcTempBus]          temp_b1_28_22_r;
wire signed [`CalcTempBus]          temp_b1_28_22_i;
wire signed [`CalcTempBus]          temp_b1_28_23_r;
wire signed [`CalcTempBus]          temp_b1_28_23_i;
wire signed [`CalcTempBus]          temp_b1_28_24_r;
wire signed [`CalcTempBus]          temp_b1_28_24_i;
wire signed [`CalcTempBus]          temp_b1_28_25_r;
wire signed [`CalcTempBus]          temp_b1_28_25_i;
wire signed [`CalcTempBus]          temp_b1_28_26_r;
wire signed [`CalcTempBus]          temp_b1_28_26_i;
wire signed [`CalcTempBus]          temp_b1_28_27_r;
wire signed [`CalcTempBus]          temp_b1_28_27_i;
wire signed [`CalcTempBus]          temp_b1_28_28_r;
wire signed [`CalcTempBus]          temp_b1_28_28_i;
wire signed [`CalcTempBus]          temp_b1_28_29_r;
wire signed [`CalcTempBus]          temp_b1_28_29_i;
wire signed [`CalcTempBus]          temp_b1_28_30_r;
wire signed [`CalcTempBus]          temp_b1_28_30_i;
wire signed [`CalcTempBus]          temp_b1_28_31_r;
wire signed [`CalcTempBus]          temp_b1_28_31_i;
wire signed [`CalcTempBus]          temp_b1_28_32_r;
wire signed [`CalcTempBus]          temp_b1_28_32_i;
wire signed [`CalcTempBus]          temp_b1_29_1_r;
wire signed [`CalcTempBus]          temp_b1_29_1_i;
wire signed [`CalcTempBus]          temp_b1_29_2_r;
wire signed [`CalcTempBus]          temp_b1_29_2_i;
wire signed [`CalcTempBus]          temp_b1_29_3_r;
wire signed [`CalcTempBus]          temp_b1_29_3_i;
wire signed [`CalcTempBus]          temp_b1_29_4_r;
wire signed [`CalcTempBus]          temp_b1_29_4_i;
wire signed [`CalcTempBus]          temp_b1_29_5_r;
wire signed [`CalcTempBus]          temp_b1_29_5_i;
wire signed [`CalcTempBus]          temp_b1_29_6_r;
wire signed [`CalcTempBus]          temp_b1_29_6_i;
wire signed [`CalcTempBus]          temp_b1_29_7_r;
wire signed [`CalcTempBus]          temp_b1_29_7_i;
wire signed [`CalcTempBus]          temp_b1_29_8_r;
wire signed [`CalcTempBus]          temp_b1_29_8_i;
wire signed [`CalcTempBus]          temp_b1_29_9_r;
wire signed [`CalcTempBus]          temp_b1_29_9_i;
wire signed [`CalcTempBus]          temp_b1_29_10_r;
wire signed [`CalcTempBus]          temp_b1_29_10_i;
wire signed [`CalcTempBus]          temp_b1_29_11_r;
wire signed [`CalcTempBus]          temp_b1_29_11_i;
wire signed [`CalcTempBus]          temp_b1_29_12_r;
wire signed [`CalcTempBus]          temp_b1_29_12_i;
wire signed [`CalcTempBus]          temp_b1_29_13_r;
wire signed [`CalcTempBus]          temp_b1_29_13_i;
wire signed [`CalcTempBus]          temp_b1_29_14_r;
wire signed [`CalcTempBus]          temp_b1_29_14_i;
wire signed [`CalcTempBus]          temp_b1_29_15_r;
wire signed [`CalcTempBus]          temp_b1_29_15_i;
wire signed [`CalcTempBus]          temp_b1_29_16_r;
wire signed [`CalcTempBus]          temp_b1_29_16_i;
wire signed [`CalcTempBus]          temp_b1_29_17_r;
wire signed [`CalcTempBus]          temp_b1_29_17_i;
wire signed [`CalcTempBus]          temp_b1_29_18_r;
wire signed [`CalcTempBus]          temp_b1_29_18_i;
wire signed [`CalcTempBus]          temp_b1_29_19_r;
wire signed [`CalcTempBus]          temp_b1_29_19_i;
wire signed [`CalcTempBus]          temp_b1_29_20_r;
wire signed [`CalcTempBus]          temp_b1_29_20_i;
wire signed [`CalcTempBus]          temp_b1_29_21_r;
wire signed [`CalcTempBus]          temp_b1_29_21_i;
wire signed [`CalcTempBus]          temp_b1_29_22_r;
wire signed [`CalcTempBus]          temp_b1_29_22_i;
wire signed [`CalcTempBus]          temp_b1_29_23_r;
wire signed [`CalcTempBus]          temp_b1_29_23_i;
wire signed [`CalcTempBus]          temp_b1_29_24_r;
wire signed [`CalcTempBus]          temp_b1_29_24_i;
wire signed [`CalcTempBus]          temp_b1_29_25_r;
wire signed [`CalcTempBus]          temp_b1_29_25_i;
wire signed [`CalcTempBus]          temp_b1_29_26_r;
wire signed [`CalcTempBus]          temp_b1_29_26_i;
wire signed [`CalcTempBus]          temp_b1_29_27_r;
wire signed [`CalcTempBus]          temp_b1_29_27_i;
wire signed [`CalcTempBus]          temp_b1_29_28_r;
wire signed [`CalcTempBus]          temp_b1_29_28_i;
wire signed [`CalcTempBus]          temp_b1_29_29_r;
wire signed [`CalcTempBus]          temp_b1_29_29_i;
wire signed [`CalcTempBus]          temp_b1_29_30_r;
wire signed [`CalcTempBus]          temp_b1_29_30_i;
wire signed [`CalcTempBus]          temp_b1_29_31_r;
wire signed [`CalcTempBus]          temp_b1_29_31_i;
wire signed [`CalcTempBus]          temp_b1_29_32_r;
wire signed [`CalcTempBus]          temp_b1_29_32_i;
wire signed [`CalcTempBus]          temp_b1_30_1_r;
wire signed [`CalcTempBus]          temp_b1_30_1_i;
wire signed [`CalcTempBus]          temp_b1_30_2_r;
wire signed [`CalcTempBus]          temp_b1_30_2_i;
wire signed [`CalcTempBus]          temp_b1_30_3_r;
wire signed [`CalcTempBus]          temp_b1_30_3_i;
wire signed [`CalcTempBus]          temp_b1_30_4_r;
wire signed [`CalcTempBus]          temp_b1_30_4_i;
wire signed [`CalcTempBus]          temp_b1_30_5_r;
wire signed [`CalcTempBus]          temp_b1_30_5_i;
wire signed [`CalcTempBus]          temp_b1_30_6_r;
wire signed [`CalcTempBus]          temp_b1_30_6_i;
wire signed [`CalcTempBus]          temp_b1_30_7_r;
wire signed [`CalcTempBus]          temp_b1_30_7_i;
wire signed [`CalcTempBus]          temp_b1_30_8_r;
wire signed [`CalcTempBus]          temp_b1_30_8_i;
wire signed [`CalcTempBus]          temp_b1_30_9_r;
wire signed [`CalcTempBus]          temp_b1_30_9_i;
wire signed [`CalcTempBus]          temp_b1_30_10_r;
wire signed [`CalcTempBus]          temp_b1_30_10_i;
wire signed [`CalcTempBus]          temp_b1_30_11_r;
wire signed [`CalcTempBus]          temp_b1_30_11_i;
wire signed [`CalcTempBus]          temp_b1_30_12_r;
wire signed [`CalcTempBus]          temp_b1_30_12_i;
wire signed [`CalcTempBus]          temp_b1_30_13_r;
wire signed [`CalcTempBus]          temp_b1_30_13_i;
wire signed [`CalcTempBus]          temp_b1_30_14_r;
wire signed [`CalcTempBus]          temp_b1_30_14_i;
wire signed [`CalcTempBus]          temp_b1_30_15_r;
wire signed [`CalcTempBus]          temp_b1_30_15_i;
wire signed [`CalcTempBus]          temp_b1_30_16_r;
wire signed [`CalcTempBus]          temp_b1_30_16_i;
wire signed [`CalcTempBus]          temp_b1_30_17_r;
wire signed [`CalcTempBus]          temp_b1_30_17_i;
wire signed [`CalcTempBus]          temp_b1_30_18_r;
wire signed [`CalcTempBus]          temp_b1_30_18_i;
wire signed [`CalcTempBus]          temp_b1_30_19_r;
wire signed [`CalcTempBus]          temp_b1_30_19_i;
wire signed [`CalcTempBus]          temp_b1_30_20_r;
wire signed [`CalcTempBus]          temp_b1_30_20_i;
wire signed [`CalcTempBus]          temp_b1_30_21_r;
wire signed [`CalcTempBus]          temp_b1_30_21_i;
wire signed [`CalcTempBus]          temp_b1_30_22_r;
wire signed [`CalcTempBus]          temp_b1_30_22_i;
wire signed [`CalcTempBus]          temp_b1_30_23_r;
wire signed [`CalcTempBus]          temp_b1_30_23_i;
wire signed [`CalcTempBus]          temp_b1_30_24_r;
wire signed [`CalcTempBus]          temp_b1_30_24_i;
wire signed [`CalcTempBus]          temp_b1_30_25_r;
wire signed [`CalcTempBus]          temp_b1_30_25_i;
wire signed [`CalcTempBus]          temp_b1_30_26_r;
wire signed [`CalcTempBus]          temp_b1_30_26_i;
wire signed [`CalcTempBus]          temp_b1_30_27_r;
wire signed [`CalcTempBus]          temp_b1_30_27_i;
wire signed [`CalcTempBus]          temp_b1_30_28_r;
wire signed [`CalcTempBus]          temp_b1_30_28_i;
wire signed [`CalcTempBus]          temp_b1_30_29_r;
wire signed [`CalcTempBus]          temp_b1_30_29_i;
wire signed [`CalcTempBus]          temp_b1_30_30_r;
wire signed [`CalcTempBus]          temp_b1_30_30_i;
wire signed [`CalcTempBus]          temp_b1_30_31_r;
wire signed [`CalcTempBus]          temp_b1_30_31_i;
wire signed [`CalcTempBus]          temp_b1_30_32_r;
wire signed [`CalcTempBus]          temp_b1_30_32_i;
wire signed [`CalcTempBus]          temp_b1_31_1_r;
wire signed [`CalcTempBus]          temp_b1_31_1_i;
wire signed [`CalcTempBus]          temp_b1_31_2_r;
wire signed [`CalcTempBus]          temp_b1_31_2_i;
wire signed [`CalcTempBus]          temp_b1_31_3_r;
wire signed [`CalcTempBus]          temp_b1_31_3_i;
wire signed [`CalcTempBus]          temp_b1_31_4_r;
wire signed [`CalcTempBus]          temp_b1_31_4_i;
wire signed [`CalcTempBus]          temp_b1_31_5_r;
wire signed [`CalcTempBus]          temp_b1_31_5_i;
wire signed [`CalcTempBus]          temp_b1_31_6_r;
wire signed [`CalcTempBus]          temp_b1_31_6_i;
wire signed [`CalcTempBus]          temp_b1_31_7_r;
wire signed [`CalcTempBus]          temp_b1_31_7_i;
wire signed [`CalcTempBus]          temp_b1_31_8_r;
wire signed [`CalcTempBus]          temp_b1_31_8_i;
wire signed [`CalcTempBus]          temp_b1_31_9_r;
wire signed [`CalcTempBus]          temp_b1_31_9_i;
wire signed [`CalcTempBus]          temp_b1_31_10_r;
wire signed [`CalcTempBus]          temp_b1_31_10_i;
wire signed [`CalcTempBus]          temp_b1_31_11_r;
wire signed [`CalcTempBus]          temp_b1_31_11_i;
wire signed [`CalcTempBus]          temp_b1_31_12_r;
wire signed [`CalcTempBus]          temp_b1_31_12_i;
wire signed [`CalcTempBus]          temp_b1_31_13_r;
wire signed [`CalcTempBus]          temp_b1_31_13_i;
wire signed [`CalcTempBus]          temp_b1_31_14_r;
wire signed [`CalcTempBus]          temp_b1_31_14_i;
wire signed [`CalcTempBus]          temp_b1_31_15_r;
wire signed [`CalcTempBus]          temp_b1_31_15_i;
wire signed [`CalcTempBus]          temp_b1_31_16_r;
wire signed [`CalcTempBus]          temp_b1_31_16_i;
wire signed [`CalcTempBus]          temp_b1_31_17_r;
wire signed [`CalcTempBus]          temp_b1_31_17_i;
wire signed [`CalcTempBus]          temp_b1_31_18_r;
wire signed [`CalcTempBus]          temp_b1_31_18_i;
wire signed [`CalcTempBus]          temp_b1_31_19_r;
wire signed [`CalcTempBus]          temp_b1_31_19_i;
wire signed [`CalcTempBus]          temp_b1_31_20_r;
wire signed [`CalcTempBus]          temp_b1_31_20_i;
wire signed [`CalcTempBus]          temp_b1_31_21_r;
wire signed [`CalcTempBus]          temp_b1_31_21_i;
wire signed [`CalcTempBus]          temp_b1_31_22_r;
wire signed [`CalcTempBus]          temp_b1_31_22_i;
wire signed [`CalcTempBus]          temp_b1_31_23_r;
wire signed [`CalcTempBus]          temp_b1_31_23_i;
wire signed [`CalcTempBus]          temp_b1_31_24_r;
wire signed [`CalcTempBus]          temp_b1_31_24_i;
wire signed [`CalcTempBus]          temp_b1_31_25_r;
wire signed [`CalcTempBus]          temp_b1_31_25_i;
wire signed [`CalcTempBus]          temp_b1_31_26_r;
wire signed [`CalcTempBus]          temp_b1_31_26_i;
wire signed [`CalcTempBus]          temp_b1_31_27_r;
wire signed [`CalcTempBus]          temp_b1_31_27_i;
wire signed [`CalcTempBus]          temp_b1_31_28_r;
wire signed [`CalcTempBus]          temp_b1_31_28_i;
wire signed [`CalcTempBus]          temp_b1_31_29_r;
wire signed [`CalcTempBus]          temp_b1_31_29_i;
wire signed [`CalcTempBus]          temp_b1_31_30_r;
wire signed [`CalcTempBus]          temp_b1_31_30_i;
wire signed [`CalcTempBus]          temp_b1_31_31_r;
wire signed [`CalcTempBus]          temp_b1_31_31_i;
wire signed [`CalcTempBus]          temp_b1_31_32_r;
wire signed [`CalcTempBus]          temp_b1_31_32_i;
wire signed [`CalcTempBus]          temp_b1_32_1_r;
wire signed [`CalcTempBus]          temp_b1_32_1_i;
wire signed [`CalcTempBus]          temp_b1_32_2_r;
wire signed [`CalcTempBus]          temp_b1_32_2_i;
wire signed [`CalcTempBus]          temp_b1_32_3_r;
wire signed [`CalcTempBus]          temp_b1_32_3_i;
wire signed [`CalcTempBus]          temp_b1_32_4_r;
wire signed [`CalcTempBus]          temp_b1_32_4_i;
wire signed [`CalcTempBus]          temp_b1_32_5_r;
wire signed [`CalcTempBus]          temp_b1_32_5_i;
wire signed [`CalcTempBus]          temp_b1_32_6_r;
wire signed [`CalcTempBus]          temp_b1_32_6_i;
wire signed [`CalcTempBus]          temp_b1_32_7_r;
wire signed [`CalcTempBus]          temp_b1_32_7_i;
wire signed [`CalcTempBus]          temp_b1_32_8_r;
wire signed [`CalcTempBus]          temp_b1_32_8_i;
wire signed [`CalcTempBus]          temp_b1_32_9_r;
wire signed [`CalcTempBus]          temp_b1_32_9_i;
wire signed [`CalcTempBus]          temp_b1_32_10_r;
wire signed [`CalcTempBus]          temp_b1_32_10_i;
wire signed [`CalcTempBus]          temp_b1_32_11_r;
wire signed [`CalcTempBus]          temp_b1_32_11_i;
wire signed [`CalcTempBus]          temp_b1_32_12_r;
wire signed [`CalcTempBus]          temp_b1_32_12_i;
wire signed [`CalcTempBus]          temp_b1_32_13_r;
wire signed [`CalcTempBus]          temp_b1_32_13_i;
wire signed [`CalcTempBus]          temp_b1_32_14_r;
wire signed [`CalcTempBus]          temp_b1_32_14_i;
wire signed [`CalcTempBus]          temp_b1_32_15_r;
wire signed [`CalcTempBus]          temp_b1_32_15_i;
wire signed [`CalcTempBus]          temp_b1_32_16_r;
wire signed [`CalcTempBus]          temp_b1_32_16_i;
wire signed [`CalcTempBus]          temp_b1_32_17_r;
wire signed [`CalcTempBus]          temp_b1_32_17_i;
wire signed [`CalcTempBus]          temp_b1_32_18_r;
wire signed [`CalcTempBus]          temp_b1_32_18_i;
wire signed [`CalcTempBus]          temp_b1_32_19_r;
wire signed [`CalcTempBus]          temp_b1_32_19_i;
wire signed [`CalcTempBus]          temp_b1_32_20_r;
wire signed [`CalcTempBus]          temp_b1_32_20_i;
wire signed [`CalcTempBus]          temp_b1_32_21_r;
wire signed [`CalcTempBus]          temp_b1_32_21_i;
wire signed [`CalcTempBus]          temp_b1_32_22_r;
wire signed [`CalcTempBus]          temp_b1_32_22_i;
wire signed [`CalcTempBus]          temp_b1_32_23_r;
wire signed [`CalcTempBus]          temp_b1_32_23_i;
wire signed [`CalcTempBus]          temp_b1_32_24_r;
wire signed [`CalcTempBus]          temp_b1_32_24_i;
wire signed [`CalcTempBus]          temp_b1_32_25_r;
wire signed [`CalcTempBus]          temp_b1_32_25_i;
wire signed [`CalcTempBus]          temp_b1_32_26_r;
wire signed [`CalcTempBus]          temp_b1_32_26_i;
wire signed [`CalcTempBus]          temp_b1_32_27_r;
wire signed [`CalcTempBus]          temp_b1_32_27_i;
wire signed [`CalcTempBus]          temp_b1_32_28_r;
wire signed [`CalcTempBus]          temp_b1_32_28_i;
wire signed [`CalcTempBus]          temp_b1_32_29_r;
wire signed [`CalcTempBus]          temp_b1_32_29_i;
wire signed [`CalcTempBus]          temp_b1_32_30_r;
wire signed [`CalcTempBus]          temp_b1_32_30_i;
wire signed [`CalcTempBus]          temp_b1_32_31_r;
wire signed [`CalcTempBus]          temp_b1_32_31_i;
wire signed [`CalcTempBus]          temp_b1_32_32_r;
wire signed [`CalcTempBus]          temp_b1_32_32_i;
wire signed [`CalcTempBus]          temp_b2_1_1_r;
wire signed [`CalcTempBus]          temp_b2_1_1_i;
wire signed [`CalcTempBus]          temp_b2_1_2_r;
wire signed [`CalcTempBus]          temp_b2_1_2_i;
wire signed [`CalcTempBus]          temp_b2_1_3_r;
wire signed [`CalcTempBus]          temp_b2_1_3_i;
wire signed [`CalcTempBus]          temp_b2_1_4_r;
wire signed [`CalcTempBus]          temp_b2_1_4_i;
wire signed [`CalcTempBus]          temp_b2_1_5_r;
wire signed [`CalcTempBus]          temp_b2_1_5_i;
wire signed [`CalcTempBus]          temp_b2_1_6_r;
wire signed [`CalcTempBus]          temp_b2_1_6_i;
wire signed [`CalcTempBus]          temp_b2_1_7_r;
wire signed [`CalcTempBus]          temp_b2_1_7_i;
wire signed [`CalcTempBus]          temp_b2_1_8_r;
wire signed [`CalcTempBus]          temp_b2_1_8_i;
wire signed [`CalcTempBus]          temp_b2_1_9_r;
wire signed [`CalcTempBus]          temp_b2_1_9_i;
wire signed [`CalcTempBus]          temp_b2_1_10_r;
wire signed [`CalcTempBus]          temp_b2_1_10_i;
wire signed [`CalcTempBus]          temp_b2_1_11_r;
wire signed [`CalcTempBus]          temp_b2_1_11_i;
wire signed [`CalcTempBus]          temp_b2_1_12_r;
wire signed [`CalcTempBus]          temp_b2_1_12_i;
wire signed [`CalcTempBus]          temp_b2_1_13_r;
wire signed [`CalcTempBus]          temp_b2_1_13_i;
wire signed [`CalcTempBus]          temp_b2_1_14_r;
wire signed [`CalcTempBus]          temp_b2_1_14_i;
wire signed [`CalcTempBus]          temp_b2_1_15_r;
wire signed [`CalcTempBus]          temp_b2_1_15_i;
wire signed [`CalcTempBus]          temp_b2_1_16_r;
wire signed [`CalcTempBus]          temp_b2_1_16_i;
wire signed [`CalcTempBus]          temp_b2_1_17_r;
wire signed [`CalcTempBus]          temp_b2_1_17_i;
wire signed [`CalcTempBus]          temp_b2_1_18_r;
wire signed [`CalcTempBus]          temp_b2_1_18_i;
wire signed [`CalcTempBus]          temp_b2_1_19_r;
wire signed [`CalcTempBus]          temp_b2_1_19_i;
wire signed [`CalcTempBus]          temp_b2_1_20_r;
wire signed [`CalcTempBus]          temp_b2_1_20_i;
wire signed [`CalcTempBus]          temp_b2_1_21_r;
wire signed [`CalcTempBus]          temp_b2_1_21_i;
wire signed [`CalcTempBus]          temp_b2_1_22_r;
wire signed [`CalcTempBus]          temp_b2_1_22_i;
wire signed [`CalcTempBus]          temp_b2_1_23_r;
wire signed [`CalcTempBus]          temp_b2_1_23_i;
wire signed [`CalcTempBus]          temp_b2_1_24_r;
wire signed [`CalcTempBus]          temp_b2_1_24_i;
wire signed [`CalcTempBus]          temp_b2_1_25_r;
wire signed [`CalcTempBus]          temp_b2_1_25_i;
wire signed [`CalcTempBus]          temp_b2_1_26_r;
wire signed [`CalcTempBus]          temp_b2_1_26_i;
wire signed [`CalcTempBus]          temp_b2_1_27_r;
wire signed [`CalcTempBus]          temp_b2_1_27_i;
wire signed [`CalcTempBus]          temp_b2_1_28_r;
wire signed [`CalcTempBus]          temp_b2_1_28_i;
wire signed [`CalcTempBus]          temp_b2_1_29_r;
wire signed [`CalcTempBus]          temp_b2_1_29_i;
wire signed [`CalcTempBus]          temp_b2_1_30_r;
wire signed [`CalcTempBus]          temp_b2_1_30_i;
wire signed [`CalcTempBus]          temp_b2_1_31_r;
wire signed [`CalcTempBus]          temp_b2_1_31_i;
wire signed [`CalcTempBus]          temp_b2_1_32_r;
wire signed [`CalcTempBus]          temp_b2_1_32_i;
wire signed [`CalcTempBus]          temp_b2_2_1_r;
wire signed [`CalcTempBus]          temp_b2_2_1_i;
wire signed [`CalcTempBus]          temp_b2_2_2_r;
wire signed [`CalcTempBus]          temp_b2_2_2_i;
wire signed [`CalcTempBus]          temp_b2_2_3_r;
wire signed [`CalcTempBus]          temp_b2_2_3_i;
wire signed [`CalcTempBus]          temp_b2_2_4_r;
wire signed [`CalcTempBus]          temp_b2_2_4_i;
wire signed [`CalcTempBus]          temp_b2_2_5_r;
wire signed [`CalcTempBus]          temp_b2_2_5_i;
wire signed [`CalcTempBus]          temp_b2_2_6_r;
wire signed [`CalcTempBus]          temp_b2_2_6_i;
wire signed [`CalcTempBus]          temp_b2_2_7_r;
wire signed [`CalcTempBus]          temp_b2_2_7_i;
wire signed [`CalcTempBus]          temp_b2_2_8_r;
wire signed [`CalcTempBus]          temp_b2_2_8_i;
wire signed [`CalcTempBus]          temp_b2_2_9_r;
wire signed [`CalcTempBus]          temp_b2_2_9_i;
wire signed [`CalcTempBus]          temp_b2_2_10_r;
wire signed [`CalcTempBus]          temp_b2_2_10_i;
wire signed [`CalcTempBus]          temp_b2_2_11_r;
wire signed [`CalcTempBus]          temp_b2_2_11_i;
wire signed [`CalcTempBus]          temp_b2_2_12_r;
wire signed [`CalcTempBus]          temp_b2_2_12_i;
wire signed [`CalcTempBus]          temp_b2_2_13_r;
wire signed [`CalcTempBus]          temp_b2_2_13_i;
wire signed [`CalcTempBus]          temp_b2_2_14_r;
wire signed [`CalcTempBus]          temp_b2_2_14_i;
wire signed [`CalcTempBus]          temp_b2_2_15_r;
wire signed [`CalcTempBus]          temp_b2_2_15_i;
wire signed [`CalcTempBus]          temp_b2_2_16_r;
wire signed [`CalcTempBus]          temp_b2_2_16_i;
wire signed [`CalcTempBus]          temp_b2_2_17_r;
wire signed [`CalcTempBus]          temp_b2_2_17_i;
wire signed [`CalcTempBus]          temp_b2_2_18_r;
wire signed [`CalcTempBus]          temp_b2_2_18_i;
wire signed [`CalcTempBus]          temp_b2_2_19_r;
wire signed [`CalcTempBus]          temp_b2_2_19_i;
wire signed [`CalcTempBus]          temp_b2_2_20_r;
wire signed [`CalcTempBus]          temp_b2_2_20_i;
wire signed [`CalcTempBus]          temp_b2_2_21_r;
wire signed [`CalcTempBus]          temp_b2_2_21_i;
wire signed [`CalcTempBus]          temp_b2_2_22_r;
wire signed [`CalcTempBus]          temp_b2_2_22_i;
wire signed [`CalcTempBus]          temp_b2_2_23_r;
wire signed [`CalcTempBus]          temp_b2_2_23_i;
wire signed [`CalcTempBus]          temp_b2_2_24_r;
wire signed [`CalcTempBus]          temp_b2_2_24_i;
wire signed [`CalcTempBus]          temp_b2_2_25_r;
wire signed [`CalcTempBus]          temp_b2_2_25_i;
wire signed [`CalcTempBus]          temp_b2_2_26_r;
wire signed [`CalcTempBus]          temp_b2_2_26_i;
wire signed [`CalcTempBus]          temp_b2_2_27_r;
wire signed [`CalcTempBus]          temp_b2_2_27_i;
wire signed [`CalcTempBus]          temp_b2_2_28_r;
wire signed [`CalcTempBus]          temp_b2_2_28_i;
wire signed [`CalcTempBus]          temp_b2_2_29_r;
wire signed [`CalcTempBus]          temp_b2_2_29_i;
wire signed [`CalcTempBus]          temp_b2_2_30_r;
wire signed [`CalcTempBus]          temp_b2_2_30_i;
wire signed [`CalcTempBus]          temp_b2_2_31_r;
wire signed [`CalcTempBus]          temp_b2_2_31_i;
wire signed [`CalcTempBus]          temp_b2_2_32_r;
wire signed [`CalcTempBus]          temp_b2_2_32_i;
wire signed [`CalcTempBus]          temp_b2_3_1_r;
wire signed [`CalcTempBus]          temp_b2_3_1_i;
wire signed [`CalcTempBus]          temp_b2_3_2_r;
wire signed [`CalcTempBus]          temp_b2_3_2_i;
wire signed [`CalcTempBus]          temp_b2_3_3_r;
wire signed [`CalcTempBus]          temp_b2_3_3_i;
wire signed [`CalcTempBus]          temp_b2_3_4_r;
wire signed [`CalcTempBus]          temp_b2_3_4_i;
wire signed [`CalcTempBus]          temp_b2_3_5_r;
wire signed [`CalcTempBus]          temp_b2_3_5_i;
wire signed [`CalcTempBus]          temp_b2_3_6_r;
wire signed [`CalcTempBus]          temp_b2_3_6_i;
wire signed [`CalcTempBus]          temp_b2_3_7_r;
wire signed [`CalcTempBus]          temp_b2_3_7_i;
wire signed [`CalcTempBus]          temp_b2_3_8_r;
wire signed [`CalcTempBus]          temp_b2_3_8_i;
wire signed [`CalcTempBus]          temp_b2_3_9_r;
wire signed [`CalcTempBus]          temp_b2_3_9_i;
wire signed [`CalcTempBus]          temp_b2_3_10_r;
wire signed [`CalcTempBus]          temp_b2_3_10_i;
wire signed [`CalcTempBus]          temp_b2_3_11_r;
wire signed [`CalcTempBus]          temp_b2_3_11_i;
wire signed [`CalcTempBus]          temp_b2_3_12_r;
wire signed [`CalcTempBus]          temp_b2_3_12_i;
wire signed [`CalcTempBus]          temp_b2_3_13_r;
wire signed [`CalcTempBus]          temp_b2_3_13_i;
wire signed [`CalcTempBus]          temp_b2_3_14_r;
wire signed [`CalcTempBus]          temp_b2_3_14_i;
wire signed [`CalcTempBus]          temp_b2_3_15_r;
wire signed [`CalcTempBus]          temp_b2_3_15_i;
wire signed [`CalcTempBus]          temp_b2_3_16_r;
wire signed [`CalcTempBus]          temp_b2_3_16_i;
wire signed [`CalcTempBus]          temp_b2_3_17_r;
wire signed [`CalcTempBus]          temp_b2_3_17_i;
wire signed [`CalcTempBus]          temp_b2_3_18_r;
wire signed [`CalcTempBus]          temp_b2_3_18_i;
wire signed [`CalcTempBus]          temp_b2_3_19_r;
wire signed [`CalcTempBus]          temp_b2_3_19_i;
wire signed [`CalcTempBus]          temp_b2_3_20_r;
wire signed [`CalcTempBus]          temp_b2_3_20_i;
wire signed [`CalcTempBus]          temp_b2_3_21_r;
wire signed [`CalcTempBus]          temp_b2_3_21_i;
wire signed [`CalcTempBus]          temp_b2_3_22_r;
wire signed [`CalcTempBus]          temp_b2_3_22_i;
wire signed [`CalcTempBus]          temp_b2_3_23_r;
wire signed [`CalcTempBus]          temp_b2_3_23_i;
wire signed [`CalcTempBus]          temp_b2_3_24_r;
wire signed [`CalcTempBus]          temp_b2_3_24_i;
wire signed [`CalcTempBus]          temp_b2_3_25_r;
wire signed [`CalcTempBus]          temp_b2_3_25_i;
wire signed [`CalcTempBus]          temp_b2_3_26_r;
wire signed [`CalcTempBus]          temp_b2_3_26_i;
wire signed [`CalcTempBus]          temp_b2_3_27_r;
wire signed [`CalcTempBus]          temp_b2_3_27_i;
wire signed [`CalcTempBus]          temp_b2_3_28_r;
wire signed [`CalcTempBus]          temp_b2_3_28_i;
wire signed [`CalcTempBus]          temp_b2_3_29_r;
wire signed [`CalcTempBus]          temp_b2_3_29_i;
wire signed [`CalcTempBus]          temp_b2_3_30_r;
wire signed [`CalcTempBus]          temp_b2_3_30_i;
wire signed [`CalcTempBus]          temp_b2_3_31_r;
wire signed [`CalcTempBus]          temp_b2_3_31_i;
wire signed [`CalcTempBus]          temp_b2_3_32_r;
wire signed [`CalcTempBus]          temp_b2_3_32_i;
wire signed [`CalcTempBus]          temp_b2_4_1_r;
wire signed [`CalcTempBus]          temp_b2_4_1_i;
wire signed [`CalcTempBus]          temp_b2_4_2_r;
wire signed [`CalcTempBus]          temp_b2_4_2_i;
wire signed [`CalcTempBus]          temp_b2_4_3_r;
wire signed [`CalcTempBus]          temp_b2_4_3_i;
wire signed [`CalcTempBus]          temp_b2_4_4_r;
wire signed [`CalcTempBus]          temp_b2_4_4_i;
wire signed [`CalcTempBus]          temp_b2_4_5_r;
wire signed [`CalcTempBus]          temp_b2_4_5_i;
wire signed [`CalcTempBus]          temp_b2_4_6_r;
wire signed [`CalcTempBus]          temp_b2_4_6_i;
wire signed [`CalcTempBus]          temp_b2_4_7_r;
wire signed [`CalcTempBus]          temp_b2_4_7_i;
wire signed [`CalcTempBus]          temp_b2_4_8_r;
wire signed [`CalcTempBus]          temp_b2_4_8_i;
wire signed [`CalcTempBus]          temp_b2_4_9_r;
wire signed [`CalcTempBus]          temp_b2_4_9_i;
wire signed [`CalcTempBus]          temp_b2_4_10_r;
wire signed [`CalcTempBus]          temp_b2_4_10_i;
wire signed [`CalcTempBus]          temp_b2_4_11_r;
wire signed [`CalcTempBus]          temp_b2_4_11_i;
wire signed [`CalcTempBus]          temp_b2_4_12_r;
wire signed [`CalcTempBus]          temp_b2_4_12_i;
wire signed [`CalcTempBus]          temp_b2_4_13_r;
wire signed [`CalcTempBus]          temp_b2_4_13_i;
wire signed [`CalcTempBus]          temp_b2_4_14_r;
wire signed [`CalcTempBus]          temp_b2_4_14_i;
wire signed [`CalcTempBus]          temp_b2_4_15_r;
wire signed [`CalcTempBus]          temp_b2_4_15_i;
wire signed [`CalcTempBus]          temp_b2_4_16_r;
wire signed [`CalcTempBus]          temp_b2_4_16_i;
wire signed [`CalcTempBus]          temp_b2_4_17_r;
wire signed [`CalcTempBus]          temp_b2_4_17_i;
wire signed [`CalcTempBus]          temp_b2_4_18_r;
wire signed [`CalcTempBus]          temp_b2_4_18_i;
wire signed [`CalcTempBus]          temp_b2_4_19_r;
wire signed [`CalcTempBus]          temp_b2_4_19_i;
wire signed [`CalcTempBus]          temp_b2_4_20_r;
wire signed [`CalcTempBus]          temp_b2_4_20_i;
wire signed [`CalcTempBus]          temp_b2_4_21_r;
wire signed [`CalcTempBus]          temp_b2_4_21_i;
wire signed [`CalcTempBus]          temp_b2_4_22_r;
wire signed [`CalcTempBus]          temp_b2_4_22_i;
wire signed [`CalcTempBus]          temp_b2_4_23_r;
wire signed [`CalcTempBus]          temp_b2_4_23_i;
wire signed [`CalcTempBus]          temp_b2_4_24_r;
wire signed [`CalcTempBus]          temp_b2_4_24_i;
wire signed [`CalcTempBus]          temp_b2_4_25_r;
wire signed [`CalcTempBus]          temp_b2_4_25_i;
wire signed [`CalcTempBus]          temp_b2_4_26_r;
wire signed [`CalcTempBus]          temp_b2_4_26_i;
wire signed [`CalcTempBus]          temp_b2_4_27_r;
wire signed [`CalcTempBus]          temp_b2_4_27_i;
wire signed [`CalcTempBus]          temp_b2_4_28_r;
wire signed [`CalcTempBus]          temp_b2_4_28_i;
wire signed [`CalcTempBus]          temp_b2_4_29_r;
wire signed [`CalcTempBus]          temp_b2_4_29_i;
wire signed [`CalcTempBus]          temp_b2_4_30_r;
wire signed [`CalcTempBus]          temp_b2_4_30_i;
wire signed [`CalcTempBus]          temp_b2_4_31_r;
wire signed [`CalcTempBus]          temp_b2_4_31_i;
wire signed [`CalcTempBus]          temp_b2_4_32_r;
wire signed [`CalcTempBus]          temp_b2_4_32_i;
wire signed [`CalcTempBus]          temp_b2_5_1_r;
wire signed [`CalcTempBus]          temp_b2_5_1_i;
wire signed [`CalcTempBus]          temp_b2_5_2_r;
wire signed [`CalcTempBus]          temp_b2_5_2_i;
wire signed [`CalcTempBus]          temp_b2_5_3_r;
wire signed [`CalcTempBus]          temp_b2_5_3_i;
wire signed [`CalcTempBus]          temp_b2_5_4_r;
wire signed [`CalcTempBus]          temp_b2_5_4_i;
wire signed [`CalcTempBus]          temp_b2_5_5_r;
wire signed [`CalcTempBus]          temp_b2_5_5_i;
wire signed [`CalcTempBus]          temp_b2_5_6_r;
wire signed [`CalcTempBus]          temp_b2_5_6_i;
wire signed [`CalcTempBus]          temp_b2_5_7_r;
wire signed [`CalcTempBus]          temp_b2_5_7_i;
wire signed [`CalcTempBus]          temp_b2_5_8_r;
wire signed [`CalcTempBus]          temp_b2_5_8_i;
wire signed [`CalcTempBus]          temp_b2_5_9_r;
wire signed [`CalcTempBus]          temp_b2_5_9_i;
wire signed [`CalcTempBus]          temp_b2_5_10_r;
wire signed [`CalcTempBus]          temp_b2_5_10_i;
wire signed [`CalcTempBus]          temp_b2_5_11_r;
wire signed [`CalcTempBus]          temp_b2_5_11_i;
wire signed [`CalcTempBus]          temp_b2_5_12_r;
wire signed [`CalcTempBus]          temp_b2_5_12_i;
wire signed [`CalcTempBus]          temp_b2_5_13_r;
wire signed [`CalcTempBus]          temp_b2_5_13_i;
wire signed [`CalcTempBus]          temp_b2_5_14_r;
wire signed [`CalcTempBus]          temp_b2_5_14_i;
wire signed [`CalcTempBus]          temp_b2_5_15_r;
wire signed [`CalcTempBus]          temp_b2_5_15_i;
wire signed [`CalcTempBus]          temp_b2_5_16_r;
wire signed [`CalcTempBus]          temp_b2_5_16_i;
wire signed [`CalcTempBus]          temp_b2_5_17_r;
wire signed [`CalcTempBus]          temp_b2_5_17_i;
wire signed [`CalcTempBus]          temp_b2_5_18_r;
wire signed [`CalcTempBus]          temp_b2_5_18_i;
wire signed [`CalcTempBus]          temp_b2_5_19_r;
wire signed [`CalcTempBus]          temp_b2_5_19_i;
wire signed [`CalcTempBus]          temp_b2_5_20_r;
wire signed [`CalcTempBus]          temp_b2_5_20_i;
wire signed [`CalcTempBus]          temp_b2_5_21_r;
wire signed [`CalcTempBus]          temp_b2_5_21_i;
wire signed [`CalcTempBus]          temp_b2_5_22_r;
wire signed [`CalcTempBus]          temp_b2_5_22_i;
wire signed [`CalcTempBus]          temp_b2_5_23_r;
wire signed [`CalcTempBus]          temp_b2_5_23_i;
wire signed [`CalcTempBus]          temp_b2_5_24_r;
wire signed [`CalcTempBus]          temp_b2_5_24_i;
wire signed [`CalcTempBus]          temp_b2_5_25_r;
wire signed [`CalcTempBus]          temp_b2_5_25_i;
wire signed [`CalcTempBus]          temp_b2_5_26_r;
wire signed [`CalcTempBus]          temp_b2_5_26_i;
wire signed [`CalcTempBus]          temp_b2_5_27_r;
wire signed [`CalcTempBus]          temp_b2_5_27_i;
wire signed [`CalcTempBus]          temp_b2_5_28_r;
wire signed [`CalcTempBus]          temp_b2_5_28_i;
wire signed [`CalcTempBus]          temp_b2_5_29_r;
wire signed [`CalcTempBus]          temp_b2_5_29_i;
wire signed [`CalcTempBus]          temp_b2_5_30_r;
wire signed [`CalcTempBus]          temp_b2_5_30_i;
wire signed [`CalcTempBus]          temp_b2_5_31_r;
wire signed [`CalcTempBus]          temp_b2_5_31_i;
wire signed [`CalcTempBus]          temp_b2_5_32_r;
wire signed [`CalcTempBus]          temp_b2_5_32_i;
wire signed [`CalcTempBus]          temp_b2_6_1_r;
wire signed [`CalcTempBus]          temp_b2_6_1_i;
wire signed [`CalcTempBus]          temp_b2_6_2_r;
wire signed [`CalcTempBus]          temp_b2_6_2_i;
wire signed [`CalcTempBus]          temp_b2_6_3_r;
wire signed [`CalcTempBus]          temp_b2_6_3_i;
wire signed [`CalcTempBus]          temp_b2_6_4_r;
wire signed [`CalcTempBus]          temp_b2_6_4_i;
wire signed [`CalcTempBus]          temp_b2_6_5_r;
wire signed [`CalcTempBus]          temp_b2_6_5_i;
wire signed [`CalcTempBus]          temp_b2_6_6_r;
wire signed [`CalcTempBus]          temp_b2_6_6_i;
wire signed [`CalcTempBus]          temp_b2_6_7_r;
wire signed [`CalcTempBus]          temp_b2_6_7_i;
wire signed [`CalcTempBus]          temp_b2_6_8_r;
wire signed [`CalcTempBus]          temp_b2_6_8_i;
wire signed [`CalcTempBus]          temp_b2_6_9_r;
wire signed [`CalcTempBus]          temp_b2_6_9_i;
wire signed [`CalcTempBus]          temp_b2_6_10_r;
wire signed [`CalcTempBus]          temp_b2_6_10_i;
wire signed [`CalcTempBus]          temp_b2_6_11_r;
wire signed [`CalcTempBus]          temp_b2_6_11_i;
wire signed [`CalcTempBus]          temp_b2_6_12_r;
wire signed [`CalcTempBus]          temp_b2_6_12_i;
wire signed [`CalcTempBus]          temp_b2_6_13_r;
wire signed [`CalcTempBus]          temp_b2_6_13_i;
wire signed [`CalcTempBus]          temp_b2_6_14_r;
wire signed [`CalcTempBus]          temp_b2_6_14_i;
wire signed [`CalcTempBus]          temp_b2_6_15_r;
wire signed [`CalcTempBus]          temp_b2_6_15_i;
wire signed [`CalcTempBus]          temp_b2_6_16_r;
wire signed [`CalcTempBus]          temp_b2_6_16_i;
wire signed [`CalcTempBus]          temp_b2_6_17_r;
wire signed [`CalcTempBus]          temp_b2_6_17_i;
wire signed [`CalcTempBus]          temp_b2_6_18_r;
wire signed [`CalcTempBus]          temp_b2_6_18_i;
wire signed [`CalcTempBus]          temp_b2_6_19_r;
wire signed [`CalcTempBus]          temp_b2_6_19_i;
wire signed [`CalcTempBus]          temp_b2_6_20_r;
wire signed [`CalcTempBus]          temp_b2_6_20_i;
wire signed [`CalcTempBus]          temp_b2_6_21_r;
wire signed [`CalcTempBus]          temp_b2_6_21_i;
wire signed [`CalcTempBus]          temp_b2_6_22_r;
wire signed [`CalcTempBus]          temp_b2_6_22_i;
wire signed [`CalcTempBus]          temp_b2_6_23_r;
wire signed [`CalcTempBus]          temp_b2_6_23_i;
wire signed [`CalcTempBus]          temp_b2_6_24_r;
wire signed [`CalcTempBus]          temp_b2_6_24_i;
wire signed [`CalcTempBus]          temp_b2_6_25_r;
wire signed [`CalcTempBus]          temp_b2_6_25_i;
wire signed [`CalcTempBus]          temp_b2_6_26_r;
wire signed [`CalcTempBus]          temp_b2_6_26_i;
wire signed [`CalcTempBus]          temp_b2_6_27_r;
wire signed [`CalcTempBus]          temp_b2_6_27_i;
wire signed [`CalcTempBus]          temp_b2_6_28_r;
wire signed [`CalcTempBus]          temp_b2_6_28_i;
wire signed [`CalcTempBus]          temp_b2_6_29_r;
wire signed [`CalcTempBus]          temp_b2_6_29_i;
wire signed [`CalcTempBus]          temp_b2_6_30_r;
wire signed [`CalcTempBus]          temp_b2_6_30_i;
wire signed [`CalcTempBus]          temp_b2_6_31_r;
wire signed [`CalcTempBus]          temp_b2_6_31_i;
wire signed [`CalcTempBus]          temp_b2_6_32_r;
wire signed [`CalcTempBus]          temp_b2_6_32_i;
wire signed [`CalcTempBus]          temp_b2_7_1_r;
wire signed [`CalcTempBus]          temp_b2_7_1_i;
wire signed [`CalcTempBus]          temp_b2_7_2_r;
wire signed [`CalcTempBus]          temp_b2_7_2_i;
wire signed [`CalcTempBus]          temp_b2_7_3_r;
wire signed [`CalcTempBus]          temp_b2_7_3_i;
wire signed [`CalcTempBus]          temp_b2_7_4_r;
wire signed [`CalcTempBus]          temp_b2_7_4_i;
wire signed [`CalcTempBus]          temp_b2_7_5_r;
wire signed [`CalcTempBus]          temp_b2_7_5_i;
wire signed [`CalcTempBus]          temp_b2_7_6_r;
wire signed [`CalcTempBus]          temp_b2_7_6_i;
wire signed [`CalcTempBus]          temp_b2_7_7_r;
wire signed [`CalcTempBus]          temp_b2_7_7_i;
wire signed [`CalcTempBus]          temp_b2_7_8_r;
wire signed [`CalcTempBus]          temp_b2_7_8_i;
wire signed [`CalcTempBus]          temp_b2_7_9_r;
wire signed [`CalcTempBus]          temp_b2_7_9_i;
wire signed [`CalcTempBus]          temp_b2_7_10_r;
wire signed [`CalcTempBus]          temp_b2_7_10_i;
wire signed [`CalcTempBus]          temp_b2_7_11_r;
wire signed [`CalcTempBus]          temp_b2_7_11_i;
wire signed [`CalcTempBus]          temp_b2_7_12_r;
wire signed [`CalcTempBus]          temp_b2_7_12_i;
wire signed [`CalcTempBus]          temp_b2_7_13_r;
wire signed [`CalcTempBus]          temp_b2_7_13_i;
wire signed [`CalcTempBus]          temp_b2_7_14_r;
wire signed [`CalcTempBus]          temp_b2_7_14_i;
wire signed [`CalcTempBus]          temp_b2_7_15_r;
wire signed [`CalcTempBus]          temp_b2_7_15_i;
wire signed [`CalcTempBus]          temp_b2_7_16_r;
wire signed [`CalcTempBus]          temp_b2_7_16_i;
wire signed [`CalcTempBus]          temp_b2_7_17_r;
wire signed [`CalcTempBus]          temp_b2_7_17_i;
wire signed [`CalcTempBus]          temp_b2_7_18_r;
wire signed [`CalcTempBus]          temp_b2_7_18_i;
wire signed [`CalcTempBus]          temp_b2_7_19_r;
wire signed [`CalcTempBus]          temp_b2_7_19_i;
wire signed [`CalcTempBus]          temp_b2_7_20_r;
wire signed [`CalcTempBus]          temp_b2_7_20_i;
wire signed [`CalcTempBus]          temp_b2_7_21_r;
wire signed [`CalcTempBus]          temp_b2_7_21_i;
wire signed [`CalcTempBus]          temp_b2_7_22_r;
wire signed [`CalcTempBus]          temp_b2_7_22_i;
wire signed [`CalcTempBus]          temp_b2_7_23_r;
wire signed [`CalcTempBus]          temp_b2_7_23_i;
wire signed [`CalcTempBus]          temp_b2_7_24_r;
wire signed [`CalcTempBus]          temp_b2_7_24_i;
wire signed [`CalcTempBus]          temp_b2_7_25_r;
wire signed [`CalcTempBus]          temp_b2_7_25_i;
wire signed [`CalcTempBus]          temp_b2_7_26_r;
wire signed [`CalcTempBus]          temp_b2_7_26_i;
wire signed [`CalcTempBus]          temp_b2_7_27_r;
wire signed [`CalcTempBus]          temp_b2_7_27_i;
wire signed [`CalcTempBus]          temp_b2_7_28_r;
wire signed [`CalcTempBus]          temp_b2_7_28_i;
wire signed [`CalcTempBus]          temp_b2_7_29_r;
wire signed [`CalcTempBus]          temp_b2_7_29_i;
wire signed [`CalcTempBus]          temp_b2_7_30_r;
wire signed [`CalcTempBus]          temp_b2_7_30_i;
wire signed [`CalcTempBus]          temp_b2_7_31_r;
wire signed [`CalcTempBus]          temp_b2_7_31_i;
wire signed [`CalcTempBus]          temp_b2_7_32_r;
wire signed [`CalcTempBus]          temp_b2_7_32_i;
wire signed [`CalcTempBus]          temp_b2_8_1_r;
wire signed [`CalcTempBus]          temp_b2_8_1_i;
wire signed [`CalcTempBus]          temp_b2_8_2_r;
wire signed [`CalcTempBus]          temp_b2_8_2_i;
wire signed [`CalcTempBus]          temp_b2_8_3_r;
wire signed [`CalcTempBus]          temp_b2_8_3_i;
wire signed [`CalcTempBus]          temp_b2_8_4_r;
wire signed [`CalcTempBus]          temp_b2_8_4_i;
wire signed [`CalcTempBus]          temp_b2_8_5_r;
wire signed [`CalcTempBus]          temp_b2_8_5_i;
wire signed [`CalcTempBus]          temp_b2_8_6_r;
wire signed [`CalcTempBus]          temp_b2_8_6_i;
wire signed [`CalcTempBus]          temp_b2_8_7_r;
wire signed [`CalcTempBus]          temp_b2_8_7_i;
wire signed [`CalcTempBus]          temp_b2_8_8_r;
wire signed [`CalcTempBus]          temp_b2_8_8_i;
wire signed [`CalcTempBus]          temp_b2_8_9_r;
wire signed [`CalcTempBus]          temp_b2_8_9_i;
wire signed [`CalcTempBus]          temp_b2_8_10_r;
wire signed [`CalcTempBus]          temp_b2_8_10_i;
wire signed [`CalcTempBus]          temp_b2_8_11_r;
wire signed [`CalcTempBus]          temp_b2_8_11_i;
wire signed [`CalcTempBus]          temp_b2_8_12_r;
wire signed [`CalcTempBus]          temp_b2_8_12_i;
wire signed [`CalcTempBus]          temp_b2_8_13_r;
wire signed [`CalcTempBus]          temp_b2_8_13_i;
wire signed [`CalcTempBus]          temp_b2_8_14_r;
wire signed [`CalcTempBus]          temp_b2_8_14_i;
wire signed [`CalcTempBus]          temp_b2_8_15_r;
wire signed [`CalcTempBus]          temp_b2_8_15_i;
wire signed [`CalcTempBus]          temp_b2_8_16_r;
wire signed [`CalcTempBus]          temp_b2_8_16_i;
wire signed [`CalcTempBus]          temp_b2_8_17_r;
wire signed [`CalcTempBus]          temp_b2_8_17_i;
wire signed [`CalcTempBus]          temp_b2_8_18_r;
wire signed [`CalcTempBus]          temp_b2_8_18_i;
wire signed [`CalcTempBus]          temp_b2_8_19_r;
wire signed [`CalcTempBus]          temp_b2_8_19_i;
wire signed [`CalcTempBus]          temp_b2_8_20_r;
wire signed [`CalcTempBus]          temp_b2_8_20_i;
wire signed [`CalcTempBus]          temp_b2_8_21_r;
wire signed [`CalcTempBus]          temp_b2_8_21_i;
wire signed [`CalcTempBus]          temp_b2_8_22_r;
wire signed [`CalcTempBus]          temp_b2_8_22_i;
wire signed [`CalcTempBus]          temp_b2_8_23_r;
wire signed [`CalcTempBus]          temp_b2_8_23_i;
wire signed [`CalcTempBus]          temp_b2_8_24_r;
wire signed [`CalcTempBus]          temp_b2_8_24_i;
wire signed [`CalcTempBus]          temp_b2_8_25_r;
wire signed [`CalcTempBus]          temp_b2_8_25_i;
wire signed [`CalcTempBus]          temp_b2_8_26_r;
wire signed [`CalcTempBus]          temp_b2_8_26_i;
wire signed [`CalcTempBus]          temp_b2_8_27_r;
wire signed [`CalcTempBus]          temp_b2_8_27_i;
wire signed [`CalcTempBus]          temp_b2_8_28_r;
wire signed [`CalcTempBus]          temp_b2_8_28_i;
wire signed [`CalcTempBus]          temp_b2_8_29_r;
wire signed [`CalcTempBus]          temp_b2_8_29_i;
wire signed [`CalcTempBus]          temp_b2_8_30_r;
wire signed [`CalcTempBus]          temp_b2_8_30_i;
wire signed [`CalcTempBus]          temp_b2_8_31_r;
wire signed [`CalcTempBus]          temp_b2_8_31_i;
wire signed [`CalcTempBus]          temp_b2_8_32_r;
wire signed [`CalcTempBus]          temp_b2_8_32_i;
wire signed [`CalcTempBus]          temp_b2_9_1_r;
wire signed [`CalcTempBus]          temp_b2_9_1_i;
wire signed [`CalcTempBus]          temp_b2_9_2_r;
wire signed [`CalcTempBus]          temp_b2_9_2_i;
wire signed [`CalcTempBus]          temp_b2_9_3_r;
wire signed [`CalcTempBus]          temp_b2_9_3_i;
wire signed [`CalcTempBus]          temp_b2_9_4_r;
wire signed [`CalcTempBus]          temp_b2_9_4_i;
wire signed [`CalcTempBus]          temp_b2_9_5_r;
wire signed [`CalcTempBus]          temp_b2_9_5_i;
wire signed [`CalcTempBus]          temp_b2_9_6_r;
wire signed [`CalcTempBus]          temp_b2_9_6_i;
wire signed [`CalcTempBus]          temp_b2_9_7_r;
wire signed [`CalcTempBus]          temp_b2_9_7_i;
wire signed [`CalcTempBus]          temp_b2_9_8_r;
wire signed [`CalcTempBus]          temp_b2_9_8_i;
wire signed [`CalcTempBus]          temp_b2_9_9_r;
wire signed [`CalcTempBus]          temp_b2_9_9_i;
wire signed [`CalcTempBus]          temp_b2_9_10_r;
wire signed [`CalcTempBus]          temp_b2_9_10_i;
wire signed [`CalcTempBus]          temp_b2_9_11_r;
wire signed [`CalcTempBus]          temp_b2_9_11_i;
wire signed [`CalcTempBus]          temp_b2_9_12_r;
wire signed [`CalcTempBus]          temp_b2_9_12_i;
wire signed [`CalcTempBus]          temp_b2_9_13_r;
wire signed [`CalcTempBus]          temp_b2_9_13_i;
wire signed [`CalcTempBus]          temp_b2_9_14_r;
wire signed [`CalcTempBus]          temp_b2_9_14_i;
wire signed [`CalcTempBus]          temp_b2_9_15_r;
wire signed [`CalcTempBus]          temp_b2_9_15_i;
wire signed [`CalcTempBus]          temp_b2_9_16_r;
wire signed [`CalcTempBus]          temp_b2_9_16_i;
wire signed [`CalcTempBus]          temp_b2_9_17_r;
wire signed [`CalcTempBus]          temp_b2_9_17_i;
wire signed [`CalcTempBus]          temp_b2_9_18_r;
wire signed [`CalcTempBus]          temp_b2_9_18_i;
wire signed [`CalcTempBus]          temp_b2_9_19_r;
wire signed [`CalcTempBus]          temp_b2_9_19_i;
wire signed [`CalcTempBus]          temp_b2_9_20_r;
wire signed [`CalcTempBus]          temp_b2_9_20_i;
wire signed [`CalcTempBus]          temp_b2_9_21_r;
wire signed [`CalcTempBus]          temp_b2_9_21_i;
wire signed [`CalcTempBus]          temp_b2_9_22_r;
wire signed [`CalcTempBus]          temp_b2_9_22_i;
wire signed [`CalcTempBus]          temp_b2_9_23_r;
wire signed [`CalcTempBus]          temp_b2_9_23_i;
wire signed [`CalcTempBus]          temp_b2_9_24_r;
wire signed [`CalcTempBus]          temp_b2_9_24_i;
wire signed [`CalcTempBus]          temp_b2_9_25_r;
wire signed [`CalcTempBus]          temp_b2_9_25_i;
wire signed [`CalcTempBus]          temp_b2_9_26_r;
wire signed [`CalcTempBus]          temp_b2_9_26_i;
wire signed [`CalcTempBus]          temp_b2_9_27_r;
wire signed [`CalcTempBus]          temp_b2_9_27_i;
wire signed [`CalcTempBus]          temp_b2_9_28_r;
wire signed [`CalcTempBus]          temp_b2_9_28_i;
wire signed [`CalcTempBus]          temp_b2_9_29_r;
wire signed [`CalcTempBus]          temp_b2_9_29_i;
wire signed [`CalcTempBus]          temp_b2_9_30_r;
wire signed [`CalcTempBus]          temp_b2_9_30_i;
wire signed [`CalcTempBus]          temp_b2_9_31_r;
wire signed [`CalcTempBus]          temp_b2_9_31_i;
wire signed [`CalcTempBus]          temp_b2_9_32_r;
wire signed [`CalcTempBus]          temp_b2_9_32_i;
wire signed [`CalcTempBus]          temp_b2_10_1_r;
wire signed [`CalcTempBus]          temp_b2_10_1_i;
wire signed [`CalcTempBus]          temp_b2_10_2_r;
wire signed [`CalcTempBus]          temp_b2_10_2_i;
wire signed [`CalcTempBus]          temp_b2_10_3_r;
wire signed [`CalcTempBus]          temp_b2_10_3_i;
wire signed [`CalcTempBus]          temp_b2_10_4_r;
wire signed [`CalcTempBus]          temp_b2_10_4_i;
wire signed [`CalcTempBus]          temp_b2_10_5_r;
wire signed [`CalcTempBus]          temp_b2_10_5_i;
wire signed [`CalcTempBus]          temp_b2_10_6_r;
wire signed [`CalcTempBus]          temp_b2_10_6_i;
wire signed [`CalcTempBus]          temp_b2_10_7_r;
wire signed [`CalcTempBus]          temp_b2_10_7_i;
wire signed [`CalcTempBus]          temp_b2_10_8_r;
wire signed [`CalcTempBus]          temp_b2_10_8_i;
wire signed [`CalcTempBus]          temp_b2_10_9_r;
wire signed [`CalcTempBus]          temp_b2_10_9_i;
wire signed [`CalcTempBus]          temp_b2_10_10_r;
wire signed [`CalcTempBus]          temp_b2_10_10_i;
wire signed [`CalcTempBus]          temp_b2_10_11_r;
wire signed [`CalcTempBus]          temp_b2_10_11_i;
wire signed [`CalcTempBus]          temp_b2_10_12_r;
wire signed [`CalcTempBus]          temp_b2_10_12_i;
wire signed [`CalcTempBus]          temp_b2_10_13_r;
wire signed [`CalcTempBus]          temp_b2_10_13_i;
wire signed [`CalcTempBus]          temp_b2_10_14_r;
wire signed [`CalcTempBus]          temp_b2_10_14_i;
wire signed [`CalcTempBus]          temp_b2_10_15_r;
wire signed [`CalcTempBus]          temp_b2_10_15_i;
wire signed [`CalcTempBus]          temp_b2_10_16_r;
wire signed [`CalcTempBus]          temp_b2_10_16_i;
wire signed [`CalcTempBus]          temp_b2_10_17_r;
wire signed [`CalcTempBus]          temp_b2_10_17_i;
wire signed [`CalcTempBus]          temp_b2_10_18_r;
wire signed [`CalcTempBus]          temp_b2_10_18_i;
wire signed [`CalcTempBus]          temp_b2_10_19_r;
wire signed [`CalcTempBus]          temp_b2_10_19_i;
wire signed [`CalcTempBus]          temp_b2_10_20_r;
wire signed [`CalcTempBus]          temp_b2_10_20_i;
wire signed [`CalcTempBus]          temp_b2_10_21_r;
wire signed [`CalcTempBus]          temp_b2_10_21_i;
wire signed [`CalcTempBus]          temp_b2_10_22_r;
wire signed [`CalcTempBus]          temp_b2_10_22_i;
wire signed [`CalcTempBus]          temp_b2_10_23_r;
wire signed [`CalcTempBus]          temp_b2_10_23_i;
wire signed [`CalcTempBus]          temp_b2_10_24_r;
wire signed [`CalcTempBus]          temp_b2_10_24_i;
wire signed [`CalcTempBus]          temp_b2_10_25_r;
wire signed [`CalcTempBus]          temp_b2_10_25_i;
wire signed [`CalcTempBus]          temp_b2_10_26_r;
wire signed [`CalcTempBus]          temp_b2_10_26_i;
wire signed [`CalcTempBus]          temp_b2_10_27_r;
wire signed [`CalcTempBus]          temp_b2_10_27_i;
wire signed [`CalcTempBus]          temp_b2_10_28_r;
wire signed [`CalcTempBus]          temp_b2_10_28_i;
wire signed [`CalcTempBus]          temp_b2_10_29_r;
wire signed [`CalcTempBus]          temp_b2_10_29_i;
wire signed [`CalcTempBus]          temp_b2_10_30_r;
wire signed [`CalcTempBus]          temp_b2_10_30_i;
wire signed [`CalcTempBus]          temp_b2_10_31_r;
wire signed [`CalcTempBus]          temp_b2_10_31_i;
wire signed [`CalcTempBus]          temp_b2_10_32_r;
wire signed [`CalcTempBus]          temp_b2_10_32_i;
wire signed [`CalcTempBus]          temp_b2_11_1_r;
wire signed [`CalcTempBus]          temp_b2_11_1_i;
wire signed [`CalcTempBus]          temp_b2_11_2_r;
wire signed [`CalcTempBus]          temp_b2_11_2_i;
wire signed [`CalcTempBus]          temp_b2_11_3_r;
wire signed [`CalcTempBus]          temp_b2_11_3_i;
wire signed [`CalcTempBus]          temp_b2_11_4_r;
wire signed [`CalcTempBus]          temp_b2_11_4_i;
wire signed [`CalcTempBus]          temp_b2_11_5_r;
wire signed [`CalcTempBus]          temp_b2_11_5_i;
wire signed [`CalcTempBus]          temp_b2_11_6_r;
wire signed [`CalcTempBus]          temp_b2_11_6_i;
wire signed [`CalcTempBus]          temp_b2_11_7_r;
wire signed [`CalcTempBus]          temp_b2_11_7_i;
wire signed [`CalcTempBus]          temp_b2_11_8_r;
wire signed [`CalcTempBus]          temp_b2_11_8_i;
wire signed [`CalcTempBus]          temp_b2_11_9_r;
wire signed [`CalcTempBus]          temp_b2_11_9_i;
wire signed [`CalcTempBus]          temp_b2_11_10_r;
wire signed [`CalcTempBus]          temp_b2_11_10_i;
wire signed [`CalcTempBus]          temp_b2_11_11_r;
wire signed [`CalcTempBus]          temp_b2_11_11_i;
wire signed [`CalcTempBus]          temp_b2_11_12_r;
wire signed [`CalcTempBus]          temp_b2_11_12_i;
wire signed [`CalcTempBus]          temp_b2_11_13_r;
wire signed [`CalcTempBus]          temp_b2_11_13_i;
wire signed [`CalcTempBus]          temp_b2_11_14_r;
wire signed [`CalcTempBus]          temp_b2_11_14_i;
wire signed [`CalcTempBus]          temp_b2_11_15_r;
wire signed [`CalcTempBus]          temp_b2_11_15_i;
wire signed [`CalcTempBus]          temp_b2_11_16_r;
wire signed [`CalcTempBus]          temp_b2_11_16_i;
wire signed [`CalcTempBus]          temp_b2_11_17_r;
wire signed [`CalcTempBus]          temp_b2_11_17_i;
wire signed [`CalcTempBus]          temp_b2_11_18_r;
wire signed [`CalcTempBus]          temp_b2_11_18_i;
wire signed [`CalcTempBus]          temp_b2_11_19_r;
wire signed [`CalcTempBus]          temp_b2_11_19_i;
wire signed [`CalcTempBus]          temp_b2_11_20_r;
wire signed [`CalcTempBus]          temp_b2_11_20_i;
wire signed [`CalcTempBus]          temp_b2_11_21_r;
wire signed [`CalcTempBus]          temp_b2_11_21_i;
wire signed [`CalcTempBus]          temp_b2_11_22_r;
wire signed [`CalcTempBus]          temp_b2_11_22_i;
wire signed [`CalcTempBus]          temp_b2_11_23_r;
wire signed [`CalcTempBus]          temp_b2_11_23_i;
wire signed [`CalcTempBus]          temp_b2_11_24_r;
wire signed [`CalcTempBus]          temp_b2_11_24_i;
wire signed [`CalcTempBus]          temp_b2_11_25_r;
wire signed [`CalcTempBus]          temp_b2_11_25_i;
wire signed [`CalcTempBus]          temp_b2_11_26_r;
wire signed [`CalcTempBus]          temp_b2_11_26_i;
wire signed [`CalcTempBus]          temp_b2_11_27_r;
wire signed [`CalcTempBus]          temp_b2_11_27_i;
wire signed [`CalcTempBus]          temp_b2_11_28_r;
wire signed [`CalcTempBus]          temp_b2_11_28_i;
wire signed [`CalcTempBus]          temp_b2_11_29_r;
wire signed [`CalcTempBus]          temp_b2_11_29_i;
wire signed [`CalcTempBus]          temp_b2_11_30_r;
wire signed [`CalcTempBus]          temp_b2_11_30_i;
wire signed [`CalcTempBus]          temp_b2_11_31_r;
wire signed [`CalcTempBus]          temp_b2_11_31_i;
wire signed [`CalcTempBus]          temp_b2_11_32_r;
wire signed [`CalcTempBus]          temp_b2_11_32_i;
wire signed [`CalcTempBus]          temp_b2_12_1_r;
wire signed [`CalcTempBus]          temp_b2_12_1_i;
wire signed [`CalcTempBus]          temp_b2_12_2_r;
wire signed [`CalcTempBus]          temp_b2_12_2_i;
wire signed [`CalcTempBus]          temp_b2_12_3_r;
wire signed [`CalcTempBus]          temp_b2_12_3_i;
wire signed [`CalcTempBus]          temp_b2_12_4_r;
wire signed [`CalcTempBus]          temp_b2_12_4_i;
wire signed [`CalcTempBus]          temp_b2_12_5_r;
wire signed [`CalcTempBus]          temp_b2_12_5_i;
wire signed [`CalcTempBus]          temp_b2_12_6_r;
wire signed [`CalcTempBus]          temp_b2_12_6_i;
wire signed [`CalcTempBus]          temp_b2_12_7_r;
wire signed [`CalcTempBus]          temp_b2_12_7_i;
wire signed [`CalcTempBus]          temp_b2_12_8_r;
wire signed [`CalcTempBus]          temp_b2_12_8_i;
wire signed [`CalcTempBus]          temp_b2_12_9_r;
wire signed [`CalcTempBus]          temp_b2_12_9_i;
wire signed [`CalcTempBus]          temp_b2_12_10_r;
wire signed [`CalcTempBus]          temp_b2_12_10_i;
wire signed [`CalcTempBus]          temp_b2_12_11_r;
wire signed [`CalcTempBus]          temp_b2_12_11_i;
wire signed [`CalcTempBus]          temp_b2_12_12_r;
wire signed [`CalcTempBus]          temp_b2_12_12_i;
wire signed [`CalcTempBus]          temp_b2_12_13_r;
wire signed [`CalcTempBus]          temp_b2_12_13_i;
wire signed [`CalcTempBus]          temp_b2_12_14_r;
wire signed [`CalcTempBus]          temp_b2_12_14_i;
wire signed [`CalcTempBus]          temp_b2_12_15_r;
wire signed [`CalcTempBus]          temp_b2_12_15_i;
wire signed [`CalcTempBus]          temp_b2_12_16_r;
wire signed [`CalcTempBus]          temp_b2_12_16_i;
wire signed [`CalcTempBus]          temp_b2_12_17_r;
wire signed [`CalcTempBus]          temp_b2_12_17_i;
wire signed [`CalcTempBus]          temp_b2_12_18_r;
wire signed [`CalcTempBus]          temp_b2_12_18_i;
wire signed [`CalcTempBus]          temp_b2_12_19_r;
wire signed [`CalcTempBus]          temp_b2_12_19_i;
wire signed [`CalcTempBus]          temp_b2_12_20_r;
wire signed [`CalcTempBus]          temp_b2_12_20_i;
wire signed [`CalcTempBus]          temp_b2_12_21_r;
wire signed [`CalcTempBus]          temp_b2_12_21_i;
wire signed [`CalcTempBus]          temp_b2_12_22_r;
wire signed [`CalcTempBus]          temp_b2_12_22_i;
wire signed [`CalcTempBus]          temp_b2_12_23_r;
wire signed [`CalcTempBus]          temp_b2_12_23_i;
wire signed [`CalcTempBus]          temp_b2_12_24_r;
wire signed [`CalcTempBus]          temp_b2_12_24_i;
wire signed [`CalcTempBus]          temp_b2_12_25_r;
wire signed [`CalcTempBus]          temp_b2_12_25_i;
wire signed [`CalcTempBus]          temp_b2_12_26_r;
wire signed [`CalcTempBus]          temp_b2_12_26_i;
wire signed [`CalcTempBus]          temp_b2_12_27_r;
wire signed [`CalcTempBus]          temp_b2_12_27_i;
wire signed [`CalcTempBus]          temp_b2_12_28_r;
wire signed [`CalcTempBus]          temp_b2_12_28_i;
wire signed [`CalcTempBus]          temp_b2_12_29_r;
wire signed [`CalcTempBus]          temp_b2_12_29_i;
wire signed [`CalcTempBus]          temp_b2_12_30_r;
wire signed [`CalcTempBus]          temp_b2_12_30_i;
wire signed [`CalcTempBus]          temp_b2_12_31_r;
wire signed [`CalcTempBus]          temp_b2_12_31_i;
wire signed [`CalcTempBus]          temp_b2_12_32_r;
wire signed [`CalcTempBus]          temp_b2_12_32_i;
wire signed [`CalcTempBus]          temp_b2_13_1_r;
wire signed [`CalcTempBus]          temp_b2_13_1_i;
wire signed [`CalcTempBus]          temp_b2_13_2_r;
wire signed [`CalcTempBus]          temp_b2_13_2_i;
wire signed [`CalcTempBus]          temp_b2_13_3_r;
wire signed [`CalcTempBus]          temp_b2_13_3_i;
wire signed [`CalcTempBus]          temp_b2_13_4_r;
wire signed [`CalcTempBus]          temp_b2_13_4_i;
wire signed [`CalcTempBus]          temp_b2_13_5_r;
wire signed [`CalcTempBus]          temp_b2_13_5_i;
wire signed [`CalcTempBus]          temp_b2_13_6_r;
wire signed [`CalcTempBus]          temp_b2_13_6_i;
wire signed [`CalcTempBus]          temp_b2_13_7_r;
wire signed [`CalcTempBus]          temp_b2_13_7_i;
wire signed [`CalcTempBus]          temp_b2_13_8_r;
wire signed [`CalcTempBus]          temp_b2_13_8_i;
wire signed [`CalcTempBus]          temp_b2_13_9_r;
wire signed [`CalcTempBus]          temp_b2_13_9_i;
wire signed [`CalcTempBus]          temp_b2_13_10_r;
wire signed [`CalcTempBus]          temp_b2_13_10_i;
wire signed [`CalcTempBus]          temp_b2_13_11_r;
wire signed [`CalcTempBus]          temp_b2_13_11_i;
wire signed [`CalcTempBus]          temp_b2_13_12_r;
wire signed [`CalcTempBus]          temp_b2_13_12_i;
wire signed [`CalcTempBus]          temp_b2_13_13_r;
wire signed [`CalcTempBus]          temp_b2_13_13_i;
wire signed [`CalcTempBus]          temp_b2_13_14_r;
wire signed [`CalcTempBus]          temp_b2_13_14_i;
wire signed [`CalcTempBus]          temp_b2_13_15_r;
wire signed [`CalcTempBus]          temp_b2_13_15_i;
wire signed [`CalcTempBus]          temp_b2_13_16_r;
wire signed [`CalcTempBus]          temp_b2_13_16_i;
wire signed [`CalcTempBus]          temp_b2_13_17_r;
wire signed [`CalcTempBus]          temp_b2_13_17_i;
wire signed [`CalcTempBus]          temp_b2_13_18_r;
wire signed [`CalcTempBus]          temp_b2_13_18_i;
wire signed [`CalcTempBus]          temp_b2_13_19_r;
wire signed [`CalcTempBus]          temp_b2_13_19_i;
wire signed [`CalcTempBus]          temp_b2_13_20_r;
wire signed [`CalcTempBus]          temp_b2_13_20_i;
wire signed [`CalcTempBus]          temp_b2_13_21_r;
wire signed [`CalcTempBus]          temp_b2_13_21_i;
wire signed [`CalcTempBus]          temp_b2_13_22_r;
wire signed [`CalcTempBus]          temp_b2_13_22_i;
wire signed [`CalcTempBus]          temp_b2_13_23_r;
wire signed [`CalcTempBus]          temp_b2_13_23_i;
wire signed [`CalcTempBus]          temp_b2_13_24_r;
wire signed [`CalcTempBus]          temp_b2_13_24_i;
wire signed [`CalcTempBus]          temp_b2_13_25_r;
wire signed [`CalcTempBus]          temp_b2_13_25_i;
wire signed [`CalcTempBus]          temp_b2_13_26_r;
wire signed [`CalcTempBus]          temp_b2_13_26_i;
wire signed [`CalcTempBus]          temp_b2_13_27_r;
wire signed [`CalcTempBus]          temp_b2_13_27_i;
wire signed [`CalcTempBus]          temp_b2_13_28_r;
wire signed [`CalcTempBus]          temp_b2_13_28_i;
wire signed [`CalcTempBus]          temp_b2_13_29_r;
wire signed [`CalcTempBus]          temp_b2_13_29_i;
wire signed [`CalcTempBus]          temp_b2_13_30_r;
wire signed [`CalcTempBus]          temp_b2_13_30_i;
wire signed [`CalcTempBus]          temp_b2_13_31_r;
wire signed [`CalcTempBus]          temp_b2_13_31_i;
wire signed [`CalcTempBus]          temp_b2_13_32_r;
wire signed [`CalcTempBus]          temp_b2_13_32_i;
wire signed [`CalcTempBus]          temp_b2_14_1_r;
wire signed [`CalcTempBus]          temp_b2_14_1_i;
wire signed [`CalcTempBus]          temp_b2_14_2_r;
wire signed [`CalcTempBus]          temp_b2_14_2_i;
wire signed [`CalcTempBus]          temp_b2_14_3_r;
wire signed [`CalcTempBus]          temp_b2_14_3_i;
wire signed [`CalcTempBus]          temp_b2_14_4_r;
wire signed [`CalcTempBus]          temp_b2_14_4_i;
wire signed [`CalcTempBus]          temp_b2_14_5_r;
wire signed [`CalcTempBus]          temp_b2_14_5_i;
wire signed [`CalcTempBus]          temp_b2_14_6_r;
wire signed [`CalcTempBus]          temp_b2_14_6_i;
wire signed [`CalcTempBus]          temp_b2_14_7_r;
wire signed [`CalcTempBus]          temp_b2_14_7_i;
wire signed [`CalcTempBus]          temp_b2_14_8_r;
wire signed [`CalcTempBus]          temp_b2_14_8_i;
wire signed [`CalcTempBus]          temp_b2_14_9_r;
wire signed [`CalcTempBus]          temp_b2_14_9_i;
wire signed [`CalcTempBus]          temp_b2_14_10_r;
wire signed [`CalcTempBus]          temp_b2_14_10_i;
wire signed [`CalcTempBus]          temp_b2_14_11_r;
wire signed [`CalcTempBus]          temp_b2_14_11_i;
wire signed [`CalcTempBus]          temp_b2_14_12_r;
wire signed [`CalcTempBus]          temp_b2_14_12_i;
wire signed [`CalcTempBus]          temp_b2_14_13_r;
wire signed [`CalcTempBus]          temp_b2_14_13_i;
wire signed [`CalcTempBus]          temp_b2_14_14_r;
wire signed [`CalcTempBus]          temp_b2_14_14_i;
wire signed [`CalcTempBus]          temp_b2_14_15_r;
wire signed [`CalcTempBus]          temp_b2_14_15_i;
wire signed [`CalcTempBus]          temp_b2_14_16_r;
wire signed [`CalcTempBus]          temp_b2_14_16_i;
wire signed [`CalcTempBus]          temp_b2_14_17_r;
wire signed [`CalcTempBus]          temp_b2_14_17_i;
wire signed [`CalcTempBus]          temp_b2_14_18_r;
wire signed [`CalcTempBus]          temp_b2_14_18_i;
wire signed [`CalcTempBus]          temp_b2_14_19_r;
wire signed [`CalcTempBus]          temp_b2_14_19_i;
wire signed [`CalcTempBus]          temp_b2_14_20_r;
wire signed [`CalcTempBus]          temp_b2_14_20_i;
wire signed [`CalcTempBus]          temp_b2_14_21_r;
wire signed [`CalcTempBus]          temp_b2_14_21_i;
wire signed [`CalcTempBus]          temp_b2_14_22_r;
wire signed [`CalcTempBus]          temp_b2_14_22_i;
wire signed [`CalcTempBus]          temp_b2_14_23_r;
wire signed [`CalcTempBus]          temp_b2_14_23_i;
wire signed [`CalcTempBus]          temp_b2_14_24_r;
wire signed [`CalcTempBus]          temp_b2_14_24_i;
wire signed [`CalcTempBus]          temp_b2_14_25_r;
wire signed [`CalcTempBus]          temp_b2_14_25_i;
wire signed [`CalcTempBus]          temp_b2_14_26_r;
wire signed [`CalcTempBus]          temp_b2_14_26_i;
wire signed [`CalcTempBus]          temp_b2_14_27_r;
wire signed [`CalcTempBus]          temp_b2_14_27_i;
wire signed [`CalcTempBus]          temp_b2_14_28_r;
wire signed [`CalcTempBus]          temp_b2_14_28_i;
wire signed [`CalcTempBus]          temp_b2_14_29_r;
wire signed [`CalcTempBus]          temp_b2_14_29_i;
wire signed [`CalcTempBus]          temp_b2_14_30_r;
wire signed [`CalcTempBus]          temp_b2_14_30_i;
wire signed [`CalcTempBus]          temp_b2_14_31_r;
wire signed [`CalcTempBus]          temp_b2_14_31_i;
wire signed [`CalcTempBus]          temp_b2_14_32_r;
wire signed [`CalcTempBus]          temp_b2_14_32_i;
wire signed [`CalcTempBus]          temp_b2_15_1_r;
wire signed [`CalcTempBus]          temp_b2_15_1_i;
wire signed [`CalcTempBus]          temp_b2_15_2_r;
wire signed [`CalcTempBus]          temp_b2_15_2_i;
wire signed [`CalcTempBus]          temp_b2_15_3_r;
wire signed [`CalcTempBus]          temp_b2_15_3_i;
wire signed [`CalcTempBus]          temp_b2_15_4_r;
wire signed [`CalcTempBus]          temp_b2_15_4_i;
wire signed [`CalcTempBus]          temp_b2_15_5_r;
wire signed [`CalcTempBus]          temp_b2_15_5_i;
wire signed [`CalcTempBus]          temp_b2_15_6_r;
wire signed [`CalcTempBus]          temp_b2_15_6_i;
wire signed [`CalcTempBus]          temp_b2_15_7_r;
wire signed [`CalcTempBus]          temp_b2_15_7_i;
wire signed [`CalcTempBus]          temp_b2_15_8_r;
wire signed [`CalcTempBus]          temp_b2_15_8_i;
wire signed [`CalcTempBus]          temp_b2_15_9_r;
wire signed [`CalcTempBus]          temp_b2_15_9_i;
wire signed [`CalcTempBus]          temp_b2_15_10_r;
wire signed [`CalcTempBus]          temp_b2_15_10_i;
wire signed [`CalcTempBus]          temp_b2_15_11_r;
wire signed [`CalcTempBus]          temp_b2_15_11_i;
wire signed [`CalcTempBus]          temp_b2_15_12_r;
wire signed [`CalcTempBus]          temp_b2_15_12_i;
wire signed [`CalcTempBus]          temp_b2_15_13_r;
wire signed [`CalcTempBus]          temp_b2_15_13_i;
wire signed [`CalcTempBus]          temp_b2_15_14_r;
wire signed [`CalcTempBus]          temp_b2_15_14_i;
wire signed [`CalcTempBus]          temp_b2_15_15_r;
wire signed [`CalcTempBus]          temp_b2_15_15_i;
wire signed [`CalcTempBus]          temp_b2_15_16_r;
wire signed [`CalcTempBus]          temp_b2_15_16_i;
wire signed [`CalcTempBus]          temp_b2_15_17_r;
wire signed [`CalcTempBus]          temp_b2_15_17_i;
wire signed [`CalcTempBus]          temp_b2_15_18_r;
wire signed [`CalcTempBus]          temp_b2_15_18_i;
wire signed [`CalcTempBus]          temp_b2_15_19_r;
wire signed [`CalcTempBus]          temp_b2_15_19_i;
wire signed [`CalcTempBus]          temp_b2_15_20_r;
wire signed [`CalcTempBus]          temp_b2_15_20_i;
wire signed [`CalcTempBus]          temp_b2_15_21_r;
wire signed [`CalcTempBus]          temp_b2_15_21_i;
wire signed [`CalcTempBus]          temp_b2_15_22_r;
wire signed [`CalcTempBus]          temp_b2_15_22_i;
wire signed [`CalcTempBus]          temp_b2_15_23_r;
wire signed [`CalcTempBus]          temp_b2_15_23_i;
wire signed [`CalcTempBus]          temp_b2_15_24_r;
wire signed [`CalcTempBus]          temp_b2_15_24_i;
wire signed [`CalcTempBus]          temp_b2_15_25_r;
wire signed [`CalcTempBus]          temp_b2_15_25_i;
wire signed [`CalcTempBus]          temp_b2_15_26_r;
wire signed [`CalcTempBus]          temp_b2_15_26_i;
wire signed [`CalcTempBus]          temp_b2_15_27_r;
wire signed [`CalcTempBus]          temp_b2_15_27_i;
wire signed [`CalcTempBus]          temp_b2_15_28_r;
wire signed [`CalcTempBus]          temp_b2_15_28_i;
wire signed [`CalcTempBus]          temp_b2_15_29_r;
wire signed [`CalcTempBus]          temp_b2_15_29_i;
wire signed [`CalcTempBus]          temp_b2_15_30_r;
wire signed [`CalcTempBus]          temp_b2_15_30_i;
wire signed [`CalcTempBus]          temp_b2_15_31_r;
wire signed [`CalcTempBus]          temp_b2_15_31_i;
wire signed [`CalcTempBus]          temp_b2_15_32_r;
wire signed [`CalcTempBus]          temp_b2_15_32_i;
wire signed [`CalcTempBus]          temp_b2_16_1_r;
wire signed [`CalcTempBus]          temp_b2_16_1_i;
wire signed [`CalcTempBus]          temp_b2_16_2_r;
wire signed [`CalcTempBus]          temp_b2_16_2_i;
wire signed [`CalcTempBus]          temp_b2_16_3_r;
wire signed [`CalcTempBus]          temp_b2_16_3_i;
wire signed [`CalcTempBus]          temp_b2_16_4_r;
wire signed [`CalcTempBus]          temp_b2_16_4_i;
wire signed [`CalcTempBus]          temp_b2_16_5_r;
wire signed [`CalcTempBus]          temp_b2_16_5_i;
wire signed [`CalcTempBus]          temp_b2_16_6_r;
wire signed [`CalcTempBus]          temp_b2_16_6_i;
wire signed [`CalcTempBus]          temp_b2_16_7_r;
wire signed [`CalcTempBus]          temp_b2_16_7_i;
wire signed [`CalcTempBus]          temp_b2_16_8_r;
wire signed [`CalcTempBus]          temp_b2_16_8_i;
wire signed [`CalcTempBus]          temp_b2_16_9_r;
wire signed [`CalcTempBus]          temp_b2_16_9_i;
wire signed [`CalcTempBus]          temp_b2_16_10_r;
wire signed [`CalcTempBus]          temp_b2_16_10_i;
wire signed [`CalcTempBus]          temp_b2_16_11_r;
wire signed [`CalcTempBus]          temp_b2_16_11_i;
wire signed [`CalcTempBus]          temp_b2_16_12_r;
wire signed [`CalcTempBus]          temp_b2_16_12_i;
wire signed [`CalcTempBus]          temp_b2_16_13_r;
wire signed [`CalcTempBus]          temp_b2_16_13_i;
wire signed [`CalcTempBus]          temp_b2_16_14_r;
wire signed [`CalcTempBus]          temp_b2_16_14_i;
wire signed [`CalcTempBus]          temp_b2_16_15_r;
wire signed [`CalcTempBus]          temp_b2_16_15_i;
wire signed [`CalcTempBus]          temp_b2_16_16_r;
wire signed [`CalcTempBus]          temp_b2_16_16_i;
wire signed [`CalcTempBus]          temp_b2_16_17_r;
wire signed [`CalcTempBus]          temp_b2_16_17_i;
wire signed [`CalcTempBus]          temp_b2_16_18_r;
wire signed [`CalcTempBus]          temp_b2_16_18_i;
wire signed [`CalcTempBus]          temp_b2_16_19_r;
wire signed [`CalcTempBus]          temp_b2_16_19_i;
wire signed [`CalcTempBus]          temp_b2_16_20_r;
wire signed [`CalcTempBus]          temp_b2_16_20_i;
wire signed [`CalcTempBus]          temp_b2_16_21_r;
wire signed [`CalcTempBus]          temp_b2_16_21_i;
wire signed [`CalcTempBus]          temp_b2_16_22_r;
wire signed [`CalcTempBus]          temp_b2_16_22_i;
wire signed [`CalcTempBus]          temp_b2_16_23_r;
wire signed [`CalcTempBus]          temp_b2_16_23_i;
wire signed [`CalcTempBus]          temp_b2_16_24_r;
wire signed [`CalcTempBus]          temp_b2_16_24_i;
wire signed [`CalcTempBus]          temp_b2_16_25_r;
wire signed [`CalcTempBus]          temp_b2_16_25_i;
wire signed [`CalcTempBus]          temp_b2_16_26_r;
wire signed [`CalcTempBus]          temp_b2_16_26_i;
wire signed [`CalcTempBus]          temp_b2_16_27_r;
wire signed [`CalcTempBus]          temp_b2_16_27_i;
wire signed [`CalcTempBus]          temp_b2_16_28_r;
wire signed [`CalcTempBus]          temp_b2_16_28_i;
wire signed [`CalcTempBus]          temp_b2_16_29_r;
wire signed [`CalcTempBus]          temp_b2_16_29_i;
wire signed [`CalcTempBus]          temp_b2_16_30_r;
wire signed [`CalcTempBus]          temp_b2_16_30_i;
wire signed [`CalcTempBus]          temp_b2_16_31_r;
wire signed [`CalcTempBus]          temp_b2_16_31_i;
wire signed [`CalcTempBus]          temp_b2_16_32_r;
wire signed [`CalcTempBus]          temp_b2_16_32_i;
wire signed [`CalcTempBus]          temp_b2_17_1_r;
wire signed [`CalcTempBus]          temp_b2_17_1_i;
wire signed [`CalcTempBus]          temp_b2_17_2_r;
wire signed [`CalcTempBus]          temp_b2_17_2_i;
wire signed [`CalcTempBus]          temp_b2_17_3_r;
wire signed [`CalcTempBus]          temp_b2_17_3_i;
wire signed [`CalcTempBus]          temp_b2_17_4_r;
wire signed [`CalcTempBus]          temp_b2_17_4_i;
wire signed [`CalcTempBus]          temp_b2_17_5_r;
wire signed [`CalcTempBus]          temp_b2_17_5_i;
wire signed [`CalcTempBus]          temp_b2_17_6_r;
wire signed [`CalcTempBus]          temp_b2_17_6_i;
wire signed [`CalcTempBus]          temp_b2_17_7_r;
wire signed [`CalcTempBus]          temp_b2_17_7_i;
wire signed [`CalcTempBus]          temp_b2_17_8_r;
wire signed [`CalcTempBus]          temp_b2_17_8_i;
wire signed [`CalcTempBus]          temp_b2_17_9_r;
wire signed [`CalcTempBus]          temp_b2_17_9_i;
wire signed [`CalcTempBus]          temp_b2_17_10_r;
wire signed [`CalcTempBus]          temp_b2_17_10_i;
wire signed [`CalcTempBus]          temp_b2_17_11_r;
wire signed [`CalcTempBus]          temp_b2_17_11_i;
wire signed [`CalcTempBus]          temp_b2_17_12_r;
wire signed [`CalcTempBus]          temp_b2_17_12_i;
wire signed [`CalcTempBus]          temp_b2_17_13_r;
wire signed [`CalcTempBus]          temp_b2_17_13_i;
wire signed [`CalcTempBus]          temp_b2_17_14_r;
wire signed [`CalcTempBus]          temp_b2_17_14_i;
wire signed [`CalcTempBus]          temp_b2_17_15_r;
wire signed [`CalcTempBus]          temp_b2_17_15_i;
wire signed [`CalcTempBus]          temp_b2_17_16_r;
wire signed [`CalcTempBus]          temp_b2_17_16_i;
wire signed [`CalcTempBus]          temp_b2_17_17_r;
wire signed [`CalcTempBus]          temp_b2_17_17_i;
wire signed [`CalcTempBus]          temp_b2_17_18_r;
wire signed [`CalcTempBus]          temp_b2_17_18_i;
wire signed [`CalcTempBus]          temp_b2_17_19_r;
wire signed [`CalcTempBus]          temp_b2_17_19_i;
wire signed [`CalcTempBus]          temp_b2_17_20_r;
wire signed [`CalcTempBus]          temp_b2_17_20_i;
wire signed [`CalcTempBus]          temp_b2_17_21_r;
wire signed [`CalcTempBus]          temp_b2_17_21_i;
wire signed [`CalcTempBus]          temp_b2_17_22_r;
wire signed [`CalcTempBus]          temp_b2_17_22_i;
wire signed [`CalcTempBus]          temp_b2_17_23_r;
wire signed [`CalcTempBus]          temp_b2_17_23_i;
wire signed [`CalcTempBus]          temp_b2_17_24_r;
wire signed [`CalcTempBus]          temp_b2_17_24_i;
wire signed [`CalcTempBus]          temp_b2_17_25_r;
wire signed [`CalcTempBus]          temp_b2_17_25_i;
wire signed [`CalcTempBus]          temp_b2_17_26_r;
wire signed [`CalcTempBus]          temp_b2_17_26_i;
wire signed [`CalcTempBus]          temp_b2_17_27_r;
wire signed [`CalcTempBus]          temp_b2_17_27_i;
wire signed [`CalcTempBus]          temp_b2_17_28_r;
wire signed [`CalcTempBus]          temp_b2_17_28_i;
wire signed [`CalcTempBus]          temp_b2_17_29_r;
wire signed [`CalcTempBus]          temp_b2_17_29_i;
wire signed [`CalcTempBus]          temp_b2_17_30_r;
wire signed [`CalcTempBus]          temp_b2_17_30_i;
wire signed [`CalcTempBus]          temp_b2_17_31_r;
wire signed [`CalcTempBus]          temp_b2_17_31_i;
wire signed [`CalcTempBus]          temp_b2_17_32_r;
wire signed [`CalcTempBus]          temp_b2_17_32_i;
wire signed [`CalcTempBus]          temp_b2_18_1_r;
wire signed [`CalcTempBus]          temp_b2_18_1_i;
wire signed [`CalcTempBus]          temp_b2_18_2_r;
wire signed [`CalcTempBus]          temp_b2_18_2_i;
wire signed [`CalcTempBus]          temp_b2_18_3_r;
wire signed [`CalcTempBus]          temp_b2_18_3_i;
wire signed [`CalcTempBus]          temp_b2_18_4_r;
wire signed [`CalcTempBus]          temp_b2_18_4_i;
wire signed [`CalcTempBus]          temp_b2_18_5_r;
wire signed [`CalcTempBus]          temp_b2_18_5_i;
wire signed [`CalcTempBus]          temp_b2_18_6_r;
wire signed [`CalcTempBus]          temp_b2_18_6_i;
wire signed [`CalcTempBus]          temp_b2_18_7_r;
wire signed [`CalcTempBus]          temp_b2_18_7_i;
wire signed [`CalcTempBus]          temp_b2_18_8_r;
wire signed [`CalcTempBus]          temp_b2_18_8_i;
wire signed [`CalcTempBus]          temp_b2_18_9_r;
wire signed [`CalcTempBus]          temp_b2_18_9_i;
wire signed [`CalcTempBus]          temp_b2_18_10_r;
wire signed [`CalcTempBus]          temp_b2_18_10_i;
wire signed [`CalcTempBus]          temp_b2_18_11_r;
wire signed [`CalcTempBus]          temp_b2_18_11_i;
wire signed [`CalcTempBus]          temp_b2_18_12_r;
wire signed [`CalcTempBus]          temp_b2_18_12_i;
wire signed [`CalcTempBus]          temp_b2_18_13_r;
wire signed [`CalcTempBus]          temp_b2_18_13_i;
wire signed [`CalcTempBus]          temp_b2_18_14_r;
wire signed [`CalcTempBus]          temp_b2_18_14_i;
wire signed [`CalcTempBus]          temp_b2_18_15_r;
wire signed [`CalcTempBus]          temp_b2_18_15_i;
wire signed [`CalcTempBus]          temp_b2_18_16_r;
wire signed [`CalcTempBus]          temp_b2_18_16_i;
wire signed [`CalcTempBus]          temp_b2_18_17_r;
wire signed [`CalcTempBus]          temp_b2_18_17_i;
wire signed [`CalcTempBus]          temp_b2_18_18_r;
wire signed [`CalcTempBus]          temp_b2_18_18_i;
wire signed [`CalcTempBus]          temp_b2_18_19_r;
wire signed [`CalcTempBus]          temp_b2_18_19_i;
wire signed [`CalcTempBus]          temp_b2_18_20_r;
wire signed [`CalcTempBus]          temp_b2_18_20_i;
wire signed [`CalcTempBus]          temp_b2_18_21_r;
wire signed [`CalcTempBus]          temp_b2_18_21_i;
wire signed [`CalcTempBus]          temp_b2_18_22_r;
wire signed [`CalcTempBus]          temp_b2_18_22_i;
wire signed [`CalcTempBus]          temp_b2_18_23_r;
wire signed [`CalcTempBus]          temp_b2_18_23_i;
wire signed [`CalcTempBus]          temp_b2_18_24_r;
wire signed [`CalcTempBus]          temp_b2_18_24_i;
wire signed [`CalcTempBus]          temp_b2_18_25_r;
wire signed [`CalcTempBus]          temp_b2_18_25_i;
wire signed [`CalcTempBus]          temp_b2_18_26_r;
wire signed [`CalcTempBus]          temp_b2_18_26_i;
wire signed [`CalcTempBus]          temp_b2_18_27_r;
wire signed [`CalcTempBus]          temp_b2_18_27_i;
wire signed [`CalcTempBus]          temp_b2_18_28_r;
wire signed [`CalcTempBus]          temp_b2_18_28_i;
wire signed [`CalcTempBus]          temp_b2_18_29_r;
wire signed [`CalcTempBus]          temp_b2_18_29_i;
wire signed [`CalcTempBus]          temp_b2_18_30_r;
wire signed [`CalcTempBus]          temp_b2_18_30_i;
wire signed [`CalcTempBus]          temp_b2_18_31_r;
wire signed [`CalcTempBus]          temp_b2_18_31_i;
wire signed [`CalcTempBus]          temp_b2_18_32_r;
wire signed [`CalcTempBus]          temp_b2_18_32_i;
wire signed [`CalcTempBus]          temp_b2_19_1_r;
wire signed [`CalcTempBus]          temp_b2_19_1_i;
wire signed [`CalcTempBus]          temp_b2_19_2_r;
wire signed [`CalcTempBus]          temp_b2_19_2_i;
wire signed [`CalcTempBus]          temp_b2_19_3_r;
wire signed [`CalcTempBus]          temp_b2_19_3_i;
wire signed [`CalcTempBus]          temp_b2_19_4_r;
wire signed [`CalcTempBus]          temp_b2_19_4_i;
wire signed [`CalcTempBus]          temp_b2_19_5_r;
wire signed [`CalcTempBus]          temp_b2_19_5_i;
wire signed [`CalcTempBus]          temp_b2_19_6_r;
wire signed [`CalcTempBus]          temp_b2_19_6_i;
wire signed [`CalcTempBus]          temp_b2_19_7_r;
wire signed [`CalcTempBus]          temp_b2_19_7_i;
wire signed [`CalcTempBus]          temp_b2_19_8_r;
wire signed [`CalcTempBus]          temp_b2_19_8_i;
wire signed [`CalcTempBus]          temp_b2_19_9_r;
wire signed [`CalcTempBus]          temp_b2_19_9_i;
wire signed [`CalcTempBus]          temp_b2_19_10_r;
wire signed [`CalcTempBus]          temp_b2_19_10_i;
wire signed [`CalcTempBus]          temp_b2_19_11_r;
wire signed [`CalcTempBus]          temp_b2_19_11_i;
wire signed [`CalcTempBus]          temp_b2_19_12_r;
wire signed [`CalcTempBus]          temp_b2_19_12_i;
wire signed [`CalcTempBus]          temp_b2_19_13_r;
wire signed [`CalcTempBus]          temp_b2_19_13_i;
wire signed [`CalcTempBus]          temp_b2_19_14_r;
wire signed [`CalcTempBus]          temp_b2_19_14_i;
wire signed [`CalcTempBus]          temp_b2_19_15_r;
wire signed [`CalcTempBus]          temp_b2_19_15_i;
wire signed [`CalcTempBus]          temp_b2_19_16_r;
wire signed [`CalcTempBus]          temp_b2_19_16_i;
wire signed [`CalcTempBus]          temp_b2_19_17_r;
wire signed [`CalcTempBus]          temp_b2_19_17_i;
wire signed [`CalcTempBus]          temp_b2_19_18_r;
wire signed [`CalcTempBus]          temp_b2_19_18_i;
wire signed [`CalcTempBus]          temp_b2_19_19_r;
wire signed [`CalcTempBus]          temp_b2_19_19_i;
wire signed [`CalcTempBus]          temp_b2_19_20_r;
wire signed [`CalcTempBus]          temp_b2_19_20_i;
wire signed [`CalcTempBus]          temp_b2_19_21_r;
wire signed [`CalcTempBus]          temp_b2_19_21_i;
wire signed [`CalcTempBus]          temp_b2_19_22_r;
wire signed [`CalcTempBus]          temp_b2_19_22_i;
wire signed [`CalcTempBus]          temp_b2_19_23_r;
wire signed [`CalcTempBus]          temp_b2_19_23_i;
wire signed [`CalcTempBus]          temp_b2_19_24_r;
wire signed [`CalcTempBus]          temp_b2_19_24_i;
wire signed [`CalcTempBus]          temp_b2_19_25_r;
wire signed [`CalcTempBus]          temp_b2_19_25_i;
wire signed [`CalcTempBus]          temp_b2_19_26_r;
wire signed [`CalcTempBus]          temp_b2_19_26_i;
wire signed [`CalcTempBus]          temp_b2_19_27_r;
wire signed [`CalcTempBus]          temp_b2_19_27_i;
wire signed [`CalcTempBus]          temp_b2_19_28_r;
wire signed [`CalcTempBus]          temp_b2_19_28_i;
wire signed [`CalcTempBus]          temp_b2_19_29_r;
wire signed [`CalcTempBus]          temp_b2_19_29_i;
wire signed [`CalcTempBus]          temp_b2_19_30_r;
wire signed [`CalcTempBus]          temp_b2_19_30_i;
wire signed [`CalcTempBus]          temp_b2_19_31_r;
wire signed [`CalcTempBus]          temp_b2_19_31_i;
wire signed [`CalcTempBus]          temp_b2_19_32_r;
wire signed [`CalcTempBus]          temp_b2_19_32_i;
wire signed [`CalcTempBus]          temp_b2_20_1_r;
wire signed [`CalcTempBus]          temp_b2_20_1_i;
wire signed [`CalcTempBus]          temp_b2_20_2_r;
wire signed [`CalcTempBus]          temp_b2_20_2_i;
wire signed [`CalcTempBus]          temp_b2_20_3_r;
wire signed [`CalcTempBus]          temp_b2_20_3_i;
wire signed [`CalcTempBus]          temp_b2_20_4_r;
wire signed [`CalcTempBus]          temp_b2_20_4_i;
wire signed [`CalcTempBus]          temp_b2_20_5_r;
wire signed [`CalcTempBus]          temp_b2_20_5_i;
wire signed [`CalcTempBus]          temp_b2_20_6_r;
wire signed [`CalcTempBus]          temp_b2_20_6_i;
wire signed [`CalcTempBus]          temp_b2_20_7_r;
wire signed [`CalcTempBus]          temp_b2_20_7_i;
wire signed [`CalcTempBus]          temp_b2_20_8_r;
wire signed [`CalcTempBus]          temp_b2_20_8_i;
wire signed [`CalcTempBus]          temp_b2_20_9_r;
wire signed [`CalcTempBus]          temp_b2_20_9_i;
wire signed [`CalcTempBus]          temp_b2_20_10_r;
wire signed [`CalcTempBus]          temp_b2_20_10_i;
wire signed [`CalcTempBus]          temp_b2_20_11_r;
wire signed [`CalcTempBus]          temp_b2_20_11_i;
wire signed [`CalcTempBus]          temp_b2_20_12_r;
wire signed [`CalcTempBus]          temp_b2_20_12_i;
wire signed [`CalcTempBus]          temp_b2_20_13_r;
wire signed [`CalcTempBus]          temp_b2_20_13_i;
wire signed [`CalcTempBus]          temp_b2_20_14_r;
wire signed [`CalcTempBus]          temp_b2_20_14_i;
wire signed [`CalcTempBus]          temp_b2_20_15_r;
wire signed [`CalcTempBus]          temp_b2_20_15_i;
wire signed [`CalcTempBus]          temp_b2_20_16_r;
wire signed [`CalcTempBus]          temp_b2_20_16_i;
wire signed [`CalcTempBus]          temp_b2_20_17_r;
wire signed [`CalcTempBus]          temp_b2_20_17_i;
wire signed [`CalcTempBus]          temp_b2_20_18_r;
wire signed [`CalcTempBus]          temp_b2_20_18_i;
wire signed [`CalcTempBus]          temp_b2_20_19_r;
wire signed [`CalcTempBus]          temp_b2_20_19_i;
wire signed [`CalcTempBus]          temp_b2_20_20_r;
wire signed [`CalcTempBus]          temp_b2_20_20_i;
wire signed [`CalcTempBus]          temp_b2_20_21_r;
wire signed [`CalcTempBus]          temp_b2_20_21_i;
wire signed [`CalcTempBus]          temp_b2_20_22_r;
wire signed [`CalcTempBus]          temp_b2_20_22_i;
wire signed [`CalcTempBus]          temp_b2_20_23_r;
wire signed [`CalcTempBus]          temp_b2_20_23_i;
wire signed [`CalcTempBus]          temp_b2_20_24_r;
wire signed [`CalcTempBus]          temp_b2_20_24_i;
wire signed [`CalcTempBus]          temp_b2_20_25_r;
wire signed [`CalcTempBus]          temp_b2_20_25_i;
wire signed [`CalcTempBus]          temp_b2_20_26_r;
wire signed [`CalcTempBus]          temp_b2_20_26_i;
wire signed [`CalcTempBus]          temp_b2_20_27_r;
wire signed [`CalcTempBus]          temp_b2_20_27_i;
wire signed [`CalcTempBus]          temp_b2_20_28_r;
wire signed [`CalcTempBus]          temp_b2_20_28_i;
wire signed [`CalcTempBus]          temp_b2_20_29_r;
wire signed [`CalcTempBus]          temp_b2_20_29_i;
wire signed [`CalcTempBus]          temp_b2_20_30_r;
wire signed [`CalcTempBus]          temp_b2_20_30_i;
wire signed [`CalcTempBus]          temp_b2_20_31_r;
wire signed [`CalcTempBus]          temp_b2_20_31_i;
wire signed [`CalcTempBus]          temp_b2_20_32_r;
wire signed [`CalcTempBus]          temp_b2_20_32_i;
wire signed [`CalcTempBus]          temp_b2_21_1_r;
wire signed [`CalcTempBus]          temp_b2_21_1_i;
wire signed [`CalcTempBus]          temp_b2_21_2_r;
wire signed [`CalcTempBus]          temp_b2_21_2_i;
wire signed [`CalcTempBus]          temp_b2_21_3_r;
wire signed [`CalcTempBus]          temp_b2_21_3_i;
wire signed [`CalcTempBus]          temp_b2_21_4_r;
wire signed [`CalcTempBus]          temp_b2_21_4_i;
wire signed [`CalcTempBus]          temp_b2_21_5_r;
wire signed [`CalcTempBus]          temp_b2_21_5_i;
wire signed [`CalcTempBus]          temp_b2_21_6_r;
wire signed [`CalcTempBus]          temp_b2_21_6_i;
wire signed [`CalcTempBus]          temp_b2_21_7_r;
wire signed [`CalcTempBus]          temp_b2_21_7_i;
wire signed [`CalcTempBus]          temp_b2_21_8_r;
wire signed [`CalcTempBus]          temp_b2_21_8_i;
wire signed [`CalcTempBus]          temp_b2_21_9_r;
wire signed [`CalcTempBus]          temp_b2_21_9_i;
wire signed [`CalcTempBus]          temp_b2_21_10_r;
wire signed [`CalcTempBus]          temp_b2_21_10_i;
wire signed [`CalcTempBus]          temp_b2_21_11_r;
wire signed [`CalcTempBus]          temp_b2_21_11_i;
wire signed [`CalcTempBus]          temp_b2_21_12_r;
wire signed [`CalcTempBus]          temp_b2_21_12_i;
wire signed [`CalcTempBus]          temp_b2_21_13_r;
wire signed [`CalcTempBus]          temp_b2_21_13_i;
wire signed [`CalcTempBus]          temp_b2_21_14_r;
wire signed [`CalcTempBus]          temp_b2_21_14_i;
wire signed [`CalcTempBus]          temp_b2_21_15_r;
wire signed [`CalcTempBus]          temp_b2_21_15_i;
wire signed [`CalcTempBus]          temp_b2_21_16_r;
wire signed [`CalcTempBus]          temp_b2_21_16_i;
wire signed [`CalcTempBus]          temp_b2_21_17_r;
wire signed [`CalcTempBus]          temp_b2_21_17_i;
wire signed [`CalcTempBus]          temp_b2_21_18_r;
wire signed [`CalcTempBus]          temp_b2_21_18_i;
wire signed [`CalcTempBus]          temp_b2_21_19_r;
wire signed [`CalcTempBus]          temp_b2_21_19_i;
wire signed [`CalcTempBus]          temp_b2_21_20_r;
wire signed [`CalcTempBus]          temp_b2_21_20_i;
wire signed [`CalcTempBus]          temp_b2_21_21_r;
wire signed [`CalcTempBus]          temp_b2_21_21_i;
wire signed [`CalcTempBus]          temp_b2_21_22_r;
wire signed [`CalcTempBus]          temp_b2_21_22_i;
wire signed [`CalcTempBus]          temp_b2_21_23_r;
wire signed [`CalcTempBus]          temp_b2_21_23_i;
wire signed [`CalcTempBus]          temp_b2_21_24_r;
wire signed [`CalcTempBus]          temp_b2_21_24_i;
wire signed [`CalcTempBus]          temp_b2_21_25_r;
wire signed [`CalcTempBus]          temp_b2_21_25_i;
wire signed [`CalcTempBus]          temp_b2_21_26_r;
wire signed [`CalcTempBus]          temp_b2_21_26_i;
wire signed [`CalcTempBus]          temp_b2_21_27_r;
wire signed [`CalcTempBus]          temp_b2_21_27_i;
wire signed [`CalcTempBus]          temp_b2_21_28_r;
wire signed [`CalcTempBus]          temp_b2_21_28_i;
wire signed [`CalcTempBus]          temp_b2_21_29_r;
wire signed [`CalcTempBus]          temp_b2_21_29_i;
wire signed [`CalcTempBus]          temp_b2_21_30_r;
wire signed [`CalcTempBus]          temp_b2_21_30_i;
wire signed [`CalcTempBus]          temp_b2_21_31_r;
wire signed [`CalcTempBus]          temp_b2_21_31_i;
wire signed [`CalcTempBus]          temp_b2_21_32_r;
wire signed [`CalcTempBus]          temp_b2_21_32_i;
wire signed [`CalcTempBus]          temp_b2_22_1_r;
wire signed [`CalcTempBus]          temp_b2_22_1_i;
wire signed [`CalcTempBus]          temp_b2_22_2_r;
wire signed [`CalcTempBus]          temp_b2_22_2_i;
wire signed [`CalcTempBus]          temp_b2_22_3_r;
wire signed [`CalcTempBus]          temp_b2_22_3_i;
wire signed [`CalcTempBus]          temp_b2_22_4_r;
wire signed [`CalcTempBus]          temp_b2_22_4_i;
wire signed [`CalcTempBus]          temp_b2_22_5_r;
wire signed [`CalcTempBus]          temp_b2_22_5_i;
wire signed [`CalcTempBus]          temp_b2_22_6_r;
wire signed [`CalcTempBus]          temp_b2_22_6_i;
wire signed [`CalcTempBus]          temp_b2_22_7_r;
wire signed [`CalcTempBus]          temp_b2_22_7_i;
wire signed [`CalcTempBus]          temp_b2_22_8_r;
wire signed [`CalcTempBus]          temp_b2_22_8_i;
wire signed [`CalcTempBus]          temp_b2_22_9_r;
wire signed [`CalcTempBus]          temp_b2_22_9_i;
wire signed [`CalcTempBus]          temp_b2_22_10_r;
wire signed [`CalcTempBus]          temp_b2_22_10_i;
wire signed [`CalcTempBus]          temp_b2_22_11_r;
wire signed [`CalcTempBus]          temp_b2_22_11_i;
wire signed [`CalcTempBus]          temp_b2_22_12_r;
wire signed [`CalcTempBus]          temp_b2_22_12_i;
wire signed [`CalcTempBus]          temp_b2_22_13_r;
wire signed [`CalcTempBus]          temp_b2_22_13_i;
wire signed [`CalcTempBus]          temp_b2_22_14_r;
wire signed [`CalcTempBus]          temp_b2_22_14_i;
wire signed [`CalcTempBus]          temp_b2_22_15_r;
wire signed [`CalcTempBus]          temp_b2_22_15_i;
wire signed [`CalcTempBus]          temp_b2_22_16_r;
wire signed [`CalcTempBus]          temp_b2_22_16_i;
wire signed [`CalcTempBus]          temp_b2_22_17_r;
wire signed [`CalcTempBus]          temp_b2_22_17_i;
wire signed [`CalcTempBus]          temp_b2_22_18_r;
wire signed [`CalcTempBus]          temp_b2_22_18_i;
wire signed [`CalcTempBus]          temp_b2_22_19_r;
wire signed [`CalcTempBus]          temp_b2_22_19_i;
wire signed [`CalcTempBus]          temp_b2_22_20_r;
wire signed [`CalcTempBus]          temp_b2_22_20_i;
wire signed [`CalcTempBus]          temp_b2_22_21_r;
wire signed [`CalcTempBus]          temp_b2_22_21_i;
wire signed [`CalcTempBus]          temp_b2_22_22_r;
wire signed [`CalcTempBus]          temp_b2_22_22_i;
wire signed [`CalcTempBus]          temp_b2_22_23_r;
wire signed [`CalcTempBus]          temp_b2_22_23_i;
wire signed [`CalcTempBus]          temp_b2_22_24_r;
wire signed [`CalcTempBus]          temp_b2_22_24_i;
wire signed [`CalcTempBus]          temp_b2_22_25_r;
wire signed [`CalcTempBus]          temp_b2_22_25_i;
wire signed [`CalcTempBus]          temp_b2_22_26_r;
wire signed [`CalcTempBus]          temp_b2_22_26_i;
wire signed [`CalcTempBus]          temp_b2_22_27_r;
wire signed [`CalcTempBus]          temp_b2_22_27_i;
wire signed [`CalcTempBus]          temp_b2_22_28_r;
wire signed [`CalcTempBus]          temp_b2_22_28_i;
wire signed [`CalcTempBus]          temp_b2_22_29_r;
wire signed [`CalcTempBus]          temp_b2_22_29_i;
wire signed [`CalcTempBus]          temp_b2_22_30_r;
wire signed [`CalcTempBus]          temp_b2_22_30_i;
wire signed [`CalcTempBus]          temp_b2_22_31_r;
wire signed [`CalcTempBus]          temp_b2_22_31_i;
wire signed [`CalcTempBus]          temp_b2_22_32_r;
wire signed [`CalcTempBus]          temp_b2_22_32_i;
wire signed [`CalcTempBus]          temp_b2_23_1_r;
wire signed [`CalcTempBus]          temp_b2_23_1_i;
wire signed [`CalcTempBus]          temp_b2_23_2_r;
wire signed [`CalcTempBus]          temp_b2_23_2_i;
wire signed [`CalcTempBus]          temp_b2_23_3_r;
wire signed [`CalcTempBus]          temp_b2_23_3_i;
wire signed [`CalcTempBus]          temp_b2_23_4_r;
wire signed [`CalcTempBus]          temp_b2_23_4_i;
wire signed [`CalcTempBus]          temp_b2_23_5_r;
wire signed [`CalcTempBus]          temp_b2_23_5_i;
wire signed [`CalcTempBus]          temp_b2_23_6_r;
wire signed [`CalcTempBus]          temp_b2_23_6_i;
wire signed [`CalcTempBus]          temp_b2_23_7_r;
wire signed [`CalcTempBus]          temp_b2_23_7_i;
wire signed [`CalcTempBus]          temp_b2_23_8_r;
wire signed [`CalcTempBus]          temp_b2_23_8_i;
wire signed [`CalcTempBus]          temp_b2_23_9_r;
wire signed [`CalcTempBus]          temp_b2_23_9_i;
wire signed [`CalcTempBus]          temp_b2_23_10_r;
wire signed [`CalcTempBus]          temp_b2_23_10_i;
wire signed [`CalcTempBus]          temp_b2_23_11_r;
wire signed [`CalcTempBus]          temp_b2_23_11_i;
wire signed [`CalcTempBus]          temp_b2_23_12_r;
wire signed [`CalcTempBus]          temp_b2_23_12_i;
wire signed [`CalcTempBus]          temp_b2_23_13_r;
wire signed [`CalcTempBus]          temp_b2_23_13_i;
wire signed [`CalcTempBus]          temp_b2_23_14_r;
wire signed [`CalcTempBus]          temp_b2_23_14_i;
wire signed [`CalcTempBus]          temp_b2_23_15_r;
wire signed [`CalcTempBus]          temp_b2_23_15_i;
wire signed [`CalcTempBus]          temp_b2_23_16_r;
wire signed [`CalcTempBus]          temp_b2_23_16_i;
wire signed [`CalcTempBus]          temp_b2_23_17_r;
wire signed [`CalcTempBus]          temp_b2_23_17_i;
wire signed [`CalcTempBus]          temp_b2_23_18_r;
wire signed [`CalcTempBus]          temp_b2_23_18_i;
wire signed [`CalcTempBus]          temp_b2_23_19_r;
wire signed [`CalcTempBus]          temp_b2_23_19_i;
wire signed [`CalcTempBus]          temp_b2_23_20_r;
wire signed [`CalcTempBus]          temp_b2_23_20_i;
wire signed [`CalcTempBus]          temp_b2_23_21_r;
wire signed [`CalcTempBus]          temp_b2_23_21_i;
wire signed [`CalcTempBus]          temp_b2_23_22_r;
wire signed [`CalcTempBus]          temp_b2_23_22_i;
wire signed [`CalcTempBus]          temp_b2_23_23_r;
wire signed [`CalcTempBus]          temp_b2_23_23_i;
wire signed [`CalcTempBus]          temp_b2_23_24_r;
wire signed [`CalcTempBus]          temp_b2_23_24_i;
wire signed [`CalcTempBus]          temp_b2_23_25_r;
wire signed [`CalcTempBus]          temp_b2_23_25_i;
wire signed [`CalcTempBus]          temp_b2_23_26_r;
wire signed [`CalcTempBus]          temp_b2_23_26_i;
wire signed [`CalcTempBus]          temp_b2_23_27_r;
wire signed [`CalcTempBus]          temp_b2_23_27_i;
wire signed [`CalcTempBus]          temp_b2_23_28_r;
wire signed [`CalcTempBus]          temp_b2_23_28_i;
wire signed [`CalcTempBus]          temp_b2_23_29_r;
wire signed [`CalcTempBus]          temp_b2_23_29_i;
wire signed [`CalcTempBus]          temp_b2_23_30_r;
wire signed [`CalcTempBus]          temp_b2_23_30_i;
wire signed [`CalcTempBus]          temp_b2_23_31_r;
wire signed [`CalcTempBus]          temp_b2_23_31_i;
wire signed [`CalcTempBus]          temp_b2_23_32_r;
wire signed [`CalcTempBus]          temp_b2_23_32_i;
wire signed [`CalcTempBus]          temp_b2_24_1_r;
wire signed [`CalcTempBus]          temp_b2_24_1_i;
wire signed [`CalcTempBus]          temp_b2_24_2_r;
wire signed [`CalcTempBus]          temp_b2_24_2_i;
wire signed [`CalcTempBus]          temp_b2_24_3_r;
wire signed [`CalcTempBus]          temp_b2_24_3_i;
wire signed [`CalcTempBus]          temp_b2_24_4_r;
wire signed [`CalcTempBus]          temp_b2_24_4_i;
wire signed [`CalcTempBus]          temp_b2_24_5_r;
wire signed [`CalcTempBus]          temp_b2_24_5_i;
wire signed [`CalcTempBus]          temp_b2_24_6_r;
wire signed [`CalcTempBus]          temp_b2_24_6_i;
wire signed [`CalcTempBus]          temp_b2_24_7_r;
wire signed [`CalcTempBus]          temp_b2_24_7_i;
wire signed [`CalcTempBus]          temp_b2_24_8_r;
wire signed [`CalcTempBus]          temp_b2_24_8_i;
wire signed [`CalcTempBus]          temp_b2_24_9_r;
wire signed [`CalcTempBus]          temp_b2_24_9_i;
wire signed [`CalcTempBus]          temp_b2_24_10_r;
wire signed [`CalcTempBus]          temp_b2_24_10_i;
wire signed [`CalcTempBus]          temp_b2_24_11_r;
wire signed [`CalcTempBus]          temp_b2_24_11_i;
wire signed [`CalcTempBus]          temp_b2_24_12_r;
wire signed [`CalcTempBus]          temp_b2_24_12_i;
wire signed [`CalcTempBus]          temp_b2_24_13_r;
wire signed [`CalcTempBus]          temp_b2_24_13_i;
wire signed [`CalcTempBus]          temp_b2_24_14_r;
wire signed [`CalcTempBus]          temp_b2_24_14_i;
wire signed [`CalcTempBus]          temp_b2_24_15_r;
wire signed [`CalcTempBus]          temp_b2_24_15_i;
wire signed [`CalcTempBus]          temp_b2_24_16_r;
wire signed [`CalcTempBus]          temp_b2_24_16_i;
wire signed [`CalcTempBus]          temp_b2_24_17_r;
wire signed [`CalcTempBus]          temp_b2_24_17_i;
wire signed [`CalcTempBus]          temp_b2_24_18_r;
wire signed [`CalcTempBus]          temp_b2_24_18_i;
wire signed [`CalcTempBus]          temp_b2_24_19_r;
wire signed [`CalcTempBus]          temp_b2_24_19_i;
wire signed [`CalcTempBus]          temp_b2_24_20_r;
wire signed [`CalcTempBus]          temp_b2_24_20_i;
wire signed [`CalcTempBus]          temp_b2_24_21_r;
wire signed [`CalcTempBus]          temp_b2_24_21_i;
wire signed [`CalcTempBus]          temp_b2_24_22_r;
wire signed [`CalcTempBus]          temp_b2_24_22_i;
wire signed [`CalcTempBus]          temp_b2_24_23_r;
wire signed [`CalcTempBus]          temp_b2_24_23_i;
wire signed [`CalcTempBus]          temp_b2_24_24_r;
wire signed [`CalcTempBus]          temp_b2_24_24_i;
wire signed [`CalcTempBus]          temp_b2_24_25_r;
wire signed [`CalcTempBus]          temp_b2_24_25_i;
wire signed [`CalcTempBus]          temp_b2_24_26_r;
wire signed [`CalcTempBus]          temp_b2_24_26_i;
wire signed [`CalcTempBus]          temp_b2_24_27_r;
wire signed [`CalcTempBus]          temp_b2_24_27_i;
wire signed [`CalcTempBus]          temp_b2_24_28_r;
wire signed [`CalcTempBus]          temp_b2_24_28_i;
wire signed [`CalcTempBus]          temp_b2_24_29_r;
wire signed [`CalcTempBus]          temp_b2_24_29_i;
wire signed [`CalcTempBus]          temp_b2_24_30_r;
wire signed [`CalcTempBus]          temp_b2_24_30_i;
wire signed [`CalcTempBus]          temp_b2_24_31_r;
wire signed [`CalcTempBus]          temp_b2_24_31_i;
wire signed [`CalcTempBus]          temp_b2_24_32_r;
wire signed [`CalcTempBus]          temp_b2_24_32_i;
wire signed [`CalcTempBus]          temp_b2_25_1_r;
wire signed [`CalcTempBus]          temp_b2_25_1_i;
wire signed [`CalcTempBus]          temp_b2_25_2_r;
wire signed [`CalcTempBus]          temp_b2_25_2_i;
wire signed [`CalcTempBus]          temp_b2_25_3_r;
wire signed [`CalcTempBus]          temp_b2_25_3_i;
wire signed [`CalcTempBus]          temp_b2_25_4_r;
wire signed [`CalcTempBus]          temp_b2_25_4_i;
wire signed [`CalcTempBus]          temp_b2_25_5_r;
wire signed [`CalcTempBus]          temp_b2_25_5_i;
wire signed [`CalcTempBus]          temp_b2_25_6_r;
wire signed [`CalcTempBus]          temp_b2_25_6_i;
wire signed [`CalcTempBus]          temp_b2_25_7_r;
wire signed [`CalcTempBus]          temp_b2_25_7_i;
wire signed [`CalcTempBus]          temp_b2_25_8_r;
wire signed [`CalcTempBus]          temp_b2_25_8_i;
wire signed [`CalcTempBus]          temp_b2_25_9_r;
wire signed [`CalcTempBus]          temp_b2_25_9_i;
wire signed [`CalcTempBus]          temp_b2_25_10_r;
wire signed [`CalcTempBus]          temp_b2_25_10_i;
wire signed [`CalcTempBus]          temp_b2_25_11_r;
wire signed [`CalcTempBus]          temp_b2_25_11_i;
wire signed [`CalcTempBus]          temp_b2_25_12_r;
wire signed [`CalcTempBus]          temp_b2_25_12_i;
wire signed [`CalcTempBus]          temp_b2_25_13_r;
wire signed [`CalcTempBus]          temp_b2_25_13_i;
wire signed [`CalcTempBus]          temp_b2_25_14_r;
wire signed [`CalcTempBus]          temp_b2_25_14_i;
wire signed [`CalcTempBus]          temp_b2_25_15_r;
wire signed [`CalcTempBus]          temp_b2_25_15_i;
wire signed [`CalcTempBus]          temp_b2_25_16_r;
wire signed [`CalcTempBus]          temp_b2_25_16_i;
wire signed [`CalcTempBus]          temp_b2_25_17_r;
wire signed [`CalcTempBus]          temp_b2_25_17_i;
wire signed [`CalcTempBus]          temp_b2_25_18_r;
wire signed [`CalcTempBus]          temp_b2_25_18_i;
wire signed [`CalcTempBus]          temp_b2_25_19_r;
wire signed [`CalcTempBus]          temp_b2_25_19_i;
wire signed [`CalcTempBus]          temp_b2_25_20_r;
wire signed [`CalcTempBus]          temp_b2_25_20_i;
wire signed [`CalcTempBus]          temp_b2_25_21_r;
wire signed [`CalcTempBus]          temp_b2_25_21_i;
wire signed [`CalcTempBus]          temp_b2_25_22_r;
wire signed [`CalcTempBus]          temp_b2_25_22_i;
wire signed [`CalcTempBus]          temp_b2_25_23_r;
wire signed [`CalcTempBus]          temp_b2_25_23_i;
wire signed [`CalcTempBus]          temp_b2_25_24_r;
wire signed [`CalcTempBus]          temp_b2_25_24_i;
wire signed [`CalcTempBus]          temp_b2_25_25_r;
wire signed [`CalcTempBus]          temp_b2_25_25_i;
wire signed [`CalcTempBus]          temp_b2_25_26_r;
wire signed [`CalcTempBus]          temp_b2_25_26_i;
wire signed [`CalcTempBus]          temp_b2_25_27_r;
wire signed [`CalcTempBus]          temp_b2_25_27_i;
wire signed [`CalcTempBus]          temp_b2_25_28_r;
wire signed [`CalcTempBus]          temp_b2_25_28_i;
wire signed [`CalcTempBus]          temp_b2_25_29_r;
wire signed [`CalcTempBus]          temp_b2_25_29_i;
wire signed [`CalcTempBus]          temp_b2_25_30_r;
wire signed [`CalcTempBus]          temp_b2_25_30_i;
wire signed [`CalcTempBus]          temp_b2_25_31_r;
wire signed [`CalcTempBus]          temp_b2_25_31_i;
wire signed [`CalcTempBus]          temp_b2_25_32_r;
wire signed [`CalcTempBus]          temp_b2_25_32_i;
wire signed [`CalcTempBus]          temp_b2_26_1_r;
wire signed [`CalcTempBus]          temp_b2_26_1_i;
wire signed [`CalcTempBus]          temp_b2_26_2_r;
wire signed [`CalcTempBus]          temp_b2_26_2_i;
wire signed [`CalcTempBus]          temp_b2_26_3_r;
wire signed [`CalcTempBus]          temp_b2_26_3_i;
wire signed [`CalcTempBus]          temp_b2_26_4_r;
wire signed [`CalcTempBus]          temp_b2_26_4_i;
wire signed [`CalcTempBus]          temp_b2_26_5_r;
wire signed [`CalcTempBus]          temp_b2_26_5_i;
wire signed [`CalcTempBus]          temp_b2_26_6_r;
wire signed [`CalcTempBus]          temp_b2_26_6_i;
wire signed [`CalcTempBus]          temp_b2_26_7_r;
wire signed [`CalcTempBus]          temp_b2_26_7_i;
wire signed [`CalcTempBus]          temp_b2_26_8_r;
wire signed [`CalcTempBus]          temp_b2_26_8_i;
wire signed [`CalcTempBus]          temp_b2_26_9_r;
wire signed [`CalcTempBus]          temp_b2_26_9_i;
wire signed [`CalcTempBus]          temp_b2_26_10_r;
wire signed [`CalcTempBus]          temp_b2_26_10_i;
wire signed [`CalcTempBus]          temp_b2_26_11_r;
wire signed [`CalcTempBus]          temp_b2_26_11_i;
wire signed [`CalcTempBus]          temp_b2_26_12_r;
wire signed [`CalcTempBus]          temp_b2_26_12_i;
wire signed [`CalcTempBus]          temp_b2_26_13_r;
wire signed [`CalcTempBus]          temp_b2_26_13_i;
wire signed [`CalcTempBus]          temp_b2_26_14_r;
wire signed [`CalcTempBus]          temp_b2_26_14_i;
wire signed [`CalcTempBus]          temp_b2_26_15_r;
wire signed [`CalcTempBus]          temp_b2_26_15_i;
wire signed [`CalcTempBus]          temp_b2_26_16_r;
wire signed [`CalcTempBus]          temp_b2_26_16_i;
wire signed [`CalcTempBus]          temp_b2_26_17_r;
wire signed [`CalcTempBus]          temp_b2_26_17_i;
wire signed [`CalcTempBus]          temp_b2_26_18_r;
wire signed [`CalcTempBus]          temp_b2_26_18_i;
wire signed [`CalcTempBus]          temp_b2_26_19_r;
wire signed [`CalcTempBus]          temp_b2_26_19_i;
wire signed [`CalcTempBus]          temp_b2_26_20_r;
wire signed [`CalcTempBus]          temp_b2_26_20_i;
wire signed [`CalcTempBus]          temp_b2_26_21_r;
wire signed [`CalcTempBus]          temp_b2_26_21_i;
wire signed [`CalcTempBus]          temp_b2_26_22_r;
wire signed [`CalcTempBus]          temp_b2_26_22_i;
wire signed [`CalcTempBus]          temp_b2_26_23_r;
wire signed [`CalcTempBus]          temp_b2_26_23_i;
wire signed [`CalcTempBus]          temp_b2_26_24_r;
wire signed [`CalcTempBus]          temp_b2_26_24_i;
wire signed [`CalcTempBus]          temp_b2_26_25_r;
wire signed [`CalcTempBus]          temp_b2_26_25_i;
wire signed [`CalcTempBus]          temp_b2_26_26_r;
wire signed [`CalcTempBus]          temp_b2_26_26_i;
wire signed [`CalcTempBus]          temp_b2_26_27_r;
wire signed [`CalcTempBus]          temp_b2_26_27_i;
wire signed [`CalcTempBus]          temp_b2_26_28_r;
wire signed [`CalcTempBus]          temp_b2_26_28_i;
wire signed [`CalcTempBus]          temp_b2_26_29_r;
wire signed [`CalcTempBus]          temp_b2_26_29_i;
wire signed [`CalcTempBus]          temp_b2_26_30_r;
wire signed [`CalcTempBus]          temp_b2_26_30_i;
wire signed [`CalcTempBus]          temp_b2_26_31_r;
wire signed [`CalcTempBus]          temp_b2_26_31_i;
wire signed [`CalcTempBus]          temp_b2_26_32_r;
wire signed [`CalcTempBus]          temp_b2_26_32_i;
wire signed [`CalcTempBus]          temp_b2_27_1_r;
wire signed [`CalcTempBus]          temp_b2_27_1_i;
wire signed [`CalcTempBus]          temp_b2_27_2_r;
wire signed [`CalcTempBus]          temp_b2_27_2_i;
wire signed [`CalcTempBus]          temp_b2_27_3_r;
wire signed [`CalcTempBus]          temp_b2_27_3_i;
wire signed [`CalcTempBus]          temp_b2_27_4_r;
wire signed [`CalcTempBus]          temp_b2_27_4_i;
wire signed [`CalcTempBus]          temp_b2_27_5_r;
wire signed [`CalcTempBus]          temp_b2_27_5_i;
wire signed [`CalcTempBus]          temp_b2_27_6_r;
wire signed [`CalcTempBus]          temp_b2_27_6_i;
wire signed [`CalcTempBus]          temp_b2_27_7_r;
wire signed [`CalcTempBus]          temp_b2_27_7_i;
wire signed [`CalcTempBus]          temp_b2_27_8_r;
wire signed [`CalcTempBus]          temp_b2_27_8_i;
wire signed [`CalcTempBus]          temp_b2_27_9_r;
wire signed [`CalcTempBus]          temp_b2_27_9_i;
wire signed [`CalcTempBus]          temp_b2_27_10_r;
wire signed [`CalcTempBus]          temp_b2_27_10_i;
wire signed [`CalcTempBus]          temp_b2_27_11_r;
wire signed [`CalcTempBus]          temp_b2_27_11_i;
wire signed [`CalcTempBus]          temp_b2_27_12_r;
wire signed [`CalcTempBus]          temp_b2_27_12_i;
wire signed [`CalcTempBus]          temp_b2_27_13_r;
wire signed [`CalcTempBus]          temp_b2_27_13_i;
wire signed [`CalcTempBus]          temp_b2_27_14_r;
wire signed [`CalcTempBus]          temp_b2_27_14_i;
wire signed [`CalcTempBus]          temp_b2_27_15_r;
wire signed [`CalcTempBus]          temp_b2_27_15_i;
wire signed [`CalcTempBus]          temp_b2_27_16_r;
wire signed [`CalcTempBus]          temp_b2_27_16_i;
wire signed [`CalcTempBus]          temp_b2_27_17_r;
wire signed [`CalcTempBus]          temp_b2_27_17_i;
wire signed [`CalcTempBus]          temp_b2_27_18_r;
wire signed [`CalcTempBus]          temp_b2_27_18_i;
wire signed [`CalcTempBus]          temp_b2_27_19_r;
wire signed [`CalcTempBus]          temp_b2_27_19_i;
wire signed [`CalcTempBus]          temp_b2_27_20_r;
wire signed [`CalcTempBus]          temp_b2_27_20_i;
wire signed [`CalcTempBus]          temp_b2_27_21_r;
wire signed [`CalcTempBus]          temp_b2_27_21_i;
wire signed [`CalcTempBus]          temp_b2_27_22_r;
wire signed [`CalcTempBus]          temp_b2_27_22_i;
wire signed [`CalcTempBus]          temp_b2_27_23_r;
wire signed [`CalcTempBus]          temp_b2_27_23_i;
wire signed [`CalcTempBus]          temp_b2_27_24_r;
wire signed [`CalcTempBus]          temp_b2_27_24_i;
wire signed [`CalcTempBus]          temp_b2_27_25_r;
wire signed [`CalcTempBus]          temp_b2_27_25_i;
wire signed [`CalcTempBus]          temp_b2_27_26_r;
wire signed [`CalcTempBus]          temp_b2_27_26_i;
wire signed [`CalcTempBus]          temp_b2_27_27_r;
wire signed [`CalcTempBus]          temp_b2_27_27_i;
wire signed [`CalcTempBus]          temp_b2_27_28_r;
wire signed [`CalcTempBus]          temp_b2_27_28_i;
wire signed [`CalcTempBus]          temp_b2_27_29_r;
wire signed [`CalcTempBus]          temp_b2_27_29_i;
wire signed [`CalcTempBus]          temp_b2_27_30_r;
wire signed [`CalcTempBus]          temp_b2_27_30_i;
wire signed [`CalcTempBus]          temp_b2_27_31_r;
wire signed [`CalcTempBus]          temp_b2_27_31_i;
wire signed [`CalcTempBus]          temp_b2_27_32_r;
wire signed [`CalcTempBus]          temp_b2_27_32_i;
wire signed [`CalcTempBus]          temp_b2_28_1_r;
wire signed [`CalcTempBus]          temp_b2_28_1_i;
wire signed [`CalcTempBus]          temp_b2_28_2_r;
wire signed [`CalcTempBus]          temp_b2_28_2_i;
wire signed [`CalcTempBus]          temp_b2_28_3_r;
wire signed [`CalcTempBus]          temp_b2_28_3_i;
wire signed [`CalcTempBus]          temp_b2_28_4_r;
wire signed [`CalcTempBus]          temp_b2_28_4_i;
wire signed [`CalcTempBus]          temp_b2_28_5_r;
wire signed [`CalcTempBus]          temp_b2_28_5_i;
wire signed [`CalcTempBus]          temp_b2_28_6_r;
wire signed [`CalcTempBus]          temp_b2_28_6_i;
wire signed [`CalcTempBus]          temp_b2_28_7_r;
wire signed [`CalcTempBus]          temp_b2_28_7_i;
wire signed [`CalcTempBus]          temp_b2_28_8_r;
wire signed [`CalcTempBus]          temp_b2_28_8_i;
wire signed [`CalcTempBus]          temp_b2_28_9_r;
wire signed [`CalcTempBus]          temp_b2_28_9_i;
wire signed [`CalcTempBus]          temp_b2_28_10_r;
wire signed [`CalcTempBus]          temp_b2_28_10_i;
wire signed [`CalcTempBus]          temp_b2_28_11_r;
wire signed [`CalcTempBus]          temp_b2_28_11_i;
wire signed [`CalcTempBus]          temp_b2_28_12_r;
wire signed [`CalcTempBus]          temp_b2_28_12_i;
wire signed [`CalcTempBus]          temp_b2_28_13_r;
wire signed [`CalcTempBus]          temp_b2_28_13_i;
wire signed [`CalcTempBus]          temp_b2_28_14_r;
wire signed [`CalcTempBus]          temp_b2_28_14_i;
wire signed [`CalcTempBus]          temp_b2_28_15_r;
wire signed [`CalcTempBus]          temp_b2_28_15_i;
wire signed [`CalcTempBus]          temp_b2_28_16_r;
wire signed [`CalcTempBus]          temp_b2_28_16_i;
wire signed [`CalcTempBus]          temp_b2_28_17_r;
wire signed [`CalcTempBus]          temp_b2_28_17_i;
wire signed [`CalcTempBus]          temp_b2_28_18_r;
wire signed [`CalcTempBus]          temp_b2_28_18_i;
wire signed [`CalcTempBus]          temp_b2_28_19_r;
wire signed [`CalcTempBus]          temp_b2_28_19_i;
wire signed [`CalcTempBus]          temp_b2_28_20_r;
wire signed [`CalcTempBus]          temp_b2_28_20_i;
wire signed [`CalcTempBus]          temp_b2_28_21_r;
wire signed [`CalcTempBus]          temp_b2_28_21_i;
wire signed [`CalcTempBus]          temp_b2_28_22_r;
wire signed [`CalcTempBus]          temp_b2_28_22_i;
wire signed [`CalcTempBus]          temp_b2_28_23_r;
wire signed [`CalcTempBus]          temp_b2_28_23_i;
wire signed [`CalcTempBus]          temp_b2_28_24_r;
wire signed [`CalcTempBus]          temp_b2_28_24_i;
wire signed [`CalcTempBus]          temp_b2_28_25_r;
wire signed [`CalcTempBus]          temp_b2_28_25_i;
wire signed [`CalcTempBus]          temp_b2_28_26_r;
wire signed [`CalcTempBus]          temp_b2_28_26_i;
wire signed [`CalcTempBus]          temp_b2_28_27_r;
wire signed [`CalcTempBus]          temp_b2_28_27_i;
wire signed [`CalcTempBus]          temp_b2_28_28_r;
wire signed [`CalcTempBus]          temp_b2_28_28_i;
wire signed [`CalcTempBus]          temp_b2_28_29_r;
wire signed [`CalcTempBus]          temp_b2_28_29_i;
wire signed [`CalcTempBus]          temp_b2_28_30_r;
wire signed [`CalcTempBus]          temp_b2_28_30_i;
wire signed [`CalcTempBus]          temp_b2_28_31_r;
wire signed [`CalcTempBus]          temp_b2_28_31_i;
wire signed [`CalcTempBus]          temp_b2_28_32_r;
wire signed [`CalcTempBus]          temp_b2_28_32_i;
wire signed [`CalcTempBus]          temp_b2_29_1_r;
wire signed [`CalcTempBus]          temp_b2_29_1_i;
wire signed [`CalcTempBus]          temp_b2_29_2_r;
wire signed [`CalcTempBus]          temp_b2_29_2_i;
wire signed [`CalcTempBus]          temp_b2_29_3_r;
wire signed [`CalcTempBus]          temp_b2_29_3_i;
wire signed [`CalcTempBus]          temp_b2_29_4_r;
wire signed [`CalcTempBus]          temp_b2_29_4_i;
wire signed [`CalcTempBus]          temp_b2_29_5_r;
wire signed [`CalcTempBus]          temp_b2_29_5_i;
wire signed [`CalcTempBus]          temp_b2_29_6_r;
wire signed [`CalcTempBus]          temp_b2_29_6_i;
wire signed [`CalcTempBus]          temp_b2_29_7_r;
wire signed [`CalcTempBus]          temp_b2_29_7_i;
wire signed [`CalcTempBus]          temp_b2_29_8_r;
wire signed [`CalcTempBus]          temp_b2_29_8_i;
wire signed [`CalcTempBus]          temp_b2_29_9_r;
wire signed [`CalcTempBus]          temp_b2_29_9_i;
wire signed [`CalcTempBus]          temp_b2_29_10_r;
wire signed [`CalcTempBus]          temp_b2_29_10_i;
wire signed [`CalcTempBus]          temp_b2_29_11_r;
wire signed [`CalcTempBus]          temp_b2_29_11_i;
wire signed [`CalcTempBus]          temp_b2_29_12_r;
wire signed [`CalcTempBus]          temp_b2_29_12_i;
wire signed [`CalcTempBus]          temp_b2_29_13_r;
wire signed [`CalcTempBus]          temp_b2_29_13_i;
wire signed [`CalcTempBus]          temp_b2_29_14_r;
wire signed [`CalcTempBus]          temp_b2_29_14_i;
wire signed [`CalcTempBus]          temp_b2_29_15_r;
wire signed [`CalcTempBus]          temp_b2_29_15_i;
wire signed [`CalcTempBus]          temp_b2_29_16_r;
wire signed [`CalcTempBus]          temp_b2_29_16_i;
wire signed [`CalcTempBus]          temp_b2_29_17_r;
wire signed [`CalcTempBus]          temp_b2_29_17_i;
wire signed [`CalcTempBus]          temp_b2_29_18_r;
wire signed [`CalcTempBus]          temp_b2_29_18_i;
wire signed [`CalcTempBus]          temp_b2_29_19_r;
wire signed [`CalcTempBus]          temp_b2_29_19_i;
wire signed [`CalcTempBus]          temp_b2_29_20_r;
wire signed [`CalcTempBus]          temp_b2_29_20_i;
wire signed [`CalcTempBus]          temp_b2_29_21_r;
wire signed [`CalcTempBus]          temp_b2_29_21_i;
wire signed [`CalcTempBus]          temp_b2_29_22_r;
wire signed [`CalcTempBus]          temp_b2_29_22_i;
wire signed [`CalcTempBus]          temp_b2_29_23_r;
wire signed [`CalcTempBus]          temp_b2_29_23_i;
wire signed [`CalcTempBus]          temp_b2_29_24_r;
wire signed [`CalcTempBus]          temp_b2_29_24_i;
wire signed [`CalcTempBus]          temp_b2_29_25_r;
wire signed [`CalcTempBus]          temp_b2_29_25_i;
wire signed [`CalcTempBus]          temp_b2_29_26_r;
wire signed [`CalcTempBus]          temp_b2_29_26_i;
wire signed [`CalcTempBus]          temp_b2_29_27_r;
wire signed [`CalcTempBus]          temp_b2_29_27_i;
wire signed [`CalcTempBus]          temp_b2_29_28_r;
wire signed [`CalcTempBus]          temp_b2_29_28_i;
wire signed [`CalcTempBus]          temp_b2_29_29_r;
wire signed [`CalcTempBus]          temp_b2_29_29_i;
wire signed [`CalcTempBus]          temp_b2_29_30_r;
wire signed [`CalcTempBus]          temp_b2_29_30_i;
wire signed [`CalcTempBus]          temp_b2_29_31_r;
wire signed [`CalcTempBus]          temp_b2_29_31_i;
wire signed [`CalcTempBus]          temp_b2_29_32_r;
wire signed [`CalcTempBus]          temp_b2_29_32_i;
wire signed [`CalcTempBus]          temp_b2_30_1_r;
wire signed [`CalcTempBus]          temp_b2_30_1_i;
wire signed [`CalcTempBus]          temp_b2_30_2_r;
wire signed [`CalcTempBus]          temp_b2_30_2_i;
wire signed [`CalcTempBus]          temp_b2_30_3_r;
wire signed [`CalcTempBus]          temp_b2_30_3_i;
wire signed [`CalcTempBus]          temp_b2_30_4_r;
wire signed [`CalcTempBus]          temp_b2_30_4_i;
wire signed [`CalcTempBus]          temp_b2_30_5_r;
wire signed [`CalcTempBus]          temp_b2_30_5_i;
wire signed [`CalcTempBus]          temp_b2_30_6_r;
wire signed [`CalcTempBus]          temp_b2_30_6_i;
wire signed [`CalcTempBus]          temp_b2_30_7_r;
wire signed [`CalcTempBus]          temp_b2_30_7_i;
wire signed [`CalcTempBus]          temp_b2_30_8_r;
wire signed [`CalcTempBus]          temp_b2_30_8_i;
wire signed [`CalcTempBus]          temp_b2_30_9_r;
wire signed [`CalcTempBus]          temp_b2_30_9_i;
wire signed [`CalcTempBus]          temp_b2_30_10_r;
wire signed [`CalcTempBus]          temp_b2_30_10_i;
wire signed [`CalcTempBus]          temp_b2_30_11_r;
wire signed [`CalcTempBus]          temp_b2_30_11_i;
wire signed [`CalcTempBus]          temp_b2_30_12_r;
wire signed [`CalcTempBus]          temp_b2_30_12_i;
wire signed [`CalcTempBus]          temp_b2_30_13_r;
wire signed [`CalcTempBus]          temp_b2_30_13_i;
wire signed [`CalcTempBus]          temp_b2_30_14_r;
wire signed [`CalcTempBus]          temp_b2_30_14_i;
wire signed [`CalcTempBus]          temp_b2_30_15_r;
wire signed [`CalcTempBus]          temp_b2_30_15_i;
wire signed [`CalcTempBus]          temp_b2_30_16_r;
wire signed [`CalcTempBus]          temp_b2_30_16_i;
wire signed [`CalcTempBus]          temp_b2_30_17_r;
wire signed [`CalcTempBus]          temp_b2_30_17_i;
wire signed [`CalcTempBus]          temp_b2_30_18_r;
wire signed [`CalcTempBus]          temp_b2_30_18_i;
wire signed [`CalcTempBus]          temp_b2_30_19_r;
wire signed [`CalcTempBus]          temp_b2_30_19_i;
wire signed [`CalcTempBus]          temp_b2_30_20_r;
wire signed [`CalcTempBus]          temp_b2_30_20_i;
wire signed [`CalcTempBus]          temp_b2_30_21_r;
wire signed [`CalcTempBus]          temp_b2_30_21_i;
wire signed [`CalcTempBus]          temp_b2_30_22_r;
wire signed [`CalcTempBus]          temp_b2_30_22_i;
wire signed [`CalcTempBus]          temp_b2_30_23_r;
wire signed [`CalcTempBus]          temp_b2_30_23_i;
wire signed [`CalcTempBus]          temp_b2_30_24_r;
wire signed [`CalcTempBus]          temp_b2_30_24_i;
wire signed [`CalcTempBus]          temp_b2_30_25_r;
wire signed [`CalcTempBus]          temp_b2_30_25_i;
wire signed [`CalcTempBus]          temp_b2_30_26_r;
wire signed [`CalcTempBus]          temp_b2_30_26_i;
wire signed [`CalcTempBus]          temp_b2_30_27_r;
wire signed [`CalcTempBus]          temp_b2_30_27_i;
wire signed [`CalcTempBus]          temp_b2_30_28_r;
wire signed [`CalcTempBus]          temp_b2_30_28_i;
wire signed [`CalcTempBus]          temp_b2_30_29_r;
wire signed [`CalcTempBus]          temp_b2_30_29_i;
wire signed [`CalcTempBus]          temp_b2_30_30_r;
wire signed [`CalcTempBus]          temp_b2_30_30_i;
wire signed [`CalcTempBus]          temp_b2_30_31_r;
wire signed [`CalcTempBus]          temp_b2_30_31_i;
wire signed [`CalcTempBus]          temp_b2_30_32_r;
wire signed [`CalcTempBus]          temp_b2_30_32_i;
wire signed [`CalcTempBus]          temp_b2_31_1_r;
wire signed [`CalcTempBus]          temp_b2_31_1_i;
wire signed [`CalcTempBus]          temp_b2_31_2_r;
wire signed [`CalcTempBus]          temp_b2_31_2_i;
wire signed [`CalcTempBus]          temp_b2_31_3_r;
wire signed [`CalcTempBus]          temp_b2_31_3_i;
wire signed [`CalcTempBus]          temp_b2_31_4_r;
wire signed [`CalcTempBus]          temp_b2_31_4_i;
wire signed [`CalcTempBus]          temp_b2_31_5_r;
wire signed [`CalcTempBus]          temp_b2_31_5_i;
wire signed [`CalcTempBus]          temp_b2_31_6_r;
wire signed [`CalcTempBus]          temp_b2_31_6_i;
wire signed [`CalcTempBus]          temp_b2_31_7_r;
wire signed [`CalcTempBus]          temp_b2_31_7_i;
wire signed [`CalcTempBus]          temp_b2_31_8_r;
wire signed [`CalcTempBus]          temp_b2_31_8_i;
wire signed [`CalcTempBus]          temp_b2_31_9_r;
wire signed [`CalcTempBus]          temp_b2_31_9_i;
wire signed [`CalcTempBus]          temp_b2_31_10_r;
wire signed [`CalcTempBus]          temp_b2_31_10_i;
wire signed [`CalcTempBus]          temp_b2_31_11_r;
wire signed [`CalcTempBus]          temp_b2_31_11_i;
wire signed [`CalcTempBus]          temp_b2_31_12_r;
wire signed [`CalcTempBus]          temp_b2_31_12_i;
wire signed [`CalcTempBus]          temp_b2_31_13_r;
wire signed [`CalcTempBus]          temp_b2_31_13_i;
wire signed [`CalcTempBus]          temp_b2_31_14_r;
wire signed [`CalcTempBus]          temp_b2_31_14_i;
wire signed [`CalcTempBus]          temp_b2_31_15_r;
wire signed [`CalcTempBus]          temp_b2_31_15_i;
wire signed [`CalcTempBus]          temp_b2_31_16_r;
wire signed [`CalcTempBus]          temp_b2_31_16_i;
wire signed [`CalcTempBus]          temp_b2_31_17_r;
wire signed [`CalcTempBus]          temp_b2_31_17_i;
wire signed [`CalcTempBus]          temp_b2_31_18_r;
wire signed [`CalcTempBus]          temp_b2_31_18_i;
wire signed [`CalcTempBus]          temp_b2_31_19_r;
wire signed [`CalcTempBus]          temp_b2_31_19_i;
wire signed [`CalcTempBus]          temp_b2_31_20_r;
wire signed [`CalcTempBus]          temp_b2_31_20_i;
wire signed [`CalcTempBus]          temp_b2_31_21_r;
wire signed [`CalcTempBus]          temp_b2_31_21_i;
wire signed [`CalcTempBus]          temp_b2_31_22_r;
wire signed [`CalcTempBus]          temp_b2_31_22_i;
wire signed [`CalcTempBus]          temp_b2_31_23_r;
wire signed [`CalcTempBus]          temp_b2_31_23_i;
wire signed [`CalcTempBus]          temp_b2_31_24_r;
wire signed [`CalcTempBus]          temp_b2_31_24_i;
wire signed [`CalcTempBus]          temp_b2_31_25_r;
wire signed [`CalcTempBus]          temp_b2_31_25_i;
wire signed [`CalcTempBus]          temp_b2_31_26_r;
wire signed [`CalcTempBus]          temp_b2_31_26_i;
wire signed [`CalcTempBus]          temp_b2_31_27_r;
wire signed [`CalcTempBus]          temp_b2_31_27_i;
wire signed [`CalcTempBus]          temp_b2_31_28_r;
wire signed [`CalcTempBus]          temp_b2_31_28_i;
wire signed [`CalcTempBus]          temp_b2_31_29_r;
wire signed [`CalcTempBus]          temp_b2_31_29_i;
wire signed [`CalcTempBus]          temp_b2_31_30_r;
wire signed [`CalcTempBus]          temp_b2_31_30_i;
wire signed [`CalcTempBus]          temp_b2_31_31_r;
wire signed [`CalcTempBus]          temp_b2_31_31_i;
wire signed [`CalcTempBus]          temp_b2_31_32_r;
wire signed [`CalcTempBus]          temp_b2_31_32_i;
wire signed [`CalcTempBus]          temp_b2_32_1_r;
wire signed [`CalcTempBus]          temp_b2_32_1_i;
wire signed [`CalcTempBus]          temp_b2_32_2_r;
wire signed [`CalcTempBus]          temp_b2_32_2_i;
wire signed [`CalcTempBus]          temp_b2_32_3_r;
wire signed [`CalcTempBus]          temp_b2_32_3_i;
wire signed [`CalcTempBus]          temp_b2_32_4_r;
wire signed [`CalcTempBus]          temp_b2_32_4_i;
wire signed [`CalcTempBus]          temp_b2_32_5_r;
wire signed [`CalcTempBus]          temp_b2_32_5_i;
wire signed [`CalcTempBus]          temp_b2_32_6_r;
wire signed [`CalcTempBus]          temp_b2_32_6_i;
wire signed [`CalcTempBus]          temp_b2_32_7_r;
wire signed [`CalcTempBus]          temp_b2_32_7_i;
wire signed [`CalcTempBus]          temp_b2_32_8_r;
wire signed [`CalcTempBus]          temp_b2_32_8_i;
wire signed [`CalcTempBus]          temp_b2_32_9_r;
wire signed [`CalcTempBus]          temp_b2_32_9_i;
wire signed [`CalcTempBus]          temp_b2_32_10_r;
wire signed [`CalcTempBus]          temp_b2_32_10_i;
wire signed [`CalcTempBus]          temp_b2_32_11_r;
wire signed [`CalcTempBus]          temp_b2_32_11_i;
wire signed [`CalcTempBus]          temp_b2_32_12_r;
wire signed [`CalcTempBus]          temp_b2_32_12_i;
wire signed [`CalcTempBus]          temp_b2_32_13_r;
wire signed [`CalcTempBus]          temp_b2_32_13_i;
wire signed [`CalcTempBus]          temp_b2_32_14_r;
wire signed [`CalcTempBus]          temp_b2_32_14_i;
wire signed [`CalcTempBus]          temp_b2_32_15_r;
wire signed [`CalcTempBus]          temp_b2_32_15_i;
wire signed [`CalcTempBus]          temp_b2_32_16_r;
wire signed [`CalcTempBus]          temp_b2_32_16_i;
wire signed [`CalcTempBus]          temp_b2_32_17_r;
wire signed [`CalcTempBus]          temp_b2_32_17_i;
wire signed [`CalcTempBus]          temp_b2_32_18_r;
wire signed [`CalcTempBus]          temp_b2_32_18_i;
wire signed [`CalcTempBus]          temp_b2_32_19_r;
wire signed [`CalcTempBus]          temp_b2_32_19_i;
wire signed [`CalcTempBus]          temp_b2_32_20_r;
wire signed [`CalcTempBus]          temp_b2_32_20_i;
wire signed [`CalcTempBus]          temp_b2_32_21_r;
wire signed [`CalcTempBus]          temp_b2_32_21_i;
wire signed [`CalcTempBus]          temp_b2_32_22_r;
wire signed [`CalcTempBus]          temp_b2_32_22_i;
wire signed [`CalcTempBus]          temp_b2_32_23_r;
wire signed [`CalcTempBus]          temp_b2_32_23_i;
wire signed [`CalcTempBus]          temp_b2_32_24_r;
wire signed [`CalcTempBus]          temp_b2_32_24_i;
wire signed [`CalcTempBus]          temp_b2_32_25_r;
wire signed [`CalcTempBus]          temp_b2_32_25_i;
wire signed [`CalcTempBus]          temp_b2_32_26_r;
wire signed [`CalcTempBus]          temp_b2_32_26_i;
wire signed [`CalcTempBus]          temp_b2_32_27_r;
wire signed [`CalcTempBus]          temp_b2_32_27_i;
wire signed [`CalcTempBus]          temp_b2_32_28_r;
wire signed [`CalcTempBus]          temp_b2_32_28_i;
wire signed [`CalcTempBus]          temp_b2_32_29_r;
wire signed [`CalcTempBus]          temp_b2_32_29_i;
wire signed [`CalcTempBus]          temp_b2_32_30_r;
wire signed [`CalcTempBus]          temp_b2_32_30_i;
wire signed [`CalcTempBus]          temp_b2_32_31_r;
wire signed [`CalcTempBus]          temp_b2_32_31_i;
wire signed [`CalcTempBus]          temp_b2_32_32_r;
wire signed [`CalcTempBus]          temp_b2_32_32_i;
wire signed [`CalcTempBus]          temp_b3_1_1_r;
wire signed [`CalcTempBus]          temp_b3_1_1_i;
wire signed [`CalcTempBus]          temp_b3_1_2_r;
wire signed [`CalcTempBus]          temp_b3_1_2_i;
wire signed [`CalcTempBus]          temp_b3_1_3_r;
wire signed [`CalcTempBus]          temp_b3_1_3_i;
wire signed [`CalcTempBus]          temp_b3_1_4_r;
wire signed [`CalcTempBus]          temp_b3_1_4_i;
wire signed [`CalcTempBus]          temp_b3_1_5_r;
wire signed [`CalcTempBus]          temp_b3_1_5_i;
wire signed [`CalcTempBus]          temp_b3_1_6_r;
wire signed [`CalcTempBus]          temp_b3_1_6_i;
wire signed [`CalcTempBus]          temp_b3_1_7_r;
wire signed [`CalcTempBus]          temp_b3_1_7_i;
wire signed [`CalcTempBus]          temp_b3_1_8_r;
wire signed [`CalcTempBus]          temp_b3_1_8_i;
wire signed [`CalcTempBus]          temp_b3_1_9_r;
wire signed [`CalcTempBus]          temp_b3_1_9_i;
wire signed [`CalcTempBus]          temp_b3_1_10_r;
wire signed [`CalcTempBus]          temp_b3_1_10_i;
wire signed [`CalcTempBus]          temp_b3_1_11_r;
wire signed [`CalcTempBus]          temp_b3_1_11_i;
wire signed [`CalcTempBus]          temp_b3_1_12_r;
wire signed [`CalcTempBus]          temp_b3_1_12_i;
wire signed [`CalcTempBus]          temp_b3_1_13_r;
wire signed [`CalcTempBus]          temp_b3_1_13_i;
wire signed [`CalcTempBus]          temp_b3_1_14_r;
wire signed [`CalcTempBus]          temp_b3_1_14_i;
wire signed [`CalcTempBus]          temp_b3_1_15_r;
wire signed [`CalcTempBus]          temp_b3_1_15_i;
wire signed [`CalcTempBus]          temp_b3_1_16_r;
wire signed [`CalcTempBus]          temp_b3_1_16_i;
wire signed [`CalcTempBus]          temp_b3_1_17_r;
wire signed [`CalcTempBus]          temp_b3_1_17_i;
wire signed [`CalcTempBus]          temp_b3_1_18_r;
wire signed [`CalcTempBus]          temp_b3_1_18_i;
wire signed [`CalcTempBus]          temp_b3_1_19_r;
wire signed [`CalcTempBus]          temp_b3_1_19_i;
wire signed [`CalcTempBus]          temp_b3_1_20_r;
wire signed [`CalcTempBus]          temp_b3_1_20_i;
wire signed [`CalcTempBus]          temp_b3_1_21_r;
wire signed [`CalcTempBus]          temp_b3_1_21_i;
wire signed [`CalcTempBus]          temp_b3_1_22_r;
wire signed [`CalcTempBus]          temp_b3_1_22_i;
wire signed [`CalcTempBus]          temp_b3_1_23_r;
wire signed [`CalcTempBus]          temp_b3_1_23_i;
wire signed [`CalcTempBus]          temp_b3_1_24_r;
wire signed [`CalcTempBus]          temp_b3_1_24_i;
wire signed [`CalcTempBus]          temp_b3_1_25_r;
wire signed [`CalcTempBus]          temp_b3_1_25_i;
wire signed [`CalcTempBus]          temp_b3_1_26_r;
wire signed [`CalcTempBus]          temp_b3_1_26_i;
wire signed [`CalcTempBus]          temp_b3_1_27_r;
wire signed [`CalcTempBus]          temp_b3_1_27_i;
wire signed [`CalcTempBus]          temp_b3_1_28_r;
wire signed [`CalcTempBus]          temp_b3_1_28_i;
wire signed [`CalcTempBus]          temp_b3_1_29_r;
wire signed [`CalcTempBus]          temp_b3_1_29_i;
wire signed [`CalcTempBus]          temp_b3_1_30_r;
wire signed [`CalcTempBus]          temp_b3_1_30_i;
wire signed [`CalcTempBus]          temp_b3_1_31_r;
wire signed [`CalcTempBus]          temp_b3_1_31_i;
wire signed [`CalcTempBus]          temp_b3_1_32_r;
wire signed [`CalcTempBus]          temp_b3_1_32_i;
wire signed [`CalcTempBus]          temp_b3_2_1_r;
wire signed [`CalcTempBus]          temp_b3_2_1_i;
wire signed [`CalcTempBus]          temp_b3_2_2_r;
wire signed [`CalcTempBus]          temp_b3_2_2_i;
wire signed [`CalcTempBus]          temp_b3_2_3_r;
wire signed [`CalcTempBus]          temp_b3_2_3_i;
wire signed [`CalcTempBus]          temp_b3_2_4_r;
wire signed [`CalcTempBus]          temp_b3_2_4_i;
wire signed [`CalcTempBus]          temp_b3_2_5_r;
wire signed [`CalcTempBus]          temp_b3_2_5_i;
wire signed [`CalcTempBus]          temp_b3_2_6_r;
wire signed [`CalcTempBus]          temp_b3_2_6_i;
wire signed [`CalcTempBus]          temp_b3_2_7_r;
wire signed [`CalcTempBus]          temp_b3_2_7_i;
wire signed [`CalcTempBus]          temp_b3_2_8_r;
wire signed [`CalcTempBus]          temp_b3_2_8_i;
wire signed [`CalcTempBus]          temp_b3_2_9_r;
wire signed [`CalcTempBus]          temp_b3_2_9_i;
wire signed [`CalcTempBus]          temp_b3_2_10_r;
wire signed [`CalcTempBus]          temp_b3_2_10_i;
wire signed [`CalcTempBus]          temp_b3_2_11_r;
wire signed [`CalcTempBus]          temp_b3_2_11_i;
wire signed [`CalcTempBus]          temp_b3_2_12_r;
wire signed [`CalcTempBus]          temp_b3_2_12_i;
wire signed [`CalcTempBus]          temp_b3_2_13_r;
wire signed [`CalcTempBus]          temp_b3_2_13_i;
wire signed [`CalcTempBus]          temp_b3_2_14_r;
wire signed [`CalcTempBus]          temp_b3_2_14_i;
wire signed [`CalcTempBus]          temp_b3_2_15_r;
wire signed [`CalcTempBus]          temp_b3_2_15_i;
wire signed [`CalcTempBus]          temp_b3_2_16_r;
wire signed [`CalcTempBus]          temp_b3_2_16_i;
wire signed [`CalcTempBus]          temp_b3_2_17_r;
wire signed [`CalcTempBus]          temp_b3_2_17_i;
wire signed [`CalcTempBus]          temp_b3_2_18_r;
wire signed [`CalcTempBus]          temp_b3_2_18_i;
wire signed [`CalcTempBus]          temp_b3_2_19_r;
wire signed [`CalcTempBus]          temp_b3_2_19_i;
wire signed [`CalcTempBus]          temp_b3_2_20_r;
wire signed [`CalcTempBus]          temp_b3_2_20_i;
wire signed [`CalcTempBus]          temp_b3_2_21_r;
wire signed [`CalcTempBus]          temp_b3_2_21_i;
wire signed [`CalcTempBus]          temp_b3_2_22_r;
wire signed [`CalcTempBus]          temp_b3_2_22_i;
wire signed [`CalcTempBus]          temp_b3_2_23_r;
wire signed [`CalcTempBus]          temp_b3_2_23_i;
wire signed [`CalcTempBus]          temp_b3_2_24_r;
wire signed [`CalcTempBus]          temp_b3_2_24_i;
wire signed [`CalcTempBus]          temp_b3_2_25_r;
wire signed [`CalcTempBus]          temp_b3_2_25_i;
wire signed [`CalcTempBus]          temp_b3_2_26_r;
wire signed [`CalcTempBus]          temp_b3_2_26_i;
wire signed [`CalcTempBus]          temp_b3_2_27_r;
wire signed [`CalcTempBus]          temp_b3_2_27_i;
wire signed [`CalcTempBus]          temp_b3_2_28_r;
wire signed [`CalcTempBus]          temp_b3_2_28_i;
wire signed [`CalcTempBus]          temp_b3_2_29_r;
wire signed [`CalcTempBus]          temp_b3_2_29_i;
wire signed [`CalcTempBus]          temp_b3_2_30_r;
wire signed [`CalcTempBus]          temp_b3_2_30_i;
wire signed [`CalcTempBus]          temp_b3_2_31_r;
wire signed [`CalcTempBus]          temp_b3_2_31_i;
wire signed [`CalcTempBus]          temp_b3_2_32_r;
wire signed [`CalcTempBus]          temp_b3_2_32_i;
wire signed [`CalcTempBus]          temp_b3_3_1_r;
wire signed [`CalcTempBus]          temp_b3_3_1_i;
wire signed [`CalcTempBus]          temp_b3_3_2_r;
wire signed [`CalcTempBus]          temp_b3_3_2_i;
wire signed [`CalcTempBus]          temp_b3_3_3_r;
wire signed [`CalcTempBus]          temp_b3_3_3_i;
wire signed [`CalcTempBus]          temp_b3_3_4_r;
wire signed [`CalcTempBus]          temp_b3_3_4_i;
wire signed [`CalcTempBus]          temp_b3_3_5_r;
wire signed [`CalcTempBus]          temp_b3_3_5_i;
wire signed [`CalcTempBus]          temp_b3_3_6_r;
wire signed [`CalcTempBus]          temp_b3_3_6_i;
wire signed [`CalcTempBus]          temp_b3_3_7_r;
wire signed [`CalcTempBus]          temp_b3_3_7_i;
wire signed [`CalcTempBus]          temp_b3_3_8_r;
wire signed [`CalcTempBus]          temp_b3_3_8_i;
wire signed [`CalcTempBus]          temp_b3_3_9_r;
wire signed [`CalcTempBus]          temp_b3_3_9_i;
wire signed [`CalcTempBus]          temp_b3_3_10_r;
wire signed [`CalcTempBus]          temp_b3_3_10_i;
wire signed [`CalcTempBus]          temp_b3_3_11_r;
wire signed [`CalcTempBus]          temp_b3_3_11_i;
wire signed [`CalcTempBus]          temp_b3_3_12_r;
wire signed [`CalcTempBus]          temp_b3_3_12_i;
wire signed [`CalcTempBus]          temp_b3_3_13_r;
wire signed [`CalcTempBus]          temp_b3_3_13_i;
wire signed [`CalcTempBus]          temp_b3_3_14_r;
wire signed [`CalcTempBus]          temp_b3_3_14_i;
wire signed [`CalcTempBus]          temp_b3_3_15_r;
wire signed [`CalcTempBus]          temp_b3_3_15_i;
wire signed [`CalcTempBus]          temp_b3_3_16_r;
wire signed [`CalcTempBus]          temp_b3_3_16_i;
wire signed [`CalcTempBus]          temp_b3_3_17_r;
wire signed [`CalcTempBus]          temp_b3_3_17_i;
wire signed [`CalcTempBus]          temp_b3_3_18_r;
wire signed [`CalcTempBus]          temp_b3_3_18_i;
wire signed [`CalcTempBus]          temp_b3_3_19_r;
wire signed [`CalcTempBus]          temp_b3_3_19_i;
wire signed [`CalcTempBus]          temp_b3_3_20_r;
wire signed [`CalcTempBus]          temp_b3_3_20_i;
wire signed [`CalcTempBus]          temp_b3_3_21_r;
wire signed [`CalcTempBus]          temp_b3_3_21_i;
wire signed [`CalcTempBus]          temp_b3_3_22_r;
wire signed [`CalcTempBus]          temp_b3_3_22_i;
wire signed [`CalcTempBus]          temp_b3_3_23_r;
wire signed [`CalcTempBus]          temp_b3_3_23_i;
wire signed [`CalcTempBus]          temp_b3_3_24_r;
wire signed [`CalcTempBus]          temp_b3_3_24_i;
wire signed [`CalcTempBus]          temp_b3_3_25_r;
wire signed [`CalcTempBus]          temp_b3_3_25_i;
wire signed [`CalcTempBus]          temp_b3_3_26_r;
wire signed [`CalcTempBus]          temp_b3_3_26_i;
wire signed [`CalcTempBus]          temp_b3_3_27_r;
wire signed [`CalcTempBus]          temp_b3_3_27_i;
wire signed [`CalcTempBus]          temp_b3_3_28_r;
wire signed [`CalcTempBus]          temp_b3_3_28_i;
wire signed [`CalcTempBus]          temp_b3_3_29_r;
wire signed [`CalcTempBus]          temp_b3_3_29_i;
wire signed [`CalcTempBus]          temp_b3_3_30_r;
wire signed [`CalcTempBus]          temp_b3_3_30_i;
wire signed [`CalcTempBus]          temp_b3_3_31_r;
wire signed [`CalcTempBus]          temp_b3_3_31_i;
wire signed [`CalcTempBus]          temp_b3_3_32_r;
wire signed [`CalcTempBus]          temp_b3_3_32_i;
wire signed [`CalcTempBus]          temp_b3_4_1_r;
wire signed [`CalcTempBus]          temp_b3_4_1_i;
wire signed [`CalcTempBus]          temp_b3_4_2_r;
wire signed [`CalcTempBus]          temp_b3_4_2_i;
wire signed [`CalcTempBus]          temp_b3_4_3_r;
wire signed [`CalcTempBus]          temp_b3_4_3_i;
wire signed [`CalcTempBus]          temp_b3_4_4_r;
wire signed [`CalcTempBus]          temp_b3_4_4_i;
wire signed [`CalcTempBus]          temp_b3_4_5_r;
wire signed [`CalcTempBus]          temp_b3_4_5_i;
wire signed [`CalcTempBus]          temp_b3_4_6_r;
wire signed [`CalcTempBus]          temp_b3_4_6_i;
wire signed [`CalcTempBus]          temp_b3_4_7_r;
wire signed [`CalcTempBus]          temp_b3_4_7_i;
wire signed [`CalcTempBus]          temp_b3_4_8_r;
wire signed [`CalcTempBus]          temp_b3_4_8_i;
wire signed [`CalcTempBus]          temp_b3_4_9_r;
wire signed [`CalcTempBus]          temp_b3_4_9_i;
wire signed [`CalcTempBus]          temp_b3_4_10_r;
wire signed [`CalcTempBus]          temp_b3_4_10_i;
wire signed [`CalcTempBus]          temp_b3_4_11_r;
wire signed [`CalcTempBus]          temp_b3_4_11_i;
wire signed [`CalcTempBus]          temp_b3_4_12_r;
wire signed [`CalcTempBus]          temp_b3_4_12_i;
wire signed [`CalcTempBus]          temp_b3_4_13_r;
wire signed [`CalcTempBus]          temp_b3_4_13_i;
wire signed [`CalcTempBus]          temp_b3_4_14_r;
wire signed [`CalcTempBus]          temp_b3_4_14_i;
wire signed [`CalcTempBus]          temp_b3_4_15_r;
wire signed [`CalcTempBus]          temp_b3_4_15_i;
wire signed [`CalcTempBus]          temp_b3_4_16_r;
wire signed [`CalcTempBus]          temp_b3_4_16_i;
wire signed [`CalcTempBus]          temp_b3_4_17_r;
wire signed [`CalcTempBus]          temp_b3_4_17_i;
wire signed [`CalcTempBus]          temp_b3_4_18_r;
wire signed [`CalcTempBus]          temp_b3_4_18_i;
wire signed [`CalcTempBus]          temp_b3_4_19_r;
wire signed [`CalcTempBus]          temp_b3_4_19_i;
wire signed [`CalcTempBus]          temp_b3_4_20_r;
wire signed [`CalcTempBus]          temp_b3_4_20_i;
wire signed [`CalcTempBus]          temp_b3_4_21_r;
wire signed [`CalcTempBus]          temp_b3_4_21_i;
wire signed [`CalcTempBus]          temp_b3_4_22_r;
wire signed [`CalcTempBus]          temp_b3_4_22_i;
wire signed [`CalcTempBus]          temp_b3_4_23_r;
wire signed [`CalcTempBus]          temp_b3_4_23_i;
wire signed [`CalcTempBus]          temp_b3_4_24_r;
wire signed [`CalcTempBus]          temp_b3_4_24_i;
wire signed [`CalcTempBus]          temp_b3_4_25_r;
wire signed [`CalcTempBus]          temp_b3_4_25_i;
wire signed [`CalcTempBus]          temp_b3_4_26_r;
wire signed [`CalcTempBus]          temp_b3_4_26_i;
wire signed [`CalcTempBus]          temp_b3_4_27_r;
wire signed [`CalcTempBus]          temp_b3_4_27_i;
wire signed [`CalcTempBus]          temp_b3_4_28_r;
wire signed [`CalcTempBus]          temp_b3_4_28_i;
wire signed [`CalcTempBus]          temp_b3_4_29_r;
wire signed [`CalcTempBus]          temp_b3_4_29_i;
wire signed [`CalcTempBus]          temp_b3_4_30_r;
wire signed [`CalcTempBus]          temp_b3_4_30_i;
wire signed [`CalcTempBus]          temp_b3_4_31_r;
wire signed [`CalcTempBus]          temp_b3_4_31_i;
wire signed [`CalcTempBus]          temp_b3_4_32_r;
wire signed [`CalcTempBus]          temp_b3_4_32_i;
wire signed [`CalcTempBus]          temp_b3_5_1_r;
wire signed [`CalcTempBus]          temp_b3_5_1_i;
wire signed [`CalcTempBus]          temp_b3_5_2_r;
wire signed [`CalcTempBus]          temp_b3_5_2_i;
wire signed [`CalcTempBus]          temp_b3_5_3_r;
wire signed [`CalcTempBus]          temp_b3_5_3_i;
wire signed [`CalcTempBus]          temp_b3_5_4_r;
wire signed [`CalcTempBus]          temp_b3_5_4_i;
wire signed [`CalcTempBus]          temp_b3_5_5_r;
wire signed [`CalcTempBus]          temp_b3_5_5_i;
wire signed [`CalcTempBus]          temp_b3_5_6_r;
wire signed [`CalcTempBus]          temp_b3_5_6_i;
wire signed [`CalcTempBus]          temp_b3_5_7_r;
wire signed [`CalcTempBus]          temp_b3_5_7_i;
wire signed [`CalcTempBus]          temp_b3_5_8_r;
wire signed [`CalcTempBus]          temp_b3_5_8_i;
wire signed [`CalcTempBus]          temp_b3_5_9_r;
wire signed [`CalcTempBus]          temp_b3_5_9_i;
wire signed [`CalcTempBus]          temp_b3_5_10_r;
wire signed [`CalcTempBus]          temp_b3_5_10_i;
wire signed [`CalcTempBus]          temp_b3_5_11_r;
wire signed [`CalcTempBus]          temp_b3_5_11_i;
wire signed [`CalcTempBus]          temp_b3_5_12_r;
wire signed [`CalcTempBus]          temp_b3_5_12_i;
wire signed [`CalcTempBus]          temp_b3_5_13_r;
wire signed [`CalcTempBus]          temp_b3_5_13_i;
wire signed [`CalcTempBus]          temp_b3_5_14_r;
wire signed [`CalcTempBus]          temp_b3_5_14_i;
wire signed [`CalcTempBus]          temp_b3_5_15_r;
wire signed [`CalcTempBus]          temp_b3_5_15_i;
wire signed [`CalcTempBus]          temp_b3_5_16_r;
wire signed [`CalcTempBus]          temp_b3_5_16_i;
wire signed [`CalcTempBus]          temp_b3_5_17_r;
wire signed [`CalcTempBus]          temp_b3_5_17_i;
wire signed [`CalcTempBus]          temp_b3_5_18_r;
wire signed [`CalcTempBus]          temp_b3_5_18_i;
wire signed [`CalcTempBus]          temp_b3_5_19_r;
wire signed [`CalcTempBus]          temp_b3_5_19_i;
wire signed [`CalcTempBus]          temp_b3_5_20_r;
wire signed [`CalcTempBus]          temp_b3_5_20_i;
wire signed [`CalcTempBus]          temp_b3_5_21_r;
wire signed [`CalcTempBus]          temp_b3_5_21_i;
wire signed [`CalcTempBus]          temp_b3_5_22_r;
wire signed [`CalcTempBus]          temp_b3_5_22_i;
wire signed [`CalcTempBus]          temp_b3_5_23_r;
wire signed [`CalcTempBus]          temp_b3_5_23_i;
wire signed [`CalcTempBus]          temp_b3_5_24_r;
wire signed [`CalcTempBus]          temp_b3_5_24_i;
wire signed [`CalcTempBus]          temp_b3_5_25_r;
wire signed [`CalcTempBus]          temp_b3_5_25_i;
wire signed [`CalcTempBus]          temp_b3_5_26_r;
wire signed [`CalcTempBus]          temp_b3_5_26_i;
wire signed [`CalcTempBus]          temp_b3_5_27_r;
wire signed [`CalcTempBus]          temp_b3_5_27_i;
wire signed [`CalcTempBus]          temp_b3_5_28_r;
wire signed [`CalcTempBus]          temp_b3_5_28_i;
wire signed [`CalcTempBus]          temp_b3_5_29_r;
wire signed [`CalcTempBus]          temp_b3_5_29_i;
wire signed [`CalcTempBus]          temp_b3_5_30_r;
wire signed [`CalcTempBus]          temp_b3_5_30_i;
wire signed [`CalcTempBus]          temp_b3_5_31_r;
wire signed [`CalcTempBus]          temp_b3_5_31_i;
wire signed [`CalcTempBus]          temp_b3_5_32_r;
wire signed [`CalcTempBus]          temp_b3_5_32_i;
wire signed [`CalcTempBus]          temp_b3_6_1_r;
wire signed [`CalcTempBus]          temp_b3_6_1_i;
wire signed [`CalcTempBus]          temp_b3_6_2_r;
wire signed [`CalcTempBus]          temp_b3_6_2_i;
wire signed [`CalcTempBus]          temp_b3_6_3_r;
wire signed [`CalcTempBus]          temp_b3_6_3_i;
wire signed [`CalcTempBus]          temp_b3_6_4_r;
wire signed [`CalcTempBus]          temp_b3_6_4_i;
wire signed [`CalcTempBus]          temp_b3_6_5_r;
wire signed [`CalcTempBus]          temp_b3_6_5_i;
wire signed [`CalcTempBus]          temp_b3_6_6_r;
wire signed [`CalcTempBus]          temp_b3_6_6_i;
wire signed [`CalcTempBus]          temp_b3_6_7_r;
wire signed [`CalcTempBus]          temp_b3_6_7_i;
wire signed [`CalcTempBus]          temp_b3_6_8_r;
wire signed [`CalcTempBus]          temp_b3_6_8_i;
wire signed [`CalcTempBus]          temp_b3_6_9_r;
wire signed [`CalcTempBus]          temp_b3_6_9_i;
wire signed [`CalcTempBus]          temp_b3_6_10_r;
wire signed [`CalcTempBus]          temp_b3_6_10_i;
wire signed [`CalcTempBus]          temp_b3_6_11_r;
wire signed [`CalcTempBus]          temp_b3_6_11_i;
wire signed [`CalcTempBus]          temp_b3_6_12_r;
wire signed [`CalcTempBus]          temp_b3_6_12_i;
wire signed [`CalcTempBus]          temp_b3_6_13_r;
wire signed [`CalcTempBus]          temp_b3_6_13_i;
wire signed [`CalcTempBus]          temp_b3_6_14_r;
wire signed [`CalcTempBus]          temp_b3_6_14_i;
wire signed [`CalcTempBus]          temp_b3_6_15_r;
wire signed [`CalcTempBus]          temp_b3_6_15_i;
wire signed [`CalcTempBus]          temp_b3_6_16_r;
wire signed [`CalcTempBus]          temp_b3_6_16_i;
wire signed [`CalcTempBus]          temp_b3_6_17_r;
wire signed [`CalcTempBus]          temp_b3_6_17_i;
wire signed [`CalcTempBus]          temp_b3_6_18_r;
wire signed [`CalcTempBus]          temp_b3_6_18_i;
wire signed [`CalcTempBus]          temp_b3_6_19_r;
wire signed [`CalcTempBus]          temp_b3_6_19_i;
wire signed [`CalcTempBus]          temp_b3_6_20_r;
wire signed [`CalcTempBus]          temp_b3_6_20_i;
wire signed [`CalcTempBus]          temp_b3_6_21_r;
wire signed [`CalcTempBus]          temp_b3_6_21_i;
wire signed [`CalcTempBus]          temp_b3_6_22_r;
wire signed [`CalcTempBus]          temp_b3_6_22_i;
wire signed [`CalcTempBus]          temp_b3_6_23_r;
wire signed [`CalcTempBus]          temp_b3_6_23_i;
wire signed [`CalcTempBus]          temp_b3_6_24_r;
wire signed [`CalcTempBus]          temp_b3_6_24_i;
wire signed [`CalcTempBus]          temp_b3_6_25_r;
wire signed [`CalcTempBus]          temp_b3_6_25_i;
wire signed [`CalcTempBus]          temp_b3_6_26_r;
wire signed [`CalcTempBus]          temp_b3_6_26_i;
wire signed [`CalcTempBus]          temp_b3_6_27_r;
wire signed [`CalcTempBus]          temp_b3_6_27_i;
wire signed [`CalcTempBus]          temp_b3_6_28_r;
wire signed [`CalcTempBus]          temp_b3_6_28_i;
wire signed [`CalcTempBus]          temp_b3_6_29_r;
wire signed [`CalcTempBus]          temp_b3_6_29_i;
wire signed [`CalcTempBus]          temp_b3_6_30_r;
wire signed [`CalcTempBus]          temp_b3_6_30_i;
wire signed [`CalcTempBus]          temp_b3_6_31_r;
wire signed [`CalcTempBus]          temp_b3_6_31_i;
wire signed [`CalcTempBus]          temp_b3_6_32_r;
wire signed [`CalcTempBus]          temp_b3_6_32_i;
wire signed [`CalcTempBus]          temp_b3_7_1_r;
wire signed [`CalcTempBus]          temp_b3_7_1_i;
wire signed [`CalcTempBus]          temp_b3_7_2_r;
wire signed [`CalcTempBus]          temp_b3_7_2_i;
wire signed [`CalcTempBus]          temp_b3_7_3_r;
wire signed [`CalcTempBus]          temp_b3_7_3_i;
wire signed [`CalcTempBus]          temp_b3_7_4_r;
wire signed [`CalcTempBus]          temp_b3_7_4_i;
wire signed [`CalcTempBus]          temp_b3_7_5_r;
wire signed [`CalcTempBus]          temp_b3_7_5_i;
wire signed [`CalcTempBus]          temp_b3_7_6_r;
wire signed [`CalcTempBus]          temp_b3_7_6_i;
wire signed [`CalcTempBus]          temp_b3_7_7_r;
wire signed [`CalcTempBus]          temp_b3_7_7_i;
wire signed [`CalcTempBus]          temp_b3_7_8_r;
wire signed [`CalcTempBus]          temp_b3_7_8_i;
wire signed [`CalcTempBus]          temp_b3_7_9_r;
wire signed [`CalcTempBus]          temp_b3_7_9_i;
wire signed [`CalcTempBus]          temp_b3_7_10_r;
wire signed [`CalcTempBus]          temp_b3_7_10_i;
wire signed [`CalcTempBus]          temp_b3_7_11_r;
wire signed [`CalcTempBus]          temp_b3_7_11_i;
wire signed [`CalcTempBus]          temp_b3_7_12_r;
wire signed [`CalcTempBus]          temp_b3_7_12_i;
wire signed [`CalcTempBus]          temp_b3_7_13_r;
wire signed [`CalcTempBus]          temp_b3_7_13_i;
wire signed [`CalcTempBus]          temp_b3_7_14_r;
wire signed [`CalcTempBus]          temp_b3_7_14_i;
wire signed [`CalcTempBus]          temp_b3_7_15_r;
wire signed [`CalcTempBus]          temp_b3_7_15_i;
wire signed [`CalcTempBus]          temp_b3_7_16_r;
wire signed [`CalcTempBus]          temp_b3_7_16_i;
wire signed [`CalcTempBus]          temp_b3_7_17_r;
wire signed [`CalcTempBus]          temp_b3_7_17_i;
wire signed [`CalcTempBus]          temp_b3_7_18_r;
wire signed [`CalcTempBus]          temp_b3_7_18_i;
wire signed [`CalcTempBus]          temp_b3_7_19_r;
wire signed [`CalcTempBus]          temp_b3_7_19_i;
wire signed [`CalcTempBus]          temp_b3_7_20_r;
wire signed [`CalcTempBus]          temp_b3_7_20_i;
wire signed [`CalcTempBus]          temp_b3_7_21_r;
wire signed [`CalcTempBus]          temp_b3_7_21_i;
wire signed [`CalcTempBus]          temp_b3_7_22_r;
wire signed [`CalcTempBus]          temp_b3_7_22_i;
wire signed [`CalcTempBus]          temp_b3_7_23_r;
wire signed [`CalcTempBus]          temp_b3_7_23_i;
wire signed [`CalcTempBus]          temp_b3_7_24_r;
wire signed [`CalcTempBus]          temp_b3_7_24_i;
wire signed [`CalcTempBus]          temp_b3_7_25_r;
wire signed [`CalcTempBus]          temp_b3_7_25_i;
wire signed [`CalcTempBus]          temp_b3_7_26_r;
wire signed [`CalcTempBus]          temp_b3_7_26_i;
wire signed [`CalcTempBus]          temp_b3_7_27_r;
wire signed [`CalcTempBus]          temp_b3_7_27_i;
wire signed [`CalcTempBus]          temp_b3_7_28_r;
wire signed [`CalcTempBus]          temp_b3_7_28_i;
wire signed [`CalcTempBus]          temp_b3_7_29_r;
wire signed [`CalcTempBus]          temp_b3_7_29_i;
wire signed [`CalcTempBus]          temp_b3_7_30_r;
wire signed [`CalcTempBus]          temp_b3_7_30_i;
wire signed [`CalcTempBus]          temp_b3_7_31_r;
wire signed [`CalcTempBus]          temp_b3_7_31_i;
wire signed [`CalcTempBus]          temp_b3_7_32_r;
wire signed [`CalcTempBus]          temp_b3_7_32_i;
wire signed [`CalcTempBus]          temp_b3_8_1_r;
wire signed [`CalcTempBus]          temp_b3_8_1_i;
wire signed [`CalcTempBus]          temp_b3_8_2_r;
wire signed [`CalcTempBus]          temp_b3_8_2_i;
wire signed [`CalcTempBus]          temp_b3_8_3_r;
wire signed [`CalcTempBus]          temp_b3_8_3_i;
wire signed [`CalcTempBus]          temp_b3_8_4_r;
wire signed [`CalcTempBus]          temp_b3_8_4_i;
wire signed [`CalcTempBus]          temp_b3_8_5_r;
wire signed [`CalcTempBus]          temp_b3_8_5_i;
wire signed [`CalcTempBus]          temp_b3_8_6_r;
wire signed [`CalcTempBus]          temp_b3_8_6_i;
wire signed [`CalcTempBus]          temp_b3_8_7_r;
wire signed [`CalcTempBus]          temp_b3_8_7_i;
wire signed [`CalcTempBus]          temp_b3_8_8_r;
wire signed [`CalcTempBus]          temp_b3_8_8_i;
wire signed [`CalcTempBus]          temp_b3_8_9_r;
wire signed [`CalcTempBus]          temp_b3_8_9_i;
wire signed [`CalcTempBus]          temp_b3_8_10_r;
wire signed [`CalcTempBus]          temp_b3_8_10_i;
wire signed [`CalcTempBus]          temp_b3_8_11_r;
wire signed [`CalcTempBus]          temp_b3_8_11_i;
wire signed [`CalcTempBus]          temp_b3_8_12_r;
wire signed [`CalcTempBus]          temp_b3_8_12_i;
wire signed [`CalcTempBus]          temp_b3_8_13_r;
wire signed [`CalcTempBus]          temp_b3_8_13_i;
wire signed [`CalcTempBus]          temp_b3_8_14_r;
wire signed [`CalcTempBus]          temp_b3_8_14_i;
wire signed [`CalcTempBus]          temp_b3_8_15_r;
wire signed [`CalcTempBus]          temp_b3_8_15_i;
wire signed [`CalcTempBus]          temp_b3_8_16_r;
wire signed [`CalcTempBus]          temp_b3_8_16_i;
wire signed [`CalcTempBus]          temp_b3_8_17_r;
wire signed [`CalcTempBus]          temp_b3_8_17_i;
wire signed [`CalcTempBus]          temp_b3_8_18_r;
wire signed [`CalcTempBus]          temp_b3_8_18_i;
wire signed [`CalcTempBus]          temp_b3_8_19_r;
wire signed [`CalcTempBus]          temp_b3_8_19_i;
wire signed [`CalcTempBus]          temp_b3_8_20_r;
wire signed [`CalcTempBus]          temp_b3_8_20_i;
wire signed [`CalcTempBus]          temp_b3_8_21_r;
wire signed [`CalcTempBus]          temp_b3_8_21_i;
wire signed [`CalcTempBus]          temp_b3_8_22_r;
wire signed [`CalcTempBus]          temp_b3_8_22_i;
wire signed [`CalcTempBus]          temp_b3_8_23_r;
wire signed [`CalcTempBus]          temp_b3_8_23_i;
wire signed [`CalcTempBus]          temp_b3_8_24_r;
wire signed [`CalcTempBus]          temp_b3_8_24_i;
wire signed [`CalcTempBus]          temp_b3_8_25_r;
wire signed [`CalcTempBus]          temp_b3_8_25_i;
wire signed [`CalcTempBus]          temp_b3_8_26_r;
wire signed [`CalcTempBus]          temp_b3_8_26_i;
wire signed [`CalcTempBus]          temp_b3_8_27_r;
wire signed [`CalcTempBus]          temp_b3_8_27_i;
wire signed [`CalcTempBus]          temp_b3_8_28_r;
wire signed [`CalcTempBus]          temp_b3_8_28_i;
wire signed [`CalcTempBus]          temp_b3_8_29_r;
wire signed [`CalcTempBus]          temp_b3_8_29_i;
wire signed [`CalcTempBus]          temp_b3_8_30_r;
wire signed [`CalcTempBus]          temp_b3_8_30_i;
wire signed [`CalcTempBus]          temp_b3_8_31_r;
wire signed [`CalcTempBus]          temp_b3_8_31_i;
wire signed [`CalcTempBus]          temp_b3_8_32_r;
wire signed [`CalcTempBus]          temp_b3_8_32_i;
wire signed [`CalcTempBus]          temp_b3_9_1_r;
wire signed [`CalcTempBus]          temp_b3_9_1_i;
wire signed [`CalcTempBus]          temp_b3_9_2_r;
wire signed [`CalcTempBus]          temp_b3_9_2_i;
wire signed [`CalcTempBus]          temp_b3_9_3_r;
wire signed [`CalcTempBus]          temp_b3_9_3_i;
wire signed [`CalcTempBus]          temp_b3_9_4_r;
wire signed [`CalcTempBus]          temp_b3_9_4_i;
wire signed [`CalcTempBus]          temp_b3_9_5_r;
wire signed [`CalcTempBus]          temp_b3_9_5_i;
wire signed [`CalcTempBus]          temp_b3_9_6_r;
wire signed [`CalcTempBus]          temp_b3_9_6_i;
wire signed [`CalcTempBus]          temp_b3_9_7_r;
wire signed [`CalcTempBus]          temp_b3_9_7_i;
wire signed [`CalcTempBus]          temp_b3_9_8_r;
wire signed [`CalcTempBus]          temp_b3_9_8_i;
wire signed [`CalcTempBus]          temp_b3_9_9_r;
wire signed [`CalcTempBus]          temp_b3_9_9_i;
wire signed [`CalcTempBus]          temp_b3_9_10_r;
wire signed [`CalcTempBus]          temp_b3_9_10_i;
wire signed [`CalcTempBus]          temp_b3_9_11_r;
wire signed [`CalcTempBus]          temp_b3_9_11_i;
wire signed [`CalcTempBus]          temp_b3_9_12_r;
wire signed [`CalcTempBus]          temp_b3_9_12_i;
wire signed [`CalcTempBus]          temp_b3_9_13_r;
wire signed [`CalcTempBus]          temp_b3_9_13_i;
wire signed [`CalcTempBus]          temp_b3_9_14_r;
wire signed [`CalcTempBus]          temp_b3_9_14_i;
wire signed [`CalcTempBus]          temp_b3_9_15_r;
wire signed [`CalcTempBus]          temp_b3_9_15_i;
wire signed [`CalcTempBus]          temp_b3_9_16_r;
wire signed [`CalcTempBus]          temp_b3_9_16_i;
wire signed [`CalcTempBus]          temp_b3_9_17_r;
wire signed [`CalcTempBus]          temp_b3_9_17_i;
wire signed [`CalcTempBus]          temp_b3_9_18_r;
wire signed [`CalcTempBus]          temp_b3_9_18_i;
wire signed [`CalcTempBus]          temp_b3_9_19_r;
wire signed [`CalcTempBus]          temp_b3_9_19_i;
wire signed [`CalcTempBus]          temp_b3_9_20_r;
wire signed [`CalcTempBus]          temp_b3_9_20_i;
wire signed [`CalcTempBus]          temp_b3_9_21_r;
wire signed [`CalcTempBus]          temp_b3_9_21_i;
wire signed [`CalcTempBus]          temp_b3_9_22_r;
wire signed [`CalcTempBus]          temp_b3_9_22_i;
wire signed [`CalcTempBus]          temp_b3_9_23_r;
wire signed [`CalcTempBus]          temp_b3_9_23_i;
wire signed [`CalcTempBus]          temp_b3_9_24_r;
wire signed [`CalcTempBus]          temp_b3_9_24_i;
wire signed [`CalcTempBus]          temp_b3_9_25_r;
wire signed [`CalcTempBus]          temp_b3_9_25_i;
wire signed [`CalcTempBus]          temp_b3_9_26_r;
wire signed [`CalcTempBus]          temp_b3_9_26_i;
wire signed [`CalcTempBus]          temp_b3_9_27_r;
wire signed [`CalcTempBus]          temp_b3_9_27_i;
wire signed [`CalcTempBus]          temp_b3_9_28_r;
wire signed [`CalcTempBus]          temp_b3_9_28_i;
wire signed [`CalcTempBus]          temp_b3_9_29_r;
wire signed [`CalcTempBus]          temp_b3_9_29_i;
wire signed [`CalcTempBus]          temp_b3_9_30_r;
wire signed [`CalcTempBus]          temp_b3_9_30_i;
wire signed [`CalcTempBus]          temp_b3_9_31_r;
wire signed [`CalcTempBus]          temp_b3_9_31_i;
wire signed [`CalcTempBus]          temp_b3_9_32_r;
wire signed [`CalcTempBus]          temp_b3_9_32_i;
wire signed [`CalcTempBus]          temp_b3_10_1_r;
wire signed [`CalcTempBus]          temp_b3_10_1_i;
wire signed [`CalcTempBus]          temp_b3_10_2_r;
wire signed [`CalcTempBus]          temp_b3_10_2_i;
wire signed [`CalcTempBus]          temp_b3_10_3_r;
wire signed [`CalcTempBus]          temp_b3_10_3_i;
wire signed [`CalcTempBus]          temp_b3_10_4_r;
wire signed [`CalcTempBus]          temp_b3_10_4_i;
wire signed [`CalcTempBus]          temp_b3_10_5_r;
wire signed [`CalcTempBus]          temp_b3_10_5_i;
wire signed [`CalcTempBus]          temp_b3_10_6_r;
wire signed [`CalcTempBus]          temp_b3_10_6_i;
wire signed [`CalcTempBus]          temp_b3_10_7_r;
wire signed [`CalcTempBus]          temp_b3_10_7_i;
wire signed [`CalcTempBus]          temp_b3_10_8_r;
wire signed [`CalcTempBus]          temp_b3_10_8_i;
wire signed [`CalcTempBus]          temp_b3_10_9_r;
wire signed [`CalcTempBus]          temp_b3_10_9_i;
wire signed [`CalcTempBus]          temp_b3_10_10_r;
wire signed [`CalcTempBus]          temp_b3_10_10_i;
wire signed [`CalcTempBus]          temp_b3_10_11_r;
wire signed [`CalcTempBus]          temp_b3_10_11_i;
wire signed [`CalcTempBus]          temp_b3_10_12_r;
wire signed [`CalcTempBus]          temp_b3_10_12_i;
wire signed [`CalcTempBus]          temp_b3_10_13_r;
wire signed [`CalcTempBus]          temp_b3_10_13_i;
wire signed [`CalcTempBus]          temp_b3_10_14_r;
wire signed [`CalcTempBus]          temp_b3_10_14_i;
wire signed [`CalcTempBus]          temp_b3_10_15_r;
wire signed [`CalcTempBus]          temp_b3_10_15_i;
wire signed [`CalcTempBus]          temp_b3_10_16_r;
wire signed [`CalcTempBus]          temp_b3_10_16_i;
wire signed [`CalcTempBus]          temp_b3_10_17_r;
wire signed [`CalcTempBus]          temp_b3_10_17_i;
wire signed [`CalcTempBus]          temp_b3_10_18_r;
wire signed [`CalcTempBus]          temp_b3_10_18_i;
wire signed [`CalcTempBus]          temp_b3_10_19_r;
wire signed [`CalcTempBus]          temp_b3_10_19_i;
wire signed [`CalcTempBus]          temp_b3_10_20_r;
wire signed [`CalcTempBus]          temp_b3_10_20_i;
wire signed [`CalcTempBus]          temp_b3_10_21_r;
wire signed [`CalcTempBus]          temp_b3_10_21_i;
wire signed [`CalcTempBus]          temp_b3_10_22_r;
wire signed [`CalcTempBus]          temp_b3_10_22_i;
wire signed [`CalcTempBus]          temp_b3_10_23_r;
wire signed [`CalcTempBus]          temp_b3_10_23_i;
wire signed [`CalcTempBus]          temp_b3_10_24_r;
wire signed [`CalcTempBus]          temp_b3_10_24_i;
wire signed [`CalcTempBus]          temp_b3_10_25_r;
wire signed [`CalcTempBus]          temp_b3_10_25_i;
wire signed [`CalcTempBus]          temp_b3_10_26_r;
wire signed [`CalcTempBus]          temp_b3_10_26_i;
wire signed [`CalcTempBus]          temp_b3_10_27_r;
wire signed [`CalcTempBus]          temp_b3_10_27_i;
wire signed [`CalcTempBus]          temp_b3_10_28_r;
wire signed [`CalcTempBus]          temp_b3_10_28_i;
wire signed [`CalcTempBus]          temp_b3_10_29_r;
wire signed [`CalcTempBus]          temp_b3_10_29_i;
wire signed [`CalcTempBus]          temp_b3_10_30_r;
wire signed [`CalcTempBus]          temp_b3_10_30_i;
wire signed [`CalcTempBus]          temp_b3_10_31_r;
wire signed [`CalcTempBus]          temp_b3_10_31_i;
wire signed [`CalcTempBus]          temp_b3_10_32_r;
wire signed [`CalcTempBus]          temp_b3_10_32_i;
wire signed [`CalcTempBus]          temp_b3_11_1_r;
wire signed [`CalcTempBus]          temp_b3_11_1_i;
wire signed [`CalcTempBus]          temp_b3_11_2_r;
wire signed [`CalcTempBus]          temp_b3_11_2_i;
wire signed [`CalcTempBus]          temp_b3_11_3_r;
wire signed [`CalcTempBus]          temp_b3_11_3_i;
wire signed [`CalcTempBus]          temp_b3_11_4_r;
wire signed [`CalcTempBus]          temp_b3_11_4_i;
wire signed [`CalcTempBus]          temp_b3_11_5_r;
wire signed [`CalcTempBus]          temp_b3_11_5_i;
wire signed [`CalcTempBus]          temp_b3_11_6_r;
wire signed [`CalcTempBus]          temp_b3_11_6_i;
wire signed [`CalcTempBus]          temp_b3_11_7_r;
wire signed [`CalcTempBus]          temp_b3_11_7_i;
wire signed [`CalcTempBus]          temp_b3_11_8_r;
wire signed [`CalcTempBus]          temp_b3_11_8_i;
wire signed [`CalcTempBus]          temp_b3_11_9_r;
wire signed [`CalcTempBus]          temp_b3_11_9_i;
wire signed [`CalcTempBus]          temp_b3_11_10_r;
wire signed [`CalcTempBus]          temp_b3_11_10_i;
wire signed [`CalcTempBus]          temp_b3_11_11_r;
wire signed [`CalcTempBus]          temp_b3_11_11_i;
wire signed [`CalcTempBus]          temp_b3_11_12_r;
wire signed [`CalcTempBus]          temp_b3_11_12_i;
wire signed [`CalcTempBus]          temp_b3_11_13_r;
wire signed [`CalcTempBus]          temp_b3_11_13_i;
wire signed [`CalcTempBus]          temp_b3_11_14_r;
wire signed [`CalcTempBus]          temp_b3_11_14_i;
wire signed [`CalcTempBus]          temp_b3_11_15_r;
wire signed [`CalcTempBus]          temp_b3_11_15_i;
wire signed [`CalcTempBus]          temp_b3_11_16_r;
wire signed [`CalcTempBus]          temp_b3_11_16_i;
wire signed [`CalcTempBus]          temp_b3_11_17_r;
wire signed [`CalcTempBus]          temp_b3_11_17_i;
wire signed [`CalcTempBus]          temp_b3_11_18_r;
wire signed [`CalcTempBus]          temp_b3_11_18_i;
wire signed [`CalcTempBus]          temp_b3_11_19_r;
wire signed [`CalcTempBus]          temp_b3_11_19_i;
wire signed [`CalcTempBus]          temp_b3_11_20_r;
wire signed [`CalcTempBus]          temp_b3_11_20_i;
wire signed [`CalcTempBus]          temp_b3_11_21_r;
wire signed [`CalcTempBus]          temp_b3_11_21_i;
wire signed [`CalcTempBus]          temp_b3_11_22_r;
wire signed [`CalcTempBus]          temp_b3_11_22_i;
wire signed [`CalcTempBus]          temp_b3_11_23_r;
wire signed [`CalcTempBus]          temp_b3_11_23_i;
wire signed [`CalcTempBus]          temp_b3_11_24_r;
wire signed [`CalcTempBus]          temp_b3_11_24_i;
wire signed [`CalcTempBus]          temp_b3_11_25_r;
wire signed [`CalcTempBus]          temp_b3_11_25_i;
wire signed [`CalcTempBus]          temp_b3_11_26_r;
wire signed [`CalcTempBus]          temp_b3_11_26_i;
wire signed [`CalcTempBus]          temp_b3_11_27_r;
wire signed [`CalcTempBus]          temp_b3_11_27_i;
wire signed [`CalcTempBus]          temp_b3_11_28_r;
wire signed [`CalcTempBus]          temp_b3_11_28_i;
wire signed [`CalcTempBus]          temp_b3_11_29_r;
wire signed [`CalcTempBus]          temp_b3_11_29_i;
wire signed [`CalcTempBus]          temp_b3_11_30_r;
wire signed [`CalcTempBus]          temp_b3_11_30_i;
wire signed [`CalcTempBus]          temp_b3_11_31_r;
wire signed [`CalcTempBus]          temp_b3_11_31_i;
wire signed [`CalcTempBus]          temp_b3_11_32_r;
wire signed [`CalcTempBus]          temp_b3_11_32_i;
wire signed [`CalcTempBus]          temp_b3_12_1_r;
wire signed [`CalcTempBus]          temp_b3_12_1_i;
wire signed [`CalcTempBus]          temp_b3_12_2_r;
wire signed [`CalcTempBus]          temp_b3_12_2_i;
wire signed [`CalcTempBus]          temp_b3_12_3_r;
wire signed [`CalcTempBus]          temp_b3_12_3_i;
wire signed [`CalcTempBus]          temp_b3_12_4_r;
wire signed [`CalcTempBus]          temp_b3_12_4_i;
wire signed [`CalcTempBus]          temp_b3_12_5_r;
wire signed [`CalcTempBus]          temp_b3_12_5_i;
wire signed [`CalcTempBus]          temp_b3_12_6_r;
wire signed [`CalcTempBus]          temp_b3_12_6_i;
wire signed [`CalcTempBus]          temp_b3_12_7_r;
wire signed [`CalcTempBus]          temp_b3_12_7_i;
wire signed [`CalcTempBus]          temp_b3_12_8_r;
wire signed [`CalcTempBus]          temp_b3_12_8_i;
wire signed [`CalcTempBus]          temp_b3_12_9_r;
wire signed [`CalcTempBus]          temp_b3_12_9_i;
wire signed [`CalcTempBus]          temp_b3_12_10_r;
wire signed [`CalcTempBus]          temp_b3_12_10_i;
wire signed [`CalcTempBus]          temp_b3_12_11_r;
wire signed [`CalcTempBus]          temp_b3_12_11_i;
wire signed [`CalcTempBus]          temp_b3_12_12_r;
wire signed [`CalcTempBus]          temp_b3_12_12_i;
wire signed [`CalcTempBus]          temp_b3_12_13_r;
wire signed [`CalcTempBus]          temp_b3_12_13_i;
wire signed [`CalcTempBus]          temp_b3_12_14_r;
wire signed [`CalcTempBus]          temp_b3_12_14_i;
wire signed [`CalcTempBus]          temp_b3_12_15_r;
wire signed [`CalcTempBus]          temp_b3_12_15_i;
wire signed [`CalcTempBus]          temp_b3_12_16_r;
wire signed [`CalcTempBus]          temp_b3_12_16_i;
wire signed [`CalcTempBus]          temp_b3_12_17_r;
wire signed [`CalcTempBus]          temp_b3_12_17_i;
wire signed [`CalcTempBus]          temp_b3_12_18_r;
wire signed [`CalcTempBus]          temp_b3_12_18_i;
wire signed [`CalcTempBus]          temp_b3_12_19_r;
wire signed [`CalcTempBus]          temp_b3_12_19_i;
wire signed [`CalcTempBus]          temp_b3_12_20_r;
wire signed [`CalcTempBus]          temp_b3_12_20_i;
wire signed [`CalcTempBus]          temp_b3_12_21_r;
wire signed [`CalcTempBus]          temp_b3_12_21_i;
wire signed [`CalcTempBus]          temp_b3_12_22_r;
wire signed [`CalcTempBus]          temp_b3_12_22_i;
wire signed [`CalcTempBus]          temp_b3_12_23_r;
wire signed [`CalcTempBus]          temp_b3_12_23_i;
wire signed [`CalcTempBus]          temp_b3_12_24_r;
wire signed [`CalcTempBus]          temp_b3_12_24_i;
wire signed [`CalcTempBus]          temp_b3_12_25_r;
wire signed [`CalcTempBus]          temp_b3_12_25_i;
wire signed [`CalcTempBus]          temp_b3_12_26_r;
wire signed [`CalcTempBus]          temp_b3_12_26_i;
wire signed [`CalcTempBus]          temp_b3_12_27_r;
wire signed [`CalcTempBus]          temp_b3_12_27_i;
wire signed [`CalcTempBus]          temp_b3_12_28_r;
wire signed [`CalcTempBus]          temp_b3_12_28_i;
wire signed [`CalcTempBus]          temp_b3_12_29_r;
wire signed [`CalcTempBus]          temp_b3_12_29_i;
wire signed [`CalcTempBus]          temp_b3_12_30_r;
wire signed [`CalcTempBus]          temp_b3_12_30_i;
wire signed [`CalcTempBus]          temp_b3_12_31_r;
wire signed [`CalcTempBus]          temp_b3_12_31_i;
wire signed [`CalcTempBus]          temp_b3_12_32_r;
wire signed [`CalcTempBus]          temp_b3_12_32_i;
wire signed [`CalcTempBus]          temp_b3_13_1_r;
wire signed [`CalcTempBus]          temp_b3_13_1_i;
wire signed [`CalcTempBus]          temp_b3_13_2_r;
wire signed [`CalcTempBus]          temp_b3_13_2_i;
wire signed [`CalcTempBus]          temp_b3_13_3_r;
wire signed [`CalcTempBus]          temp_b3_13_3_i;
wire signed [`CalcTempBus]          temp_b3_13_4_r;
wire signed [`CalcTempBus]          temp_b3_13_4_i;
wire signed [`CalcTempBus]          temp_b3_13_5_r;
wire signed [`CalcTempBus]          temp_b3_13_5_i;
wire signed [`CalcTempBus]          temp_b3_13_6_r;
wire signed [`CalcTempBus]          temp_b3_13_6_i;
wire signed [`CalcTempBus]          temp_b3_13_7_r;
wire signed [`CalcTempBus]          temp_b3_13_7_i;
wire signed [`CalcTempBus]          temp_b3_13_8_r;
wire signed [`CalcTempBus]          temp_b3_13_8_i;
wire signed [`CalcTempBus]          temp_b3_13_9_r;
wire signed [`CalcTempBus]          temp_b3_13_9_i;
wire signed [`CalcTempBus]          temp_b3_13_10_r;
wire signed [`CalcTempBus]          temp_b3_13_10_i;
wire signed [`CalcTempBus]          temp_b3_13_11_r;
wire signed [`CalcTempBus]          temp_b3_13_11_i;
wire signed [`CalcTempBus]          temp_b3_13_12_r;
wire signed [`CalcTempBus]          temp_b3_13_12_i;
wire signed [`CalcTempBus]          temp_b3_13_13_r;
wire signed [`CalcTempBus]          temp_b3_13_13_i;
wire signed [`CalcTempBus]          temp_b3_13_14_r;
wire signed [`CalcTempBus]          temp_b3_13_14_i;
wire signed [`CalcTempBus]          temp_b3_13_15_r;
wire signed [`CalcTempBus]          temp_b3_13_15_i;
wire signed [`CalcTempBus]          temp_b3_13_16_r;
wire signed [`CalcTempBus]          temp_b3_13_16_i;
wire signed [`CalcTempBus]          temp_b3_13_17_r;
wire signed [`CalcTempBus]          temp_b3_13_17_i;
wire signed [`CalcTempBus]          temp_b3_13_18_r;
wire signed [`CalcTempBus]          temp_b3_13_18_i;
wire signed [`CalcTempBus]          temp_b3_13_19_r;
wire signed [`CalcTempBus]          temp_b3_13_19_i;
wire signed [`CalcTempBus]          temp_b3_13_20_r;
wire signed [`CalcTempBus]          temp_b3_13_20_i;
wire signed [`CalcTempBus]          temp_b3_13_21_r;
wire signed [`CalcTempBus]          temp_b3_13_21_i;
wire signed [`CalcTempBus]          temp_b3_13_22_r;
wire signed [`CalcTempBus]          temp_b3_13_22_i;
wire signed [`CalcTempBus]          temp_b3_13_23_r;
wire signed [`CalcTempBus]          temp_b3_13_23_i;
wire signed [`CalcTempBus]          temp_b3_13_24_r;
wire signed [`CalcTempBus]          temp_b3_13_24_i;
wire signed [`CalcTempBus]          temp_b3_13_25_r;
wire signed [`CalcTempBus]          temp_b3_13_25_i;
wire signed [`CalcTempBus]          temp_b3_13_26_r;
wire signed [`CalcTempBus]          temp_b3_13_26_i;
wire signed [`CalcTempBus]          temp_b3_13_27_r;
wire signed [`CalcTempBus]          temp_b3_13_27_i;
wire signed [`CalcTempBus]          temp_b3_13_28_r;
wire signed [`CalcTempBus]          temp_b3_13_28_i;
wire signed [`CalcTempBus]          temp_b3_13_29_r;
wire signed [`CalcTempBus]          temp_b3_13_29_i;
wire signed [`CalcTempBus]          temp_b3_13_30_r;
wire signed [`CalcTempBus]          temp_b3_13_30_i;
wire signed [`CalcTempBus]          temp_b3_13_31_r;
wire signed [`CalcTempBus]          temp_b3_13_31_i;
wire signed [`CalcTempBus]          temp_b3_13_32_r;
wire signed [`CalcTempBus]          temp_b3_13_32_i;
wire signed [`CalcTempBus]          temp_b3_14_1_r;
wire signed [`CalcTempBus]          temp_b3_14_1_i;
wire signed [`CalcTempBus]          temp_b3_14_2_r;
wire signed [`CalcTempBus]          temp_b3_14_2_i;
wire signed [`CalcTempBus]          temp_b3_14_3_r;
wire signed [`CalcTempBus]          temp_b3_14_3_i;
wire signed [`CalcTempBus]          temp_b3_14_4_r;
wire signed [`CalcTempBus]          temp_b3_14_4_i;
wire signed [`CalcTempBus]          temp_b3_14_5_r;
wire signed [`CalcTempBus]          temp_b3_14_5_i;
wire signed [`CalcTempBus]          temp_b3_14_6_r;
wire signed [`CalcTempBus]          temp_b3_14_6_i;
wire signed [`CalcTempBus]          temp_b3_14_7_r;
wire signed [`CalcTempBus]          temp_b3_14_7_i;
wire signed [`CalcTempBus]          temp_b3_14_8_r;
wire signed [`CalcTempBus]          temp_b3_14_8_i;
wire signed [`CalcTempBus]          temp_b3_14_9_r;
wire signed [`CalcTempBus]          temp_b3_14_9_i;
wire signed [`CalcTempBus]          temp_b3_14_10_r;
wire signed [`CalcTempBus]          temp_b3_14_10_i;
wire signed [`CalcTempBus]          temp_b3_14_11_r;
wire signed [`CalcTempBus]          temp_b3_14_11_i;
wire signed [`CalcTempBus]          temp_b3_14_12_r;
wire signed [`CalcTempBus]          temp_b3_14_12_i;
wire signed [`CalcTempBus]          temp_b3_14_13_r;
wire signed [`CalcTempBus]          temp_b3_14_13_i;
wire signed [`CalcTempBus]          temp_b3_14_14_r;
wire signed [`CalcTempBus]          temp_b3_14_14_i;
wire signed [`CalcTempBus]          temp_b3_14_15_r;
wire signed [`CalcTempBus]          temp_b3_14_15_i;
wire signed [`CalcTempBus]          temp_b3_14_16_r;
wire signed [`CalcTempBus]          temp_b3_14_16_i;
wire signed [`CalcTempBus]          temp_b3_14_17_r;
wire signed [`CalcTempBus]          temp_b3_14_17_i;
wire signed [`CalcTempBus]          temp_b3_14_18_r;
wire signed [`CalcTempBus]          temp_b3_14_18_i;
wire signed [`CalcTempBus]          temp_b3_14_19_r;
wire signed [`CalcTempBus]          temp_b3_14_19_i;
wire signed [`CalcTempBus]          temp_b3_14_20_r;
wire signed [`CalcTempBus]          temp_b3_14_20_i;
wire signed [`CalcTempBus]          temp_b3_14_21_r;
wire signed [`CalcTempBus]          temp_b3_14_21_i;
wire signed [`CalcTempBus]          temp_b3_14_22_r;
wire signed [`CalcTempBus]          temp_b3_14_22_i;
wire signed [`CalcTempBus]          temp_b3_14_23_r;
wire signed [`CalcTempBus]          temp_b3_14_23_i;
wire signed [`CalcTempBus]          temp_b3_14_24_r;
wire signed [`CalcTempBus]          temp_b3_14_24_i;
wire signed [`CalcTempBus]          temp_b3_14_25_r;
wire signed [`CalcTempBus]          temp_b3_14_25_i;
wire signed [`CalcTempBus]          temp_b3_14_26_r;
wire signed [`CalcTempBus]          temp_b3_14_26_i;
wire signed [`CalcTempBus]          temp_b3_14_27_r;
wire signed [`CalcTempBus]          temp_b3_14_27_i;
wire signed [`CalcTempBus]          temp_b3_14_28_r;
wire signed [`CalcTempBus]          temp_b3_14_28_i;
wire signed [`CalcTempBus]          temp_b3_14_29_r;
wire signed [`CalcTempBus]          temp_b3_14_29_i;
wire signed [`CalcTempBus]          temp_b3_14_30_r;
wire signed [`CalcTempBus]          temp_b3_14_30_i;
wire signed [`CalcTempBus]          temp_b3_14_31_r;
wire signed [`CalcTempBus]          temp_b3_14_31_i;
wire signed [`CalcTempBus]          temp_b3_14_32_r;
wire signed [`CalcTempBus]          temp_b3_14_32_i;
wire signed [`CalcTempBus]          temp_b3_15_1_r;
wire signed [`CalcTempBus]          temp_b3_15_1_i;
wire signed [`CalcTempBus]          temp_b3_15_2_r;
wire signed [`CalcTempBus]          temp_b3_15_2_i;
wire signed [`CalcTempBus]          temp_b3_15_3_r;
wire signed [`CalcTempBus]          temp_b3_15_3_i;
wire signed [`CalcTempBus]          temp_b3_15_4_r;
wire signed [`CalcTempBus]          temp_b3_15_4_i;
wire signed [`CalcTempBus]          temp_b3_15_5_r;
wire signed [`CalcTempBus]          temp_b3_15_5_i;
wire signed [`CalcTempBus]          temp_b3_15_6_r;
wire signed [`CalcTempBus]          temp_b3_15_6_i;
wire signed [`CalcTempBus]          temp_b3_15_7_r;
wire signed [`CalcTempBus]          temp_b3_15_7_i;
wire signed [`CalcTempBus]          temp_b3_15_8_r;
wire signed [`CalcTempBus]          temp_b3_15_8_i;
wire signed [`CalcTempBus]          temp_b3_15_9_r;
wire signed [`CalcTempBus]          temp_b3_15_9_i;
wire signed [`CalcTempBus]          temp_b3_15_10_r;
wire signed [`CalcTempBus]          temp_b3_15_10_i;
wire signed [`CalcTempBus]          temp_b3_15_11_r;
wire signed [`CalcTempBus]          temp_b3_15_11_i;
wire signed [`CalcTempBus]          temp_b3_15_12_r;
wire signed [`CalcTempBus]          temp_b3_15_12_i;
wire signed [`CalcTempBus]          temp_b3_15_13_r;
wire signed [`CalcTempBus]          temp_b3_15_13_i;
wire signed [`CalcTempBus]          temp_b3_15_14_r;
wire signed [`CalcTempBus]          temp_b3_15_14_i;
wire signed [`CalcTempBus]          temp_b3_15_15_r;
wire signed [`CalcTempBus]          temp_b3_15_15_i;
wire signed [`CalcTempBus]          temp_b3_15_16_r;
wire signed [`CalcTempBus]          temp_b3_15_16_i;
wire signed [`CalcTempBus]          temp_b3_15_17_r;
wire signed [`CalcTempBus]          temp_b3_15_17_i;
wire signed [`CalcTempBus]          temp_b3_15_18_r;
wire signed [`CalcTempBus]          temp_b3_15_18_i;
wire signed [`CalcTempBus]          temp_b3_15_19_r;
wire signed [`CalcTempBus]          temp_b3_15_19_i;
wire signed [`CalcTempBus]          temp_b3_15_20_r;
wire signed [`CalcTempBus]          temp_b3_15_20_i;
wire signed [`CalcTempBus]          temp_b3_15_21_r;
wire signed [`CalcTempBus]          temp_b3_15_21_i;
wire signed [`CalcTempBus]          temp_b3_15_22_r;
wire signed [`CalcTempBus]          temp_b3_15_22_i;
wire signed [`CalcTempBus]          temp_b3_15_23_r;
wire signed [`CalcTempBus]          temp_b3_15_23_i;
wire signed [`CalcTempBus]          temp_b3_15_24_r;
wire signed [`CalcTempBus]          temp_b3_15_24_i;
wire signed [`CalcTempBus]          temp_b3_15_25_r;
wire signed [`CalcTempBus]          temp_b3_15_25_i;
wire signed [`CalcTempBus]          temp_b3_15_26_r;
wire signed [`CalcTempBus]          temp_b3_15_26_i;
wire signed [`CalcTempBus]          temp_b3_15_27_r;
wire signed [`CalcTempBus]          temp_b3_15_27_i;
wire signed [`CalcTempBus]          temp_b3_15_28_r;
wire signed [`CalcTempBus]          temp_b3_15_28_i;
wire signed [`CalcTempBus]          temp_b3_15_29_r;
wire signed [`CalcTempBus]          temp_b3_15_29_i;
wire signed [`CalcTempBus]          temp_b3_15_30_r;
wire signed [`CalcTempBus]          temp_b3_15_30_i;
wire signed [`CalcTempBus]          temp_b3_15_31_r;
wire signed [`CalcTempBus]          temp_b3_15_31_i;
wire signed [`CalcTempBus]          temp_b3_15_32_r;
wire signed [`CalcTempBus]          temp_b3_15_32_i;
wire signed [`CalcTempBus]          temp_b3_16_1_r;
wire signed [`CalcTempBus]          temp_b3_16_1_i;
wire signed [`CalcTempBus]          temp_b3_16_2_r;
wire signed [`CalcTempBus]          temp_b3_16_2_i;
wire signed [`CalcTempBus]          temp_b3_16_3_r;
wire signed [`CalcTempBus]          temp_b3_16_3_i;
wire signed [`CalcTempBus]          temp_b3_16_4_r;
wire signed [`CalcTempBus]          temp_b3_16_4_i;
wire signed [`CalcTempBus]          temp_b3_16_5_r;
wire signed [`CalcTempBus]          temp_b3_16_5_i;
wire signed [`CalcTempBus]          temp_b3_16_6_r;
wire signed [`CalcTempBus]          temp_b3_16_6_i;
wire signed [`CalcTempBus]          temp_b3_16_7_r;
wire signed [`CalcTempBus]          temp_b3_16_7_i;
wire signed [`CalcTempBus]          temp_b3_16_8_r;
wire signed [`CalcTempBus]          temp_b3_16_8_i;
wire signed [`CalcTempBus]          temp_b3_16_9_r;
wire signed [`CalcTempBus]          temp_b3_16_9_i;
wire signed [`CalcTempBus]          temp_b3_16_10_r;
wire signed [`CalcTempBus]          temp_b3_16_10_i;
wire signed [`CalcTempBus]          temp_b3_16_11_r;
wire signed [`CalcTempBus]          temp_b3_16_11_i;
wire signed [`CalcTempBus]          temp_b3_16_12_r;
wire signed [`CalcTempBus]          temp_b3_16_12_i;
wire signed [`CalcTempBus]          temp_b3_16_13_r;
wire signed [`CalcTempBus]          temp_b3_16_13_i;
wire signed [`CalcTempBus]          temp_b3_16_14_r;
wire signed [`CalcTempBus]          temp_b3_16_14_i;
wire signed [`CalcTempBus]          temp_b3_16_15_r;
wire signed [`CalcTempBus]          temp_b3_16_15_i;
wire signed [`CalcTempBus]          temp_b3_16_16_r;
wire signed [`CalcTempBus]          temp_b3_16_16_i;
wire signed [`CalcTempBus]          temp_b3_16_17_r;
wire signed [`CalcTempBus]          temp_b3_16_17_i;
wire signed [`CalcTempBus]          temp_b3_16_18_r;
wire signed [`CalcTempBus]          temp_b3_16_18_i;
wire signed [`CalcTempBus]          temp_b3_16_19_r;
wire signed [`CalcTempBus]          temp_b3_16_19_i;
wire signed [`CalcTempBus]          temp_b3_16_20_r;
wire signed [`CalcTempBus]          temp_b3_16_20_i;
wire signed [`CalcTempBus]          temp_b3_16_21_r;
wire signed [`CalcTempBus]          temp_b3_16_21_i;
wire signed [`CalcTempBus]          temp_b3_16_22_r;
wire signed [`CalcTempBus]          temp_b3_16_22_i;
wire signed [`CalcTempBus]          temp_b3_16_23_r;
wire signed [`CalcTempBus]          temp_b3_16_23_i;
wire signed [`CalcTempBus]          temp_b3_16_24_r;
wire signed [`CalcTempBus]          temp_b3_16_24_i;
wire signed [`CalcTempBus]          temp_b3_16_25_r;
wire signed [`CalcTempBus]          temp_b3_16_25_i;
wire signed [`CalcTempBus]          temp_b3_16_26_r;
wire signed [`CalcTempBus]          temp_b3_16_26_i;
wire signed [`CalcTempBus]          temp_b3_16_27_r;
wire signed [`CalcTempBus]          temp_b3_16_27_i;
wire signed [`CalcTempBus]          temp_b3_16_28_r;
wire signed [`CalcTempBus]          temp_b3_16_28_i;
wire signed [`CalcTempBus]          temp_b3_16_29_r;
wire signed [`CalcTempBus]          temp_b3_16_29_i;
wire signed [`CalcTempBus]          temp_b3_16_30_r;
wire signed [`CalcTempBus]          temp_b3_16_30_i;
wire signed [`CalcTempBus]          temp_b3_16_31_r;
wire signed [`CalcTempBus]          temp_b3_16_31_i;
wire signed [`CalcTempBus]          temp_b3_16_32_r;
wire signed [`CalcTempBus]          temp_b3_16_32_i;
wire signed [`CalcTempBus]          temp_b3_17_1_r;
wire signed [`CalcTempBus]          temp_b3_17_1_i;
wire signed [`CalcTempBus]          temp_b3_17_2_r;
wire signed [`CalcTempBus]          temp_b3_17_2_i;
wire signed [`CalcTempBus]          temp_b3_17_3_r;
wire signed [`CalcTempBus]          temp_b3_17_3_i;
wire signed [`CalcTempBus]          temp_b3_17_4_r;
wire signed [`CalcTempBus]          temp_b3_17_4_i;
wire signed [`CalcTempBus]          temp_b3_17_5_r;
wire signed [`CalcTempBus]          temp_b3_17_5_i;
wire signed [`CalcTempBus]          temp_b3_17_6_r;
wire signed [`CalcTempBus]          temp_b3_17_6_i;
wire signed [`CalcTempBus]          temp_b3_17_7_r;
wire signed [`CalcTempBus]          temp_b3_17_7_i;
wire signed [`CalcTempBus]          temp_b3_17_8_r;
wire signed [`CalcTempBus]          temp_b3_17_8_i;
wire signed [`CalcTempBus]          temp_b3_17_9_r;
wire signed [`CalcTempBus]          temp_b3_17_9_i;
wire signed [`CalcTempBus]          temp_b3_17_10_r;
wire signed [`CalcTempBus]          temp_b3_17_10_i;
wire signed [`CalcTempBus]          temp_b3_17_11_r;
wire signed [`CalcTempBus]          temp_b3_17_11_i;
wire signed [`CalcTempBus]          temp_b3_17_12_r;
wire signed [`CalcTempBus]          temp_b3_17_12_i;
wire signed [`CalcTempBus]          temp_b3_17_13_r;
wire signed [`CalcTempBus]          temp_b3_17_13_i;
wire signed [`CalcTempBus]          temp_b3_17_14_r;
wire signed [`CalcTempBus]          temp_b3_17_14_i;
wire signed [`CalcTempBus]          temp_b3_17_15_r;
wire signed [`CalcTempBus]          temp_b3_17_15_i;
wire signed [`CalcTempBus]          temp_b3_17_16_r;
wire signed [`CalcTempBus]          temp_b3_17_16_i;
wire signed [`CalcTempBus]          temp_b3_17_17_r;
wire signed [`CalcTempBus]          temp_b3_17_17_i;
wire signed [`CalcTempBus]          temp_b3_17_18_r;
wire signed [`CalcTempBus]          temp_b3_17_18_i;
wire signed [`CalcTempBus]          temp_b3_17_19_r;
wire signed [`CalcTempBus]          temp_b3_17_19_i;
wire signed [`CalcTempBus]          temp_b3_17_20_r;
wire signed [`CalcTempBus]          temp_b3_17_20_i;
wire signed [`CalcTempBus]          temp_b3_17_21_r;
wire signed [`CalcTempBus]          temp_b3_17_21_i;
wire signed [`CalcTempBus]          temp_b3_17_22_r;
wire signed [`CalcTempBus]          temp_b3_17_22_i;
wire signed [`CalcTempBus]          temp_b3_17_23_r;
wire signed [`CalcTempBus]          temp_b3_17_23_i;
wire signed [`CalcTempBus]          temp_b3_17_24_r;
wire signed [`CalcTempBus]          temp_b3_17_24_i;
wire signed [`CalcTempBus]          temp_b3_17_25_r;
wire signed [`CalcTempBus]          temp_b3_17_25_i;
wire signed [`CalcTempBus]          temp_b3_17_26_r;
wire signed [`CalcTempBus]          temp_b3_17_26_i;
wire signed [`CalcTempBus]          temp_b3_17_27_r;
wire signed [`CalcTempBus]          temp_b3_17_27_i;
wire signed [`CalcTempBus]          temp_b3_17_28_r;
wire signed [`CalcTempBus]          temp_b3_17_28_i;
wire signed [`CalcTempBus]          temp_b3_17_29_r;
wire signed [`CalcTempBus]          temp_b3_17_29_i;
wire signed [`CalcTempBus]          temp_b3_17_30_r;
wire signed [`CalcTempBus]          temp_b3_17_30_i;
wire signed [`CalcTempBus]          temp_b3_17_31_r;
wire signed [`CalcTempBus]          temp_b3_17_31_i;
wire signed [`CalcTempBus]          temp_b3_17_32_r;
wire signed [`CalcTempBus]          temp_b3_17_32_i;
wire signed [`CalcTempBus]          temp_b3_18_1_r;
wire signed [`CalcTempBus]          temp_b3_18_1_i;
wire signed [`CalcTempBus]          temp_b3_18_2_r;
wire signed [`CalcTempBus]          temp_b3_18_2_i;
wire signed [`CalcTempBus]          temp_b3_18_3_r;
wire signed [`CalcTempBus]          temp_b3_18_3_i;
wire signed [`CalcTempBus]          temp_b3_18_4_r;
wire signed [`CalcTempBus]          temp_b3_18_4_i;
wire signed [`CalcTempBus]          temp_b3_18_5_r;
wire signed [`CalcTempBus]          temp_b3_18_5_i;
wire signed [`CalcTempBus]          temp_b3_18_6_r;
wire signed [`CalcTempBus]          temp_b3_18_6_i;
wire signed [`CalcTempBus]          temp_b3_18_7_r;
wire signed [`CalcTempBus]          temp_b3_18_7_i;
wire signed [`CalcTempBus]          temp_b3_18_8_r;
wire signed [`CalcTempBus]          temp_b3_18_8_i;
wire signed [`CalcTempBus]          temp_b3_18_9_r;
wire signed [`CalcTempBus]          temp_b3_18_9_i;
wire signed [`CalcTempBus]          temp_b3_18_10_r;
wire signed [`CalcTempBus]          temp_b3_18_10_i;
wire signed [`CalcTempBus]          temp_b3_18_11_r;
wire signed [`CalcTempBus]          temp_b3_18_11_i;
wire signed [`CalcTempBus]          temp_b3_18_12_r;
wire signed [`CalcTempBus]          temp_b3_18_12_i;
wire signed [`CalcTempBus]          temp_b3_18_13_r;
wire signed [`CalcTempBus]          temp_b3_18_13_i;
wire signed [`CalcTempBus]          temp_b3_18_14_r;
wire signed [`CalcTempBus]          temp_b3_18_14_i;
wire signed [`CalcTempBus]          temp_b3_18_15_r;
wire signed [`CalcTempBus]          temp_b3_18_15_i;
wire signed [`CalcTempBus]          temp_b3_18_16_r;
wire signed [`CalcTempBus]          temp_b3_18_16_i;
wire signed [`CalcTempBus]          temp_b3_18_17_r;
wire signed [`CalcTempBus]          temp_b3_18_17_i;
wire signed [`CalcTempBus]          temp_b3_18_18_r;
wire signed [`CalcTempBus]          temp_b3_18_18_i;
wire signed [`CalcTempBus]          temp_b3_18_19_r;
wire signed [`CalcTempBus]          temp_b3_18_19_i;
wire signed [`CalcTempBus]          temp_b3_18_20_r;
wire signed [`CalcTempBus]          temp_b3_18_20_i;
wire signed [`CalcTempBus]          temp_b3_18_21_r;
wire signed [`CalcTempBus]          temp_b3_18_21_i;
wire signed [`CalcTempBus]          temp_b3_18_22_r;
wire signed [`CalcTempBus]          temp_b3_18_22_i;
wire signed [`CalcTempBus]          temp_b3_18_23_r;
wire signed [`CalcTempBus]          temp_b3_18_23_i;
wire signed [`CalcTempBus]          temp_b3_18_24_r;
wire signed [`CalcTempBus]          temp_b3_18_24_i;
wire signed [`CalcTempBus]          temp_b3_18_25_r;
wire signed [`CalcTempBus]          temp_b3_18_25_i;
wire signed [`CalcTempBus]          temp_b3_18_26_r;
wire signed [`CalcTempBus]          temp_b3_18_26_i;
wire signed [`CalcTempBus]          temp_b3_18_27_r;
wire signed [`CalcTempBus]          temp_b3_18_27_i;
wire signed [`CalcTempBus]          temp_b3_18_28_r;
wire signed [`CalcTempBus]          temp_b3_18_28_i;
wire signed [`CalcTempBus]          temp_b3_18_29_r;
wire signed [`CalcTempBus]          temp_b3_18_29_i;
wire signed [`CalcTempBus]          temp_b3_18_30_r;
wire signed [`CalcTempBus]          temp_b3_18_30_i;
wire signed [`CalcTempBus]          temp_b3_18_31_r;
wire signed [`CalcTempBus]          temp_b3_18_31_i;
wire signed [`CalcTempBus]          temp_b3_18_32_r;
wire signed [`CalcTempBus]          temp_b3_18_32_i;
wire signed [`CalcTempBus]          temp_b3_19_1_r;
wire signed [`CalcTempBus]          temp_b3_19_1_i;
wire signed [`CalcTempBus]          temp_b3_19_2_r;
wire signed [`CalcTempBus]          temp_b3_19_2_i;
wire signed [`CalcTempBus]          temp_b3_19_3_r;
wire signed [`CalcTempBus]          temp_b3_19_3_i;
wire signed [`CalcTempBus]          temp_b3_19_4_r;
wire signed [`CalcTempBus]          temp_b3_19_4_i;
wire signed [`CalcTempBus]          temp_b3_19_5_r;
wire signed [`CalcTempBus]          temp_b3_19_5_i;
wire signed [`CalcTempBus]          temp_b3_19_6_r;
wire signed [`CalcTempBus]          temp_b3_19_6_i;
wire signed [`CalcTempBus]          temp_b3_19_7_r;
wire signed [`CalcTempBus]          temp_b3_19_7_i;
wire signed [`CalcTempBus]          temp_b3_19_8_r;
wire signed [`CalcTempBus]          temp_b3_19_8_i;
wire signed [`CalcTempBus]          temp_b3_19_9_r;
wire signed [`CalcTempBus]          temp_b3_19_9_i;
wire signed [`CalcTempBus]          temp_b3_19_10_r;
wire signed [`CalcTempBus]          temp_b3_19_10_i;
wire signed [`CalcTempBus]          temp_b3_19_11_r;
wire signed [`CalcTempBus]          temp_b3_19_11_i;
wire signed [`CalcTempBus]          temp_b3_19_12_r;
wire signed [`CalcTempBus]          temp_b3_19_12_i;
wire signed [`CalcTempBus]          temp_b3_19_13_r;
wire signed [`CalcTempBus]          temp_b3_19_13_i;
wire signed [`CalcTempBus]          temp_b3_19_14_r;
wire signed [`CalcTempBus]          temp_b3_19_14_i;
wire signed [`CalcTempBus]          temp_b3_19_15_r;
wire signed [`CalcTempBus]          temp_b3_19_15_i;
wire signed [`CalcTempBus]          temp_b3_19_16_r;
wire signed [`CalcTempBus]          temp_b3_19_16_i;
wire signed [`CalcTempBus]          temp_b3_19_17_r;
wire signed [`CalcTempBus]          temp_b3_19_17_i;
wire signed [`CalcTempBus]          temp_b3_19_18_r;
wire signed [`CalcTempBus]          temp_b3_19_18_i;
wire signed [`CalcTempBus]          temp_b3_19_19_r;
wire signed [`CalcTempBus]          temp_b3_19_19_i;
wire signed [`CalcTempBus]          temp_b3_19_20_r;
wire signed [`CalcTempBus]          temp_b3_19_20_i;
wire signed [`CalcTempBus]          temp_b3_19_21_r;
wire signed [`CalcTempBus]          temp_b3_19_21_i;
wire signed [`CalcTempBus]          temp_b3_19_22_r;
wire signed [`CalcTempBus]          temp_b3_19_22_i;
wire signed [`CalcTempBus]          temp_b3_19_23_r;
wire signed [`CalcTempBus]          temp_b3_19_23_i;
wire signed [`CalcTempBus]          temp_b3_19_24_r;
wire signed [`CalcTempBus]          temp_b3_19_24_i;
wire signed [`CalcTempBus]          temp_b3_19_25_r;
wire signed [`CalcTempBus]          temp_b3_19_25_i;
wire signed [`CalcTempBus]          temp_b3_19_26_r;
wire signed [`CalcTempBus]          temp_b3_19_26_i;
wire signed [`CalcTempBus]          temp_b3_19_27_r;
wire signed [`CalcTempBus]          temp_b3_19_27_i;
wire signed [`CalcTempBus]          temp_b3_19_28_r;
wire signed [`CalcTempBus]          temp_b3_19_28_i;
wire signed [`CalcTempBus]          temp_b3_19_29_r;
wire signed [`CalcTempBus]          temp_b3_19_29_i;
wire signed [`CalcTempBus]          temp_b3_19_30_r;
wire signed [`CalcTempBus]          temp_b3_19_30_i;
wire signed [`CalcTempBus]          temp_b3_19_31_r;
wire signed [`CalcTempBus]          temp_b3_19_31_i;
wire signed [`CalcTempBus]          temp_b3_19_32_r;
wire signed [`CalcTempBus]          temp_b3_19_32_i;
wire signed [`CalcTempBus]          temp_b3_20_1_r;
wire signed [`CalcTempBus]          temp_b3_20_1_i;
wire signed [`CalcTempBus]          temp_b3_20_2_r;
wire signed [`CalcTempBus]          temp_b3_20_2_i;
wire signed [`CalcTempBus]          temp_b3_20_3_r;
wire signed [`CalcTempBus]          temp_b3_20_3_i;
wire signed [`CalcTempBus]          temp_b3_20_4_r;
wire signed [`CalcTempBus]          temp_b3_20_4_i;
wire signed [`CalcTempBus]          temp_b3_20_5_r;
wire signed [`CalcTempBus]          temp_b3_20_5_i;
wire signed [`CalcTempBus]          temp_b3_20_6_r;
wire signed [`CalcTempBus]          temp_b3_20_6_i;
wire signed [`CalcTempBus]          temp_b3_20_7_r;
wire signed [`CalcTempBus]          temp_b3_20_7_i;
wire signed [`CalcTempBus]          temp_b3_20_8_r;
wire signed [`CalcTempBus]          temp_b3_20_8_i;
wire signed [`CalcTempBus]          temp_b3_20_9_r;
wire signed [`CalcTempBus]          temp_b3_20_9_i;
wire signed [`CalcTempBus]          temp_b3_20_10_r;
wire signed [`CalcTempBus]          temp_b3_20_10_i;
wire signed [`CalcTempBus]          temp_b3_20_11_r;
wire signed [`CalcTempBus]          temp_b3_20_11_i;
wire signed [`CalcTempBus]          temp_b3_20_12_r;
wire signed [`CalcTempBus]          temp_b3_20_12_i;
wire signed [`CalcTempBus]          temp_b3_20_13_r;
wire signed [`CalcTempBus]          temp_b3_20_13_i;
wire signed [`CalcTempBus]          temp_b3_20_14_r;
wire signed [`CalcTempBus]          temp_b3_20_14_i;
wire signed [`CalcTempBus]          temp_b3_20_15_r;
wire signed [`CalcTempBus]          temp_b3_20_15_i;
wire signed [`CalcTempBus]          temp_b3_20_16_r;
wire signed [`CalcTempBus]          temp_b3_20_16_i;
wire signed [`CalcTempBus]          temp_b3_20_17_r;
wire signed [`CalcTempBus]          temp_b3_20_17_i;
wire signed [`CalcTempBus]          temp_b3_20_18_r;
wire signed [`CalcTempBus]          temp_b3_20_18_i;
wire signed [`CalcTempBus]          temp_b3_20_19_r;
wire signed [`CalcTempBus]          temp_b3_20_19_i;
wire signed [`CalcTempBus]          temp_b3_20_20_r;
wire signed [`CalcTempBus]          temp_b3_20_20_i;
wire signed [`CalcTempBus]          temp_b3_20_21_r;
wire signed [`CalcTempBus]          temp_b3_20_21_i;
wire signed [`CalcTempBus]          temp_b3_20_22_r;
wire signed [`CalcTempBus]          temp_b3_20_22_i;
wire signed [`CalcTempBus]          temp_b3_20_23_r;
wire signed [`CalcTempBus]          temp_b3_20_23_i;
wire signed [`CalcTempBus]          temp_b3_20_24_r;
wire signed [`CalcTempBus]          temp_b3_20_24_i;
wire signed [`CalcTempBus]          temp_b3_20_25_r;
wire signed [`CalcTempBus]          temp_b3_20_25_i;
wire signed [`CalcTempBus]          temp_b3_20_26_r;
wire signed [`CalcTempBus]          temp_b3_20_26_i;
wire signed [`CalcTempBus]          temp_b3_20_27_r;
wire signed [`CalcTempBus]          temp_b3_20_27_i;
wire signed [`CalcTempBus]          temp_b3_20_28_r;
wire signed [`CalcTempBus]          temp_b3_20_28_i;
wire signed [`CalcTempBus]          temp_b3_20_29_r;
wire signed [`CalcTempBus]          temp_b3_20_29_i;
wire signed [`CalcTempBus]          temp_b3_20_30_r;
wire signed [`CalcTempBus]          temp_b3_20_30_i;
wire signed [`CalcTempBus]          temp_b3_20_31_r;
wire signed [`CalcTempBus]          temp_b3_20_31_i;
wire signed [`CalcTempBus]          temp_b3_20_32_r;
wire signed [`CalcTempBus]          temp_b3_20_32_i;
wire signed [`CalcTempBus]          temp_b3_21_1_r;
wire signed [`CalcTempBus]          temp_b3_21_1_i;
wire signed [`CalcTempBus]          temp_b3_21_2_r;
wire signed [`CalcTempBus]          temp_b3_21_2_i;
wire signed [`CalcTempBus]          temp_b3_21_3_r;
wire signed [`CalcTempBus]          temp_b3_21_3_i;
wire signed [`CalcTempBus]          temp_b3_21_4_r;
wire signed [`CalcTempBus]          temp_b3_21_4_i;
wire signed [`CalcTempBus]          temp_b3_21_5_r;
wire signed [`CalcTempBus]          temp_b3_21_5_i;
wire signed [`CalcTempBus]          temp_b3_21_6_r;
wire signed [`CalcTempBus]          temp_b3_21_6_i;
wire signed [`CalcTempBus]          temp_b3_21_7_r;
wire signed [`CalcTempBus]          temp_b3_21_7_i;
wire signed [`CalcTempBus]          temp_b3_21_8_r;
wire signed [`CalcTempBus]          temp_b3_21_8_i;
wire signed [`CalcTempBus]          temp_b3_21_9_r;
wire signed [`CalcTempBus]          temp_b3_21_9_i;
wire signed [`CalcTempBus]          temp_b3_21_10_r;
wire signed [`CalcTempBus]          temp_b3_21_10_i;
wire signed [`CalcTempBus]          temp_b3_21_11_r;
wire signed [`CalcTempBus]          temp_b3_21_11_i;
wire signed [`CalcTempBus]          temp_b3_21_12_r;
wire signed [`CalcTempBus]          temp_b3_21_12_i;
wire signed [`CalcTempBus]          temp_b3_21_13_r;
wire signed [`CalcTempBus]          temp_b3_21_13_i;
wire signed [`CalcTempBus]          temp_b3_21_14_r;
wire signed [`CalcTempBus]          temp_b3_21_14_i;
wire signed [`CalcTempBus]          temp_b3_21_15_r;
wire signed [`CalcTempBus]          temp_b3_21_15_i;
wire signed [`CalcTempBus]          temp_b3_21_16_r;
wire signed [`CalcTempBus]          temp_b3_21_16_i;
wire signed [`CalcTempBus]          temp_b3_21_17_r;
wire signed [`CalcTempBus]          temp_b3_21_17_i;
wire signed [`CalcTempBus]          temp_b3_21_18_r;
wire signed [`CalcTempBus]          temp_b3_21_18_i;
wire signed [`CalcTempBus]          temp_b3_21_19_r;
wire signed [`CalcTempBus]          temp_b3_21_19_i;
wire signed [`CalcTempBus]          temp_b3_21_20_r;
wire signed [`CalcTempBus]          temp_b3_21_20_i;
wire signed [`CalcTempBus]          temp_b3_21_21_r;
wire signed [`CalcTempBus]          temp_b3_21_21_i;
wire signed [`CalcTempBus]          temp_b3_21_22_r;
wire signed [`CalcTempBus]          temp_b3_21_22_i;
wire signed [`CalcTempBus]          temp_b3_21_23_r;
wire signed [`CalcTempBus]          temp_b3_21_23_i;
wire signed [`CalcTempBus]          temp_b3_21_24_r;
wire signed [`CalcTempBus]          temp_b3_21_24_i;
wire signed [`CalcTempBus]          temp_b3_21_25_r;
wire signed [`CalcTempBus]          temp_b3_21_25_i;
wire signed [`CalcTempBus]          temp_b3_21_26_r;
wire signed [`CalcTempBus]          temp_b3_21_26_i;
wire signed [`CalcTempBus]          temp_b3_21_27_r;
wire signed [`CalcTempBus]          temp_b3_21_27_i;
wire signed [`CalcTempBus]          temp_b3_21_28_r;
wire signed [`CalcTempBus]          temp_b3_21_28_i;
wire signed [`CalcTempBus]          temp_b3_21_29_r;
wire signed [`CalcTempBus]          temp_b3_21_29_i;
wire signed [`CalcTempBus]          temp_b3_21_30_r;
wire signed [`CalcTempBus]          temp_b3_21_30_i;
wire signed [`CalcTempBus]          temp_b3_21_31_r;
wire signed [`CalcTempBus]          temp_b3_21_31_i;
wire signed [`CalcTempBus]          temp_b3_21_32_r;
wire signed [`CalcTempBus]          temp_b3_21_32_i;
wire signed [`CalcTempBus]          temp_b3_22_1_r;
wire signed [`CalcTempBus]          temp_b3_22_1_i;
wire signed [`CalcTempBus]          temp_b3_22_2_r;
wire signed [`CalcTempBus]          temp_b3_22_2_i;
wire signed [`CalcTempBus]          temp_b3_22_3_r;
wire signed [`CalcTempBus]          temp_b3_22_3_i;
wire signed [`CalcTempBus]          temp_b3_22_4_r;
wire signed [`CalcTempBus]          temp_b3_22_4_i;
wire signed [`CalcTempBus]          temp_b3_22_5_r;
wire signed [`CalcTempBus]          temp_b3_22_5_i;
wire signed [`CalcTempBus]          temp_b3_22_6_r;
wire signed [`CalcTempBus]          temp_b3_22_6_i;
wire signed [`CalcTempBus]          temp_b3_22_7_r;
wire signed [`CalcTempBus]          temp_b3_22_7_i;
wire signed [`CalcTempBus]          temp_b3_22_8_r;
wire signed [`CalcTempBus]          temp_b3_22_8_i;
wire signed [`CalcTempBus]          temp_b3_22_9_r;
wire signed [`CalcTempBus]          temp_b3_22_9_i;
wire signed [`CalcTempBus]          temp_b3_22_10_r;
wire signed [`CalcTempBus]          temp_b3_22_10_i;
wire signed [`CalcTempBus]          temp_b3_22_11_r;
wire signed [`CalcTempBus]          temp_b3_22_11_i;
wire signed [`CalcTempBus]          temp_b3_22_12_r;
wire signed [`CalcTempBus]          temp_b3_22_12_i;
wire signed [`CalcTempBus]          temp_b3_22_13_r;
wire signed [`CalcTempBus]          temp_b3_22_13_i;
wire signed [`CalcTempBus]          temp_b3_22_14_r;
wire signed [`CalcTempBus]          temp_b3_22_14_i;
wire signed [`CalcTempBus]          temp_b3_22_15_r;
wire signed [`CalcTempBus]          temp_b3_22_15_i;
wire signed [`CalcTempBus]          temp_b3_22_16_r;
wire signed [`CalcTempBus]          temp_b3_22_16_i;
wire signed [`CalcTempBus]          temp_b3_22_17_r;
wire signed [`CalcTempBus]          temp_b3_22_17_i;
wire signed [`CalcTempBus]          temp_b3_22_18_r;
wire signed [`CalcTempBus]          temp_b3_22_18_i;
wire signed [`CalcTempBus]          temp_b3_22_19_r;
wire signed [`CalcTempBus]          temp_b3_22_19_i;
wire signed [`CalcTempBus]          temp_b3_22_20_r;
wire signed [`CalcTempBus]          temp_b3_22_20_i;
wire signed [`CalcTempBus]          temp_b3_22_21_r;
wire signed [`CalcTempBus]          temp_b3_22_21_i;
wire signed [`CalcTempBus]          temp_b3_22_22_r;
wire signed [`CalcTempBus]          temp_b3_22_22_i;
wire signed [`CalcTempBus]          temp_b3_22_23_r;
wire signed [`CalcTempBus]          temp_b3_22_23_i;
wire signed [`CalcTempBus]          temp_b3_22_24_r;
wire signed [`CalcTempBus]          temp_b3_22_24_i;
wire signed [`CalcTempBus]          temp_b3_22_25_r;
wire signed [`CalcTempBus]          temp_b3_22_25_i;
wire signed [`CalcTempBus]          temp_b3_22_26_r;
wire signed [`CalcTempBus]          temp_b3_22_26_i;
wire signed [`CalcTempBus]          temp_b3_22_27_r;
wire signed [`CalcTempBus]          temp_b3_22_27_i;
wire signed [`CalcTempBus]          temp_b3_22_28_r;
wire signed [`CalcTempBus]          temp_b3_22_28_i;
wire signed [`CalcTempBus]          temp_b3_22_29_r;
wire signed [`CalcTempBus]          temp_b3_22_29_i;
wire signed [`CalcTempBus]          temp_b3_22_30_r;
wire signed [`CalcTempBus]          temp_b3_22_30_i;
wire signed [`CalcTempBus]          temp_b3_22_31_r;
wire signed [`CalcTempBus]          temp_b3_22_31_i;
wire signed [`CalcTempBus]          temp_b3_22_32_r;
wire signed [`CalcTempBus]          temp_b3_22_32_i;
wire signed [`CalcTempBus]          temp_b3_23_1_r;
wire signed [`CalcTempBus]          temp_b3_23_1_i;
wire signed [`CalcTempBus]          temp_b3_23_2_r;
wire signed [`CalcTempBus]          temp_b3_23_2_i;
wire signed [`CalcTempBus]          temp_b3_23_3_r;
wire signed [`CalcTempBus]          temp_b3_23_3_i;
wire signed [`CalcTempBus]          temp_b3_23_4_r;
wire signed [`CalcTempBus]          temp_b3_23_4_i;
wire signed [`CalcTempBus]          temp_b3_23_5_r;
wire signed [`CalcTempBus]          temp_b3_23_5_i;
wire signed [`CalcTempBus]          temp_b3_23_6_r;
wire signed [`CalcTempBus]          temp_b3_23_6_i;
wire signed [`CalcTempBus]          temp_b3_23_7_r;
wire signed [`CalcTempBus]          temp_b3_23_7_i;
wire signed [`CalcTempBus]          temp_b3_23_8_r;
wire signed [`CalcTempBus]          temp_b3_23_8_i;
wire signed [`CalcTempBus]          temp_b3_23_9_r;
wire signed [`CalcTempBus]          temp_b3_23_9_i;
wire signed [`CalcTempBus]          temp_b3_23_10_r;
wire signed [`CalcTempBus]          temp_b3_23_10_i;
wire signed [`CalcTempBus]          temp_b3_23_11_r;
wire signed [`CalcTempBus]          temp_b3_23_11_i;
wire signed [`CalcTempBus]          temp_b3_23_12_r;
wire signed [`CalcTempBus]          temp_b3_23_12_i;
wire signed [`CalcTempBus]          temp_b3_23_13_r;
wire signed [`CalcTempBus]          temp_b3_23_13_i;
wire signed [`CalcTempBus]          temp_b3_23_14_r;
wire signed [`CalcTempBus]          temp_b3_23_14_i;
wire signed [`CalcTempBus]          temp_b3_23_15_r;
wire signed [`CalcTempBus]          temp_b3_23_15_i;
wire signed [`CalcTempBus]          temp_b3_23_16_r;
wire signed [`CalcTempBus]          temp_b3_23_16_i;
wire signed [`CalcTempBus]          temp_b3_23_17_r;
wire signed [`CalcTempBus]          temp_b3_23_17_i;
wire signed [`CalcTempBus]          temp_b3_23_18_r;
wire signed [`CalcTempBus]          temp_b3_23_18_i;
wire signed [`CalcTempBus]          temp_b3_23_19_r;
wire signed [`CalcTempBus]          temp_b3_23_19_i;
wire signed [`CalcTempBus]          temp_b3_23_20_r;
wire signed [`CalcTempBus]          temp_b3_23_20_i;
wire signed [`CalcTempBus]          temp_b3_23_21_r;
wire signed [`CalcTempBus]          temp_b3_23_21_i;
wire signed [`CalcTempBus]          temp_b3_23_22_r;
wire signed [`CalcTempBus]          temp_b3_23_22_i;
wire signed [`CalcTempBus]          temp_b3_23_23_r;
wire signed [`CalcTempBus]          temp_b3_23_23_i;
wire signed [`CalcTempBus]          temp_b3_23_24_r;
wire signed [`CalcTempBus]          temp_b3_23_24_i;
wire signed [`CalcTempBus]          temp_b3_23_25_r;
wire signed [`CalcTempBus]          temp_b3_23_25_i;
wire signed [`CalcTempBus]          temp_b3_23_26_r;
wire signed [`CalcTempBus]          temp_b3_23_26_i;
wire signed [`CalcTempBus]          temp_b3_23_27_r;
wire signed [`CalcTempBus]          temp_b3_23_27_i;
wire signed [`CalcTempBus]          temp_b3_23_28_r;
wire signed [`CalcTempBus]          temp_b3_23_28_i;
wire signed [`CalcTempBus]          temp_b3_23_29_r;
wire signed [`CalcTempBus]          temp_b3_23_29_i;
wire signed [`CalcTempBus]          temp_b3_23_30_r;
wire signed [`CalcTempBus]          temp_b3_23_30_i;
wire signed [`CalcTempBus]          temp_b3_23_31_r;
wire signed [`CalcTempBus]          temp_b3_23_31_i;
wire signed [`CalcTempBus]          temp_b3_23_32_r;
wire signed [`CalcTempBus]          temp_b3_23_32_i;
wire signed [`CalcTempBus]          temp_b3_24_1_r;
wire signed [`CalcTempBus]          temp_b3_24_1_i;
wire signed [`CalcTempBus]          temp_b3_24_2_r;
wire signed [`CalcTempBus]          temp_b3_24_2_i;
wire signed [`CalcTempBus]          temp_b3_24_3_r;
wire signed [`CalcTempBus]          temp_b3_24_3_i;
wire signed [`CalcTempBus]          temp_b3_24_4_r;
wire signed [`CalcTempBus]          temp_b3_24_4_i;
wire signed [`CalcTempBus]          temp_b3_24_5_r;
wire signed [`CalcTempBus]          temp_b3_24_5_i;
wire signed [`CalcTempBus]          temp_b3_24_6_r;
wire signed [`CalcTempBus]          temp_b3_24_6_i;
wire signed [`CalcTempBus]          temp_b3_24_7_r;
wire signed [`CalcTempBus]          temp_b3_24_7_i;
wire signed [`CalcTempBus]          temp_b3_24_8_r;
wire signed [`CalcTempBus]          temp_b3_24_8_i;
wire signed [`CalcTempBus]          temp_b3_24_9_r;
wire signed [`CalcTempBus]          temp_b3_24_9_i;
wire signed [`CalcTempBus]          temp_b3_24_10_r;
wire signed [`CalcTempBus]          temp_b3_24_10_i;
wire signed [`CalcTempBus]          temp_b3_24_11_r;
wire signed [`CalcTempBus]          temp_b3_24_11_i;
wire signed [`CalcTempBus]          temp_b3_24_12_r;
wire signed [`CalcTempBus]          temp_b3_24_12_i;
wire signed [`CalcTempBus]          temp_b3_24_13_r;
wire signed [`CalcTempBus]          temp_b3_24_13_i;
wire signed [`CalcTempBus]          temp_b3_24_14_r;
wire signed [`CalcTempBus]          temp_b3_24_14_i;
wire signed [`CalcTempBus]          temp_b3_24_15_r;
wire signed [`CalcTempBus]          temp_b3_24_15_i;
wire signed [`CalcTempBus]          temp_b3_24_16_r;
wire signed [`CalcTempBus]          temp_b3_24_16_i;
wire signed [`CalcTempBus]          temp_b3_24_17_r;
wire signed [`CalcTempBus]          temp_b3_24_17_i;
wire signed [`CalcTempBus]          temp_b3_24_18_r;
wire signed [`CalcTempBus]          temp_b3_24_18_i;
wire signed [`CalcTempBus]          temp_b3_24_19_r;
wire signed [`CalcTempBus]          temp_b3_24_19_i;
wire signed [`CalcTempBus]          temp_b3_24_20_r;
wire signed [`CalcTempBus]          temp_b3_24_20_i;
wire signed [`CalcTempBus]          temp_b3_24_21_r;
wire signed [`CalcTempBus]          temp_b3_24_21_i;
wire signed [`CalcTempBus]          temp_b3_24_22_r;
wire signed [`CalcTempBus]          temp_b3_24_22_i;
wire signed [`CalcTempBus]          temp_b3_24_23_r;
wire signed [`CalcTempBus]          temp_b3_24_23_i;
wire signed [`CalcTempBus]          temp_b3_24_24_r;
wire signed [`CalcTempBus]          temp_b3_24_24_i;
wire signed [`CalcTempBus]          temp_b3_24_25_r;
wire signed [`CalcTempBus]          temp_b3_24_25_i;
wire signed [`CalcTempBus]          temp_b3_24_26_r;
wire signed [`CalcTempBus]          temp_b3_24_26_i;
wire signed [`CalcTempBus]          temp_b3_24_27_r;
wire signed [`CalcTempBus]          temp_b3_24_27_i;
wire signed [`CalcTempBus]          temp_b3_24_28_r;
wire signed [`CalcTempBus]          temp_b3_24_28_i;
wire signed [`CalcTempBus]          temp_b3_24_29_r;
wire signed [`CalcTempBus]          temp_b3_24_29_i;
wire signed [`CalcTempBus]          temp_b3_24_30_r;
wire signed [`CalcTempBus]          temp_b3_24_30_i;
wire signed [`CalcTempBus]          temp_b3_24_31_r;
wire signed [`CalcTempBus]          temp_b3_24_31_i;
wire signed [`CalcTempBus]          temp_b3_24_32_r;
wire signed [`CalcTempBus]          temp_b3_24_32_i;
wire signed [`CalcTempBus]          temp_b3_25_1_r;
wire signed [`CalcTempBus]          temp_b3_25_1_i;
wire signed [`CalcTempBus]          temp_b3_25_2_r;
wire signed [`CalcTempBus]          temp_b3_25_2_i;
wire signed [`CalcTempBus]          temp_b3_25_3_r;
wire signed [`CalcTempBus]          temp_b3_25_3_i;
wire signed [`CalcTempBus]          temp_b3_25_4_r;
wire signed [`CalcTempBus]          temp_b3_25_4_i;
wire signed [`CalcTempBus]          temp_b3_25_5_r;
wire signed [`CalcTempBus]          temp_b3_25_5_i;
wire signed [`CalcTempBus]          temp_b3_25_6_r;
wire signed [`CalcTempBus]          temp_b3_25_6_i;
wire signed [`CalcTempBus]          temp_b3_25_7_r;
wire signed [`CalcTempBus]          temp_b3_25_7_i;
wire signed [`CalcTempBus]          temp_b3_25_8_r;
wire signed [`CalcTempBus]          temp_b3_25_8_i;
wire signed [`CalcTempBus]          temp_b3_25_9_r;
wire signed [`CalcTempBus]          temp_b3_25_9_i;
wire signed [`CalcTempBus]          temp_b3_25_10_r;
wire signed [`CalcTempBus]          temp_b3_25_10_i;
wire signed [`CalcTempBus]          temp_b3_25_11_r;
wire signed [`CalcTempBus]          temp_b3_25_11_i;
wire signed [`CalcTempBus]          temp_b3_25_12_r;
wire signed [`CalcTempBus]          temp_b3_25_12_i;
wire signed [`CalcTempBus]          temp_b3_25_13_r;
wire signed [`CalcTempBus]          temp_b3_25_13_i;
wire signed [`CalcTempBus]          temp_b3_25_14_r;
wire signed [`CalcTempBus]          temp_b3_25_14_i;
wire signed [`CalcTempBus]          temp_b3_25_15_r;
wire signed [`CalcTempBus]          temp_b3_25_15_i;
wire signed [`CalcTempBus]          temp_b3_25_16_r;
wire signed [`CalcTempBus]          temp_b3_25_16_i;
wire signed [`CalcTempBus]          temp_b3_25_17_r;
wire signed [`CalcTempBus]          temp_b3_25_17_i;
wire signed [`CalcTempBus]          temp_b3_25_18_r;
wire signed [`CalcTempBus]          temp_b3_25_18_i;
wire signed [`CalcTempBus]          temp_b3_25_19_r;
wire signed [`CalcTempBus]          temp_b3_25_19_i;
wire signed [`CalcTempBus]          temp_b3_25_20_r;
wire signed [`CalcTempBus]          temp_b3_25_20_i;
wire signed [`CalcTempBus]          temp_b3_25_21_r;
wire signed [`CalcTempBus]          temp_b3_25_21_i;
wire signed [`CalcTempBus]          temp_b3_25_22_r;
wire signed [`CalcTempBus]          temp_b3_25_22_i;
wire signed [`CalcTempBus]          temp_b3_25_23_r;
wire signed [`CalcTempBus]          temp_b3_25_23_i;
wire signed [`CalcTempBus]          temp_b3_25_24_r;
wire signed [`CalcTempBus]          temp_b3_25_24_i;
wire signed [`CalcTempBus]          temp_b3_25_25_r;
wire signed [`CalcTempBus]          temp_b3_25_25_i;
wire signed [`CalcTempBus]          temp_b3_25_26_r;
wire signed [`CalcTempBus]          temp_b3_25_26_i;
wire signed [`CalcTempBus]          temp_b3_25_27_r;
wire signed [`CalcTempBus]          temp_b3_25_27_i;
wire signed [`CalcTempBus]          temp_b3_25_28_r;
wire signed [`CalcTempBus]          temp_b3_25_28_i;
wire signed [`CalcTempBus]          temp_b3_25_29_r;
wire signed [`CalcTempBus]          temp_b3_25_29_i;
wire signed [`CalcTempBus]          temp_b3_25_30_r;
wire signed [`CalcTempBus]          temp_b3_25_30_i;
wire signed [`CalcTempBus]          temp_b3_25_31_r;
wire signed [`CalcTempBus]          temp_b3_25_31_i;
wire signed [`CalcTempBus]          temp_b3_25_32_r;
wire signed [`CalcTempBus]          temp_b3_25_32_i;
wire signed [`CalcTempBus]          temp_b3_26_1_r;
wire signed [`CalcTempBus]          temp_b3_26_1_i;
wire signed [`CalcTempBus]          temp_b3_26_2_r;
wire signed [`CalcTempBus]          temp_b3_26_2_i;
wire signed [`CalcTempBus]          temp_b3_26_3_r;
wire signed [`CalcTempBus]          temp_b3_26_3_i;
wire signed [`CalcTempBus]          temp_b3_26_4_r;
wire signed [`CalcTempBus]          temp_b3_26_4_i;
wire signed [`CalcTempBus]          temp_b3_26_5_r;
wire signed [`CalcTempBus]          temp_b3_26_5_i;
wire signed [`CalcTempBus]          temp_b3_26_6_r;
wire signed [`CalcTempBus]          temp_b3_26_6_i;
wire signed [`CalcTempBus]          temp_b3_26_7_r;
wire signed [`CalcTempBus]          temp_b3_26_7_i;
wire signed [`CalcTempBus]          temp_b3_26_8_r;
wire signed [`CalcTempBus]          temp_b3_26_8_i;
wire signed [`CalcTempBus]          temp_b3_26_9_r;
wire signed [`CalcTempBus]          temp_b3_26_9_i;
wire signed [`CalcTempBus]          temp_b3_26_10_r;
wire signed [`CalcTempBus]          temp_b3_26_10_i;
wire signed [`CalcTempBus]          temp_b3_26_11_r;
wire signed [`CalcTempBus]          temp_b3_26_11_i;
wire signed [`CalcTempBus]          temp_b3_26_12_r;
wire signed [`CalcTempBus]          temp_b3_26_12_i;
wire signed [`CalcTempBus]          temp_b3_26_13_r;
wire signed [`CalcTempBus]          temp_b3_26_13_i;
wire signed [`CalcTempBus]          temp_b3_26_14_r;
wire signed [`CalcTempBus]          temp_b3_26_14_i;
wire signed [`CalcTempBus]          temp_b3_26_15_r;
wire signed [`CalcTempBus]          temp_b3_26_15_i;
wire signed [`CalcTempBus]          temp_b3_26_16_r;
wire signed [`CalcTempBus]          temp_b3_26_16_i;
wire signed [`CalcTempBus]          temp_b3_26_17_r;
wire signed [`CalcTempBus]          temp_b3_26_17_i;
wire signed [`CalcTempBus]          temp_b3_26_18_r;
wire signed [`CalcTempBus]          temp_b3_26_18_i;
wire signed [`CalcTempBus]          temp_b3_26_19_r;
wire signed [`CalcTempBus]          temp_b3_26_19_i;
wire signed [`CalcTempBus]          temp_b3_26_20_r;
wire signed [`CalcTempBus]          temp_b3_26_20_i;
wire signed [`CalcTempBus]          temp_b3_26_21_r;
wire signed [`CalcTempBus]          temp_b3_26_21_i;
wire signed [`CalcTempBus]          temp_b3_26_22_r;
wire signed [`CalcTempBus]          temp_b3_26_22_i;
wire signed [`CalcTempBus]          temp_b3_26_23_r;
wire signed [`CalcTempBus]          temp_b3_26_23_i;
wire signed [`CalcTempBus]          temp_b3_26_24_r;
wire signed [`CalcTempBus]          temp_b3_26_24_i;
wire signed [`CalcTempBus]          temp_b3_26_25_r;
wire signed [`CalcTempBus]          temp_b3_26_25_i;
wire signed [`CalcTempBus]          temp_b3_26_26_r;
wire signed [`CalcTempBus]          temp_b3_26_26_i;
wire signed [`CalcTempBus]          temp_b3_26_27_r;
wire signed [`CalcTempBus]          temp_b3_26_27_i;
wire signed [`CalcTempBus]          temp_b3_26_28_r;
wire signed [`CalcTempBus]          temp_b3_26_28_i;
wire signed [`CalcTempBus]          temp_b3_26_29_r;
wire signed [`CalcTempBus]          temp_b3_26_29_i;
wire signed [`CalcTempBus]          temp_b3_26_30_r;
wire signed [`CalcTempBus]          temp_b3_26_30_i;
wire signed [`CalcTempBus]          temp_b3_26_31_r;
wire signed [`CalcTempBus]          temp_b3_26_31_i;
wire signed [`CalcTempBus]          temp_b3_26_32_r;
wire signed [`CalcTempBus]          temp_b3_26_32_i;
wire signed [`CalcTempBus]          temp_b3_27_1_r;
wire signed [`CalcTempBus]          temp_b3_27_1_i;
wire signed [`CalcTempBus]          temp_b3_27_2_r;
wire signed [`CalcTempBus]          temp_b3_27_2_i;
wire signed [`CalcTempBus]          temp_b3_27_3_r;
wire signed [`CalcTempBus]          temp_b3_27_3_i;
wire signed [`CalcTempBus]          temp_b3_27_4_r;
wire signed [`CalcTempBus]          temp_b3_27_4_i;
wire signed [`CalcTempBus]          temp_b3_27_5_r;
wire signed [`CalcTempBus]          temp_b3_27_5_i;
wire signed [`CalcTempBus]          temp_b3_27_6_r;
wire signed [`CalcTempBus]          temp_b3_27_6_i;
wire signed [`CalcTempBus]          temp_b3_27_7_r;
wire signed [`CalcTempBus]          temp_b3_27_7_i;
wire signed [`CalcTempBus]          temp_b3_27_8_r;
wire signed [`CalcTempBus]          temp_b3_27_8_i;
wire signed [`CalcTempBus]          temp_b3_27_9_r;
wire signed [`CalcTempBus]          temp_b3_27_9_i;
wire signed [`CalcTempBus]          temp_b3_27_10_r;
wire signed [`CalcTempBus]          temp_b3_27_10_i;
wire signed [`CalcTempBus]          temp_b3_27_11_r;
wire signed [`CalcTempBus]          temp_b3_27_11_i;
wire signed [`CalcTempBus]          temp_b3_27_12_r;
wire signed [`CalcTempBus]          temp_b3_27_12_i;
wire signed [`CalcTempBus]          temp_b3_27_13_r;
wire signed [`CalcTempBus]          temp_b3_27_13_i;
wire signed [`CalcTempBus]          temp_b3_27_14_r;
wire signed [`CalcTempBus]          temp_b3_27_14_i;
wire signed [`CalcTempBus]          temp_b3_27_15_r;
wire signed [`CalcTempBus]          temp_b3_27_15_i;
wire signed [`CalcTempBus]          temp_b3_27_16_r;
wire signed [`CalcTempBus]          temp_b3_27_16_i;
wire signed [`CalcTempBus]          temp_b3_27_17_r;
wire signed [`CalcTempBus]          temp_b3_27_17_i;
wire signed [`CalcTempBus]          temp_b3_27_18_r;
wire signed [`CalcTempBus]          temp_b3_27_18_i;
wire signed [`CalcTempBus]          temp_b3_27_19_r;
wire signed [`CalcTempBus]          temp_b3_27_19_i;
wire signed [`CalcTempBus]          temp_b3_27_20_r;
wire signed [`CalcTempBus]          temp_b3_27_20_i;
wire signed [`CalcTempBus]          temp_b3_27_21_r;
wire signed [`CalcTempBus]          temp_b3_27_21_i;
wire signed [`CalcTempBus]          temp_b3_27_22_r;
wire signed [`CalcTempBus]          temp_b3_27_22_i;
wire signed [`CalcTempBus]          temp_b3_27_23_r;
wire signed [`CalcTempBus]          temp_b3_27_23_i;
wire signed [`CalcTempBus]          temp_b3_27_24_r;
wire signed [`CalcTempBus]          temp_b3_27_24_i;
wire signed [`CalcTempBus]          temp_b3_27_25_r;
wire signed [`CalcTempBus]          temp_b3_27_25_i;
wire signed [`CalcTempBus]          temp_b3_27_26_r;
wire signed [`CalcTempBus]          temp_b3_27_26_i;
wire signed [`CalcTempBus]          temp_b3_27_27_r;
wire signed [`CalcTempBus]          temp_b3_27_27_i;
wire signed [`CalcTempBus]          temp_b3_27_28_r;
wire signed [`CalcTempBus]          temp_b3_27_28_i;
wire signed [`CalcTempBus]          temp_b3_27_29_r;
wire signed [`CalcTempBus]          temp_b3_27_29_i;
wire signed [`CalcTempBus]          temp_b3_27_30_r;
wire signed [`CalcTempBus]          temp_b3_27_30_i;
wire signed [`CalcTempBus]          temp_b3_27_31_r;
wire signed [`CalcTempBus]          temp_b3_27_31_i;
wire signed [`CalcTempBus]          temp_b3_27_32_r;
wire signed [`CalcTempBus]          temp_b3_27_32_i;
wire signed [`CalcTempBus]          temp_b3_28_1_r;
wire signed [`CalcTempBus]          temp_b3_28_1_i;
wire signed [`CalcTempBus]          temp_b3_28_2_r;
wire signed [`CalcTempBus]          temp_b3_28_2_i;
wire signed [`CalcTempBus]          temp_b3_28_3_r;
wire signed [`CalcTempBus]          temp_b3_28_3_i;
wire signed [`CalcTempBus]          temp_b3_28_4_r;
wire signed [`CalcTempBus]          temp_b3_28_4_i;
wire signed [`CalcTempBus]          temp_b3_28_5_r;
wire signed [`CalcTempBus]          temp_b3_28_5_i;
wire signed [`CalcTempBus]          temp_b3_28_6_r;
wire signed [`CalcTempBus]          temp_b3_28_6_i;
wire signed [`CalcTempBus]          temp_b3_28_7_r;
wire signed [`CalcTempBus]          temp_b3_28_7_i;
wire signed [`CalcTempBus]          temp_b3_28_8_r;
wire signed [`CalcTempBus]          temp_b3_28_8_i;
wire signed [`CalcTempBus]          temp_b3_28_9_r;
wire signed [`CalcTempBus]          temp_b3_28_9_i;
wire signed [`CalcTempBus]          temp_b3_28_10_r;
wire signed [`CalcTempBus]          temp_b3_28_10_i;
wire signed [`CalcTempBus]          temp_b3_28_11_r;
wire signed [`CalcTempBus]          temp_b3_28_11_i;
wire signed [`CalcTempBus]          temp_b3_28_12_r;
wire signed [`CalcTempBus]          temp_b3_28_12_i;
wire signed [`CalcTempBus]          temp_b3_28_13_r;
wire signed [`CalcTempBus]          temp_b3_28_13_i;
wire signed [`CalcTempBus]          temp_b3_28_14_r;
wire signed [`CalcTempBus]          temp_b3_28_14_i;
wire signed [`CalcTempBus]          temp_b3_28_15_r;
wire signed [`CalcTempBus]          temp_b3_28_15_i;
wire signed [`CalcTempBus]          temp_b3_28_16_r;
wire signed [`CalcTempBus]          temp_b3_28_16_i;
wire signed [`CalcTempBus]          temp_b3_28_17_r;
wire signed [`CalcTempBus]          temp_b3_28_17_i;
wire signed [`CalcTempBus]          temp_b3_28_18_r;
wire signed [`CalcTempBus]          temp_b3_28_18_i;
wire signed [`CalcTempBus]          temp_b3_28_19_r;
wire signed [`CalcTempBus]          temp_b3_28_19_i;
wire signed [`CalcTempBus]          temp_b3_28_20_r;
wire signed [`CalcTempBus]          temp_b3_28_20_i;
wire signed [`CalcTempBus]          temp_b3_28_21_r;
wire signed [`CalcTempBus]          temp_b3_28_21_i;
wire signed [`CalcTempBus]          temp_b3_28_22_r;
wire signed [`CalcTempBus]          temp_b3_28_22_i;
wire signed [`CalcTempBus]          temp_b3_28_23_r;
wire signed [`CalcTempBus]          temp_b3_28_23_i;
wire signed [`CalcTempBus]          temp_b3_28_24_r;
wire signed [`CalcTempBus]          temp_b3_28_24_i;
wire signed [`CalcTempBus]          temp_b3_28_25_r;
wire signed [`CalcTempBus]          temp_b3_28_25_i;
wire signed [`CalcTempBus]          temp_b3_28_26_r;
wire signed [`CalcTempBus]          temp_b3_28_26_i;
wire signed [`CalcTempBus]          temp_b3_28_27_r;
wire signed [`CalcTempBus]          temp_b3_28_27_i;
wire signed [`CalcTempBus]          temp_b3_28_28_r;
wire signed [`CalcTempBus]          temp_b3_28_28_i;
wire signed [`CalcTempBus]          temp_b3_28_29_r;
wire signed [`CalcTempBus]          temp_b3_28_29_i;
wire signed [`CalcTempBus]          temp_b3_28_30_r;
wire signed [`CalcTempBus]          temp_b3_28_30_i;
wire signed [`CalcTempBus]          temp_b3_28_31_r;
wire signed [`CalcTempBus]          temp_b3_28_31_i;
wire signed [`CalcTempBus]          temp_b3_28_32_r;
wire signed [`CalcTempBus]          temp_b3_28_32_i;
wire signed [`CalcTempBus]          temp_b3_29_1_r;
wire signed [`CalcTempBus]          temp_b3_29_1_i;
wire signed [`CalcTempBus]          temp_b3_29_2_r;
wire signed [`CalcTempBus]          temp_b3_29_2_i;
wire signed [`CalcTempBus]          temp_b3_29_3_r;
wire signed [`CalcTempBus]          temp_b3_29_3_i;
wire signed [`CalcTempBus]          temp_b3_29_4_r;
wire signed [`CalcTempBus]          temp_b3_29_4_i;
wire signed [`CalcTempBus]          temp_b3_29_5_r;
wire signed [`CalcTempBus]          temp_b3_29_5_i;
wire signed [`CalcTempBus]          temp_b3_29_6_r;
wire signed [`CalcTempBus]          temp_b3_29_6_i;
wire signed [`CalcTempBus]          temp_b3_29_7_r;
wire signed [`CalcTempBus]          temp_b3_29_7_i;
wire signed [`CalcTempBus]          temp_b3_29_8_r;
wire signed [`CalcTempBus]          temp_b3_29_8_i;
wire signed [`CalcTempBus]          temp_b3_29_9_r;
wire signed [`CalcTempBus]          temp_b3_29_9_i;
wire signed [`CalcTempBus]          temp_b3_29_10_r;
wire signed [`CalcTempBus]          temp_b3_29_10_i;
wire signed [`CalcTempBus]          temp_b3_29_11_r;
wire signed [`CalcTempBus]          temp_b3_29_11_i;
wire signed [`CalcTempBus]          temp_b3_29_12_r;
wire signed [`CalcTempBus]          temp_b3_29_12_i;
wire signed [`CalcTempBus]          temp_b3_29_13_r;
wire signed [`CalcTempBus]          temp_b3_29_13_i;
wire signed [`CalcTempBus]          temp_b3_29_14_r;
wire signed [`CalcTempBus]          temp_b3_29_14_i;
wire signed [`CalcTempBus]          temp_b3_29_15_r;
wire signed [`CalcTempBus]          temp_b3_29_15_i;
wire signed [`CalcTempBus]          temp_b3_29_16_r;
wire signed [`CalcTempBus]          temp_b3_29_16_i;
wire signed [`CalcTempBus]          temp_b3_29_17_r;
wire signed [`CalcTempBus]          temp_b3_29_17_i;
wire signed [`CalcTempBus]          temp_b3_29_18_r;
wire signed [`CalcTempBus]          temp_b3_29_18_i;
wire signed [`CalcTempBus]          temp_b3_29_19_r;
wire signed [`CalcTempBus]          temp_b3_29_19_i;
wire signed [`CalcTempBus]          temp_b3_29_20_r;
wire signed [`CalcTempBus]          temp_b3_29_20_i;
wire signed [`CalcTempBus]          temp_b3_29_21_r;
wire signed [`CalcTempBus]          temp_b3_29_21_i;
wire signed [`CalcTempBus]          temp_b3_29_22_r;
wire signed [`CalcTempBus]          temp_b3_29_22_i;
wire signed [`CalcTempBus]          temp_b3_29_23_r;
wire signed [`CalcTempBus]          temp_b3_29_23_i;
wire signed [`CalcTempBus]          temp_b3_29_24_r;
wire signed [`CalcTempBus]          temp_b3_29_24_i;
wire signed [`CalcTempBus]          temp_b3_29_25_r;
wire signed [`CalcTempBus]          temp_b3_29_25_i;
wire signed [`CalcTempBus]          temp_b3_29_26_r;
wire signed [`CalcTempBus]          temp_b3_29_26_i;
wire signed [`CalcTempBus]          temp_b3_29_27_r;
wire signed [`CalcTempBus]          temp_b3_29_27_i;
wire signed [`CalcTempBus]          temp_b3_29_28_r;
wire signed [`CalcTempBus]          temp_b3_29_28_i;
wire signed [`CalcTempBus]          temp_b3_29_29_r;
wire signed [`CalcTempBus]          temp_b3_29_29_i;
wire signed [`CalcTempBus]          temp_b3_29_30_r;
wire signed [`CalcTempBus]          temp_b3_29_30_i;
wire signed [`CalcTempBus]          temp_b3_29_31_r;
wire signed [`CalcTempBus]          temp_b3_29_31_i;
wire signed [`CalcTempBus]          temp_b3_29_32_r;
wire signed [`CalcTempBus]          temp_b3_29_32_i;
wire signed [`CalcTempBus]          temp_b3_30_1_r;
wire signed [`CalcTempBus]          temp_b3_30_1_i;
wire signed [`CalcTempBus]          temp_b3_30_2_r;
wire signed [`CalcTempBus]          temp_b3_30_2_i;
wire signed [`CalcTempBus]          temp_b3_30_3_r;
wire signed [`CalcTempBus]          temp_b3_30_3_i;
wire signed [`CalcTempBus]          temp_b3_30_4_r;
wire signed [`CalcTempBus]          temp_b3_30_4_i;
wire signed [`CalcTempBus]          temp_b3_30_5_r;
wire signed [`CalcTempBus]          temp_b3_30_5_i;
wire signed [`CalcTempBus]          temp_b3_30_6_r;
wire signed [`CalcTempBus]          temp_b3_30_6_i;
wire signed [`CalcTempBus]          temp_b3_30_7_r;
wire signed [`CalcTempBus]          temp_b3_30_7_i;
wire signed [`CalcTempBus]          temp_b3_30_8_r;
wire signed [`CalcTempBus]          temp_b3_30_8_i;
wire signed [`CalcTempBus]          temp_b3_30_9_r;
wire signed [`CalcTempBus]          temp_b3_30_9_i;
wire signed [`CalcTempBus]          temp_b3_30_10_r;
wire signed [`CalcTempBus]          temp_b3_30_10_i;
wire signed [`CalcTempBus]          temp_b3_30_11_r;
wire signed [`CalcTempBus]          temp_b3_30_11_i;
wire signed [`CalcTempBus]          temp_b3_30_12_r;
wire signed [`CalcTempBus]          temp_b3_30_12_i;
wire signed [`CalcTempBus]          temp_b3_30_13_r;
wire signed [`CalcTempBus]          temp_b3_30_13_i;
wire signed [`CalcTempBus]          temp_b3_30_14_r;
wire signed [`CalcTempBus]          temp_b3_30_14_i;
wire signed [`CalcTempBus]          temp_b3_30_15_r;
wire signed [`CalcTempBus]          temp_b3_30_15_i;
wire signed [`CalcTempBus]          temp_b3_30_16_r;
wire signed [`CalcTempBus]          temp_b3_30_16_i;
wire signed [`CalcTempBus]          temp_b3_30_17_r;
wire signed [`CalcTempBus]          temp_b3_30_17_i;
wire signed [`CalcTempBus]          temp_b3_30_18_r;
wire signed [`CalcTempBus]          temp_b3_30_18_i;
wire signed [`CalcTempBus]          temp_b3_30_19_r;
wire signed [`CalcTempBus]          temp_b3_30_19_i;
wire signed [`CalcTempBus]          temp_b3_30_20_r;
wire signed [`CalcTempBus]          temp_b3_30_20_i;
wire signed [`CalcTempBus]          temp_b3_30_21_r;
wire signed [`CalcTempBus]          temp_b3_30_21_i;
wire signed [`CalcTempBus]          temp_b3_30_22_r;
wire signed [`CalcTempBus]          temp_b3_30_22_i;
wire signed [`CalcTempBus]          temp_b3_30_23_r;
wire signed [`CalcTempBus]          temp_b3_30_23_i;
wire signed [`CalcTempBus]          temp_b3_30_24_r;
wire signed [`CalcTempBus]          temp_b3_30_24_i;
wire signed [`CalcTempBus]          temp_b3_30_25_r;
wire signed [`CalcTempBus]          temp_b3_30_25_i;
wire signed [`CalcTempBus]          temp_b3_30_26_r;
wire signed [`CalcTempBus]          temp_b3_30_26_i;
wire signed [`CalcTempBus]          temp_b3_30_27_r;
wire signed [`CalcTempBus]          temp_b3_30_27_i;
wire signed [`CalcTempBus]          temp_b3_30_28_r;
wire signed [`CalcTempBus]          temp_b3_30_28_i;
wire signed [`CalcTempBus]          temp_b3_30_29_r;
wire signed [`CalcTempBus]          temp_b3_30_29_i;
wire signed [`CalcTempBus]          temp_b3_30_30_r;
wire signed [`CalcTempBus]          temp_b3_30_30_i;
wire signed [`CalcTempBus]          temp_b3_30_31_r;
wire signed [`CalcTempBus]          temp_b3_30_31_i;
wire signed [`CalcTempBus]          temp_b3_30_32_r;
wire signed [`CalcTempBus]          temp_b3_30_32_i;
wire signed [`CalcTempBus]          temp_b3_31_1_r;
wire signed [`CalcTempBus]          temp_b3_31_1_i;
wire signed [`CalcTempBus]          temp_b3_31_2_r;
wire signed [`CalcTempBus]          temp_b3_31_2_i;
wire signed [`CalcTempBus]          temp_b3_31_3_r;
wire signed [`CalcTempBus]          temp_b3_31_3_i;
wire signed [`CalcTempBus]          temp_b3_31_4_r;
wire signed [`CalcTempBus]          temp_b3_31_4_i;
wire signed [`CalcTempBus]          temp_b3_31_5_r;
wire signed [`CalcTempBus]          temp_b3_31_5_i;
wire signed [`CalcTempBus]          temp_b3_31_6_r;
wire signed [`CalcTempBus]          temp_b3_31_6_i;
wire signed [`CalcTempBus]          temp_b3_31_7_r;
wire signed [`CalcTempBus]          temp_b3_31_7_i;
wire signed [`CalcTempBus]          temp_b3_31_8_r;
wire signed [`CalcTempBus]          temp_b3_31_8_i;
wire signed [`CalcTempBus]          temp_b3_31_9_r;
wire signed [`CalcTempBus]          temp_b3_31_9_i;
wire signed [`CalcTempBus]          temp_b3_31_10_r;
wire signed [`CalcTempBus]          temp_b3_31_10_i;
wire signed [`CalcTempBus]          temp_b3_31_11_r;
wire signed [`CalcTempBus]          temp_b3_31_11_i;
wire signed [`CalcTempBus]          temp_b3_31_12_r;
wire signed [`CalcTempBus]          temp_b3_31_12_i;
wire signed [`CalcTempBus]          temp_b3_31_13_r;
wire signed [`CalcTempBus]          temp_b3_31_13_i;
wire signed [`CalcTempBus]          temp_b3_31_14_r;
wire signed [`CalcTempBus]          temp_b3_31_14_i;
wire signed [`CalcTempBus]          temp_b3_31_15_r;
wire signed [`CalcTempBus]          temp_b3_31_15_i;
wire signed [`CalcTempBus]          temp_b3_31_16_r;
wire signed [`CalcTempBus]          temp_b3_31_16_i;
wire signed [`CalcTempBus]          temp_b3_31_17_r;
wire signed [`CalcTempBus]          temp_b3_31_17_i;
wire signed [`CalcTempBus]          temp_b3_31_18_r;
wire signed [`CalcTempBus]          temp_b3_31_18_i;
wire signed [`CalcTempBus]          temp_b3_31_19_r;
wire signed [`CalcTempBus]          temp_b3_31_19_i;
wire signed [`CalcTempBus]          temp_b3_31_20_r;
wire signed [`CalcTempBus]          temp_b3_31_20_i;
wire signed [`CalcTempBus]          temp_b3_31_21_r;
wire signed [`CalcTempBus]          temp_b3_31_21_i;
wire signed [`CalcTempBus]          temp_b3_31_22_r;
wire signed [`CalcTempBus]          temp_b3_31_22_i;
wire signed [`CalcTempBus]          temp_b3_31_23_r;
wire signed [`CalcTempBus]          temp_b3_31_23_i;
wire signed [`CalcTempBus]          temp_b3_31_24_r;
wire signed [`CalcTempBus]          temp_b3_31_24_i;
wire signed [`CalcTempBus]          temp_b3_31_25_r;
wire signed [`CalcTempBus]          temp_b3_31_25_i;
wire signed [`CalcTempBus]          temp_b3_31_26_r;
wire signed [`CalcTempBus]          temp_b3_31_26_i;
wire signed [`CalcTempBus]          temp_b3_31_27_r;
wire signed [`CalcTempBus]          temp_b3_31_27_i;
wire signed [`CalcTempBus]          temp_b3_31_28_r;
wire signed [`CalcTempBus]          temp_b3_31_28_i;
wire signed [`CalcTempBus]          temp_b3_31_29_r;
wire signed [`CalcTempBus]          temp_b3_31_29_i;
wire signed [`CalcTempBus]          temp_b3_31_30_r;
wire signed [`CalcTempBus]          temp_b3_31_30_i;
wire signed [`CalcTempBus]          temp_b3_31_31_r;
wire signed [`CalcTempBus]          temp_b3_31_31_i;
wire signed [`CalcTempBus]          temp_b3_31_32_r;
wire signed [`CalcTempBus]          temp_b3_31_32_i;
wire signed [`CalcTempBus]          temp_b3_32_1_r;
wire signed [`CalcTempBus]          temp_b3_32_1_i;
wire signed [`CalcTempBus]          temp_b3_32_2_r;
wire signed [`CalcTempBus]          temp_b3_32_2_i;
wire signed [`CalcTempBus]          temp_b3_32_3_r;
wire signed [`CalcTempBus]          temp_b3_32_3_i;
wire signed [`CalcTempBus]          temp_b3_32_4_r;
wire signed [`CalcTempBus]          temp_b3_32_4_i;
wire signed [`CalcTempBus]          temp_b3_32_5_r;
wire signed [`CalcTempBus]          temp_b3_32_5_i;
wire signed [`CalcTempBus]          temp_b3_32_6_r;
wire signed [`CalcTempBus]          temp_b3_32_6_i;
wire signed [`CalcTempBus]          temp_b3_32_7_r;
wire signed [`CalcTempBus]          temp_b3_32_7_i;
wire signed [`CalcTempBus]          temp_b3_32_8_r;
wire signed [`CalcTempBus]          temp_b3_32_8_i;
wire signed [`CalcTempBus]          temp_b3_32_9_r;
wire signed [`CalcTempBus]          temp_b3_32_9_i;
wire signed [`CalcTempBus]          temp_b3_32_10_r;
wire signed [`CalcTempBus]          temp_b3_32_10_i;
wire signed [`CalcTempBus]          temp_b3_32_11_r;
wire signed [`CalcTempBus]          temp_b3_32_11_i;
wire signed [`CalcTempBus]          temp_b3_32_12_r;
wire signed [`CalcTempBus]          temp_b3_32_12_i;
wire signed [`CalcTempBus]          temp_b3_32_13_r;
wire signed [`CalcTempBus]          temp_b3_32_13_i;
wire signed [`CalcTempBus]          temp_b3_32_14_r;
wire signed [`CalcTempBus]          temp_b3_32_14_i;
wire signed [`CalcTempBus]          temp_b3_32_15_r;
wire signed [`CalcTempBus]          temp_b3_32_15_i;
wire signed [`CalcTempBus]          temp_b3_32_16_r;
wire signed [`CalcTempBus]          temp_b3_32_16_i;
wire signed [`CalcTempBus]          temp_b3_32_17_r;
wire signed [`CalcTempBus]          temp_b3_32_17_i;
wire signed [`CalcTempBus]          temp_b3_32_18_r;
wire signed [`CalcTempBus]          temp_b3_32_18_i;
wire signed [`CalcTempBus]          temp_b3_32_19_r;
wire signed [`CalcTempBus]          temp_b3_32_19_i;
wire signed [`CalcTempBus]          temp_b3_32_20_r;
wire signed [`CalcTempBus]          temp_b3_32_20_i;
wire signed [`CalcTempBus]          temp_b3_32_21_r;
wire signed [`CalcTempBus]          temp_b3_32_21_i;
wire signed [`CalcTempBus]          temp_b3_32_22_r;
wire signed [`CalcTempBus]          temp_b3_32_22_i;
wire signed [`CalcTempBus]          temp_b3_32_23_r;
wire signed [`CalcTempBus]          temp_b3_32_23_i;
wire signed [`CalcTempBus]          temp_b3_32_24_r;
wire signed [`CalcTempBus]          temp_b3_32_24_i;
wire signed [`CalcTempBus]          temp_b3_32_25_r;
wire signed [`CalcTempBus]          temp_b3_32_25_i;
wire signed [`CalcTempBus]          temp_b3_32_26_r;
wire signed [`CalcTempBus]          temp_b3_32_26_i;
wire signed [`CalcTempBus]          temp_b3_32_27_r;
wire signed [`CalcTempBus]          temp_b3_32_27_i;
wire signed [`CalcTempBus]          temp_b3_32_28_r;
wire signed [`CalcTempBus]          temp_b3_32_28_i;
wire signed [`CalcTempBus]          temp_b3_32_29_r;
wire signed [`CalcTempBus]          temp_b3_32_29_i;
wire signed [`CalcTempBus]          temp_b3_32_30_r;
wire signed [`CalcTempBus]          temp_b3_32_30_i;
wire signed [`CalcTempBus]          temp_b3_32_31_r;
wire signed [`CalcTempBus]          temp_b3_32_31_i;
wire signed [`CalcTempBus]          temp_b3_32_32_r;
wire signed [`CalcTempBus]          temp_b3_32_32_i;
wire signed [`CalcTempBus]          temp_b4_1_1_r;
wire signed [`CalcTempBus]          temp_b4_1_1_i;
wire signed [`CalcTempBus]          temp_b4_1_2_r;
wire signed [`CalcTempBus]          temp_b4_1_2_i;
wire signed [`CalcTempBus]          temp_b4_1_3_r;
wire signed [`CalcTempBus]          temp_b4_1_3_i;
wire signed [`CalcTempBus]          temp_b4_1_4_r;
wire signed [`CalcTempBus]          temp_b4_1_4_i;
wire signed [`CalcTempBus]          temp_b4_1_5_r;
wire signed [`CalcTempBus]          temp_b4_1_5_i;
wire signed [`CalcTempBus]          temp_b4_1_6_r;
wire signed [`CalcTempBus]          temp_b4_1_6_i;
wire signed [`CalcTempBus]          temp_b4_1_7_r;
wire signed [`CalcTempBus]          temp_b4_1_7_i;
wire signed [`CalcTempBus]          temp_b4_1_8_r;
wire signed [`CalcTempBus]          temp_b4_1_8_i;
wire signed [`CalcTempBus]          temp_b4_1_9_r;
wire signed [`CalcTempBus]          temp_b4_1_9_i;
wire signed [`CalcTempBus]          temp_b4_1_10_r;
wire signed [`CalcTempBus]          temp_b4_1_10_i;
wire signed [`CalcTempBus]          temp_b4_1_11_r;
wire signed [`CalcTempBus]          temp_b4_1_11_i;
wire signed [`CalcTempBus]          temp_b4_1_12_r;
wire signed [`CalcTempBus]          temp_b4_1_12_i;
wire signed [`CalcTempBus]          temp_b4_1_13_r;
wire signed [`CalcTempBus]          temp_b4_1_13_i;
wire signed [`CalcTempBus]          temp_b4_1_14_r;
wire signed [`CalcTempBus]          temp_b4_1_14_i;
wire signed [`CalcTempBus]          temp_b4_1_15_r;
wire signed [`CalcTempBus]          temp_b4_1_15_i;
wire signed [`CalcTempBus]          temp_b4_1_16_r;
wire signed [`CalcTempBus]          temp_b4_1_16_i;
wire signed [`CalcTempBus]          temp_b4_1_17_r;
wire signed [`CalcTempBus]          temp_b4_1_17_i;
wire signed [`CalcTempBus]          temp_b4_1_18_r;
wire signed [`CalcTempBus]          temp_b4_1_18_i;
wire signed [`CalcTempBus]          temp_b4_1_19_r;
wire signed [`CalcTempBus]          temp_b4_1_19_i;
wire signed [`CalcTempBus]          temp_b4_1_20_r;
wire signed [`CalcTempBus]          temp_b4_1_20_i;
wire signed [`CalcTempBus]          temp_b4_1_21_r;
wire signed [`CalcTempBus]          temp_b4_1_21_i;
wire signed [`CalcTempBus]          temp_b4_1_22_r;
wire signed [`CalcTempBus]          temp_b4_1_22_i;
wire signed [`CalcTempBus]          temp_b4_1_23_r;
wire signed [`CalcTempBus]          temp_b4_1_23_i;
wire signed [`CalcTempBus]          temp_b4_1_24_r;
wire signed [`CalcTempBus]          temp_b4_1_24_i;
wire signed [`CalcTempBus]          temp_b4_1_25_r;
wire signed [`CalcTempBus]          temp_b4_1_25_i;
wire signed [`CalcTempBus]          temp_b4_1_26_r;
wire signed [`CalcTempBus]          temp_b4_1_26_i;
wire signed [`CalcTempBus]          temp_b4_1_27_r;
wire signed [`CalcTempBus]          temp_b4_1_27_i;
wire signed [`CalcTempBus]          temp_b4_1_28_r;
wire signed [`CalcTempBus]          temp_b4_1_28_i;
wire signed [`CalcTempBus]          temp_b4_1_29_r;
wire signed [`CalcTempBus]          temp_b4_1_29_i;
wire signed [`CalcTempBus]          temp_b4_1_30_r;
wire signed [`CalcTempBus]          temp_b4_1_30_i;
wire signed [`CalcTempBus]          temp_b4_1_31_r;
wire signed [`CalcTempBus]          temp_b4_1_31_i;
wire signed [`CalcTempBus]          temp_b4_1_32_r;
wire signed [`CalcTempBus]          temp_b4_1_32_i;
wire signed [`CalcTempBus]          temp_b4_2_1_r;
wire signed [`CalcTempBus]          temp_b4_2_1_i;
wire signed [`CalcTempBus]          temp_b4_2_2_r;
wire signed [`CalcTempBus]          temp_b4_2_2_i;
wire signed [`CalcTempBus]          temp_b4_2_3_r;
wire signed [`CalcTempBus]          temp_b4_2_3_i;
wire signed [`CalcTempBus]          temp_b4_2_4_r;
wire signed [`CalcTempBus]          temp_b4_2_4_i;
wire signed [`CalcTempBus]          temp_b4_2_5_r;
wire signed [`CalcTempBus]          temp_b4_2_5_i;
wire signed [`CalcTempBus]          temp_b4_2_6_r;
wire signed [`CalcTempBus]          temp_b4_2_6_i;
wire signed [`CalcTempBus]          temp_b4_2_7_r;
wire signed [`CalcTempBus]          temp_b4_2_7_i;
wire signed [`CalcTempBus]          temp_b4_2_8_r;
wire signed [`CalcTempBus]          temp_b4_2_8_i;
wire signed [`CalcTempBus]          temp_b4_2_9_r;
wire signed [`CalcTempBus]          temp_b4_2_9_i;
wire signed [`CalcTempBus]          temp_b4_2_10_r;
wire signed [`CalcTempBus]          temp_b4_2_10_i;
wire signed [`CalcTempBus]          temp_b4_2_11_r;
wire signed [`CalcTempBus]          temp_b4_2_11_i;
wire signed [`CalcTempBus]          temp_b4_2_12_r;
wire signed [`CalcTempBus]          temp_b4_2_12_i;
wire signed [`CalcTempBus]          temp_b4_2_13_r;
wire signed [`CalcTempBus]          temp_b4_2_13_i;
wire signed [`CalcTempBus]          temp_b4_2_14_r;
wire signed [`CalcTempBus]          temp_b4_2_14_i;
wire signed [`CalcTempBus]          temp_b4_2_15_r;
wire signed [`CalcTempBus]          temp_b4_2_15_i;
wire signed [`CalcTempBus]          temp_b4_2_16_r;
wire signed [`CalcTempBus]          temp_b4_2_16_i;
wire signed [`CalcTempBus]          temp_b4_2_17_r;
wire signed [`CalcTempBus]          temp_b4_2_17_i;
wire signed [`CalcTempBus]          temp_b4_2_18_r;
wire signed [`CalcTempBus]          temp_b4_2_18_i;
wire signed [`CalcTempBus]          temp_b4_2_19_r;
wire signed [`CalcTempBus]          temp_b4_2_19_i;
wire signed [`CalcTempBus]          temp_b4_2_20_r;
wire signed [`CalcTempBus]          temp_b4_2_20_i;
wire signed [`CalcTempBus]          temp_b4_2_21_r;
wire signed [`CalcTempBus]          temp_b4_2_21_i;
wire signed [`CalcTempBus]          temp_b4_2_22_r;
wire signed [`CalcTempBus]          temp_b4_2_22_i;
wire signed [`CalcTempBus]          temp_b4_2_23_r;
wire signed [`CalcTempBus]          temp_b4_2_23_i;
wire signed [`CalcTempBus]          temp_b4_2_24_r;
wire signed [`CalcTempBus]          temp_b4_2_24_i;
wire signed [`CalcTempBus]          temp_b4_2_25_r;
wire signed [`CalcTempBus]          temp_b4_2_25_i;
wire signed [`CalcTempBus]          temp_b4_2_26_r;
wire signed [`CalcTempBus]          temp_b4_2_26_i;
wire signed [`CalcTempBus]          temp_b4_2_27_r;
wire signed [`CalcTempBus]          temp_b4_2_27_i;
wire signed [`CalcTempBus]          temp_b4_2_28_r;
wire signed [`CalcTempBus]          temp_b4_2_28_i;
wire signed [`CalcTempBus]          temp_b4_2_29_r;
wire signed [`CalcTempBus]          temp_b4_2_29_i;
wire signed [`CalcTempBus]          temp_b4_2_30_r;
wire signed [`CalcTempBus]          temp_b4_2_30_i;
wire signed [`CalcTempBus]          temp_b4_2_31_r;
wire signed [`CalcTempBus]          temp_b4_2_31_i;
wire signed [`CalcTempBus]          temp_b4_2_32_r;
wire signed [`CalcTempBus]          temp_b4_2_32_i;
wire signed [`CalcTempBus]          temp_b4_3_1_r;
wire signed [`CalcTempBus]          temp_b4_3_1_i;
wire signed [`CalcTempBus]          temp_b4_3_2_r;
wire signed [`CalcTempBus]          temp_b4_3_2_i;
wire signed [`CalcTempBus]          temp_b4_3_3_r;
wire signed [`CalcTempBus]          temp_b4_3_3_i;
wire signed [`CalcTempBus]          temp_b4_3_4_r;
wire signed [`CalcTempBus]          temp_b4_3_4_i;
wire signed [`CalcTempBus]          temp_b4_3_5_r;
wire signed [`CalcTempBus]          temp_b4_3_5_i;
wire signed [`CalcTempBus]          temp_b4_3_6_r;
wire signed [`CalcTempBus]          temp_b4_3_6_i;
wire signed [`CalcTempBus]          temp_b4_3_7_r;
wire signed [`CalcTempBus]          temp_b4_3_7_i;
wire signed [`CalcTempBus]          temp_b4_3_8_r;
wire signed [`CalcTempBus]          temp_b4_3_8_i;
wire signed [`CalcTempBus]          temp_b4_3_9_r;
wire signed [`CalcTempBus]          temp_b4_3_9_i;
wire signed [`CalcTempBus]          temp_b4_3_10_r;
wire signed [`CalcTempBus]          temp_b4_3_10_i;
wire signed [`CalcTempBus]          temp_b4_3_11_r;
wire signed [`CalcTempBus]          temp_b4_3_11_i;
wire signed [`CalcTempBus]          temp_b4_3_12_r;
wire signed [`CalcTempBus]          temp_b4_3_12_i;
wire signed [`CalcTempBus]          temp_b4_3_13_r;
wire signed [`CalcTempBus]          temp_b4_3_13_i;
wire signed [`CalcTempBus]          temp_b4_3_14_r;
wire signed [`CalcTempBus]          temp_b4_3_14_i;
wire signed [`CalcTempBus]          temp_b4_3_15_r;
wire signed [`CalcTempBus]          temp_b4_3_15_i;
wire signed [`CalcTempBus]          temp_b4_3_16_r;
wire signed [`CalcTempBus]          temp_b4_3_16_i;
wire signed [`CalcTempBus]          temp_b4_3_17_r;
wire signed [`CalcTempBus]          temp_b4_3_17_i;
wire signed [`CalcTempBus]          temp_b4_3_18_r;
wire signed [`CalcTempBus]          temp_b4_3_18_i;
wire signed [`CalcTempBus]          temp_b4_3_19_r;
wire signed [`CalcTempBus]          temp_b4_3_19_i;
wire signed [`CalcTempBus]          temp_b4_3_20_r;
wire signed [`CalcTempBus]          temp_b4_3_20_i;
wire signed [`CalcTempBus]          temp_b4_3_21_r;
wire signed [`CalcTempBus]          temp_b4_3_21_i;
wire signed [`CalcTempBus]          temp_b4_3_22_r;
wire signed [`CalcTempBus]          temp_b4_3_22_i;
wire signed [`CalcTempBus]          temp_b4_3_23_r;
wire signed [`CalcTempBus]          temp_b4_3_23_i;
wire signed [`CalcTempBus]          temp_b4_3_24_r;
wire signed [`CalcTempBus]          temp_b4_3_24_i;
wire signed [`CalcTempBus]          temp_b4_3_25_r;
wire signed [`CalcTempBus]          temp_b4_3_25_i;
wire signed [`CalcTempBus]          temp_b4_3_26_r;
wire signed [`CalcTempBus]          temp_b4_3_26_i;
wire signed [`CalcTempBus]          temp_b4_3_27_r;
wire signed [`CalcTempBus]          temp_b4_3_27_i;
wire signed [`CalcTempBus]          temp_b4_3_28_r;
wire signed [`CalcTempBus]          temp_b4_3_28_i;
wire signed [`CalcTempBus]          temp_b4_3_29_r;
wire signed [`CalcTempBus]          temp_b4_3_29_i;
wire signed [`CalcTempBus]          temp_b4_3_30_r;
wire signed [`CalcTempBus]          temp_b4_3_30_i;
wire signed [`CalcTempBus]          temp_b4_3_31_r;
wire signed [`CalcTempBus]          temp_b4_3_31_i;
wire signed [`CalcTempBus]          temp_b4_3_32_r;
wire signed [`CalcTempBus]          temp_b4_3_32_i;
wire signed [`CalcTempBus]          temp_b4_4_1_r;
wire signed [`CalcTempBus]          temp_b4_4_1_i;
wire signed [`CalcTempBus]          temp_b4_4_2_r;
wire signed [`CalcTempBus]          temp_b4_4_2_i;
wire signed [`CalcTempBus]          temp_b4_4_3_r;
wire signed [`CalcTempBus]          temp_b4_4_3_i;
wire signed [`CalcTempBus]          temp_b4_4_4_r;
wire signed [`CalcTempBus]          temp_b4_4_4_i;
wire signed [`CalcTempBus]          temp_b4_4_5_r;
wire signed [`CalcTempBus]          temp_b4_4_5_i;
wire signed [`CalcTempBus]          temp_b4_4_6_r;
wire signed [`CalcTempBus]          temp_b4_4_6_i;
wire signed [`CalcTempBus]          temp_b4_4_7_r;
wire signed [`CalcTempBus]          temp_b4_4_7_i;
wire signed [`CalcTempBus]          temp_b4_4_8_r;
wire signed [`CalcTempBus]          temp_b4_4_8_i;
wire signed [`CalcTempBus]          temp_b4_4_9_r;
wire signed [`CalcTempBus]          temp_b4_4_9_i;
wire signed [`CalcTempBus]          temp_b4_4_10_r;
wire signed [`CalcTempBus]          temp_b4_4_10_i;
wire signed [`CalcTempBus]          temp_b4_4_11_r;
wire signed [`CalcTempBus]          temp_b4_4_11_i;
wire signed [`CalcTempBus]          temp_b4_4_12_r;
wire signed [`CalcTempBus]          temp_b4_4_12_i;
wire signed [`CalcTempBus]          temp_b4_4_13_r;
wire signed [`CalcTempBus]          temp_b4_4_13_i;
wire signed [`CalcTempBus]          temp_b4_4_14_r;
wire signed [`CalcTempBus]          temp_b4_4_14_i;
wire signed [`CalcTempBus]          temp_b4_4_15_r;
wire signed [`CalcTempBus]          temp_b4_4_15_i;
wire signed [`CalcTempBus]          temp_b4_4_16_r;
wire signed [`CalcTempBus]          temp_b4_4_16_i;
wire signed [`CalcTempBus]          temp_b4_4_17_r;
wire signed [`CalcTempBus]          temp_b4_4_17_i;
wire signed [`CalcTempBus]          temp_b4_4_18_r;
wire signed [`CalcTempBus]          temp_b4_4_18_i;
wire signed [`CalcTempBus]          temp_b4_4_19_r;
wire signed [`CalcTempBus]          temp_b4_4_19_i;
wire signed [`CalcTempBus]          temp_b4_4_20_r;
wire signed [`CalcTempBus]          temp_b4_4_20_i;
wire signed [`CalcTempBus]          temp_b4_4_21_r;
wire signed [`CalcTempBus]          temp_b4_4_21_i;
wire signed [`CalcTempBus]          temp_b4_4_22_r;
wire signed [`CalcTempBus]          temp_b4_4_22_i;
wire signed [`CalcTempBus]          temp_b4_4_23_r;
wire signed [`CalcTempBus]          temp_b4_4_23_i;
wire signed [`CalcTempBus]          temp_b4_4_24_r;
wire signed [`CalcTempBus]          temp_b4_4_24_i;
wire signed [`CalcTempBus]          temp_b4_4_25_r;
wire signed [`CalcTempBus]          temp_b4_4_25_i;
wire signed [`CalcTempBus]          temp_b4_4_26_r;
wire signed [`CalcTempBus]          temp_b4_4_26_i;
wire signed [`CalcTempBus]          temp_b4_4_27_r;
wire signed [`CalcTempBus]          temp_b4_4_27_i;
wire signed [`CalcTempBus]          temp_b4_4_28_r;
wire signed [`CalcTempBus]          temp_b4_4_28_i;
wire signed [`CalcTempBus]          temp_b4_4_29_r;
wire signed [`CalcTempBus]          temp_b4_4_29_i;
wire signed [`CalcTempBus]          temp_b4_4_30_r;
wire signed [`CalcTempBus]          temp_b4_4_30_i;
wire signed [`CalcTempBus]          temp_b4_4_31_r;
wire signed [`CalcTempBus]          temp_b4_4_31_i;
wire signed [`CalcTempBus]          temp_b4_4_32_r;
wire signed [`CalcTempBus]          temp_b4_4_32_i;
wire signed [`CalcTempBus]          temp_b4_5_1_r;
wire signed [`CalcTempBus]          temp_b4_5_1_i;
wire signed [`CalcTempBus]          temp_b4_5_2_r;
wire signed [`CalcTempBus]          temp_b4_5_2_i;
wire signed [`CalcTempBus]          temp_b4_5_3_r;
wire signed [`CalcTempBus]          temp_b4_5_3_i;
wire signed [`CalcTempBus]          temp_b4_5_4_r;
wire signed [`CalcTempBus]          temp_b4_5_4_i;
wire signed [`CalcTempBus]          temp_b4_5_5_r;
wire signed [`CalcTempBus]          temp_b4_5_5_i;
wire signed [`CalcTempBus]          temp_b4_5_6_r;
wire signed [`CalcTempBus]          temp_b4_5_6_i;
wire signed [`CalcTempBus]          temp_b4_5_7_r;
wire signed [`CalcTempBus]          temp_b4_5_7_i;
wire signed [`CalcTempBus]          temp_b4_5_8_r;
wire signed [`CalcTempBus]          temp_b4_5_8_i;
wire signed [`CalcTempBus]          temp_b4_5_9_r;
wire signed [`CalcTempBus]          temp_b4_5_9_i;
wire signed [`CalcTempBus]          temp_b4_5_10_r;
wire signed [`CalcTempBus]          temp_b4_5_10_i;
wire signed [`CalcTempBus]          temp_b4_5_11_r;
wire signed [`CalcTempBus]          temp_b4_5_11_i;
wire signed [`CalcTempBus]          temp_b4_5_12_r;
wire signed [`CalcTempBus]          temp_b4_5_12_i;
wire signed [`CalcTempBus]          temp_b4_5_13_r;
wire signed [`CalcTempBus]          temp_b4_5_13_i;
wire signed [`CalcTempBus]          temp_b4_5_14_r;
wire signed [`CalcTempBus]          temp_b4_5_14_i;
wire signed [`CalcTempBus]          temp_b4_5_15_r;
wire signed [`CalcTempBus]          temp_b4_5_15_i;
wire signed [`CalcTempBus]          temp_b4_5_16_r;
wire signed [`CalcTempBus]          temp_b4_5_16_i;
wire signed [`CalcTempBus]          temp_b4_5_17_r;
wire signed [`CalcTempBus]          temp_b4_5_17_i;
wire signed [`CalcTempBus]          temp_b4_5_18_r;
wire signed [`CalcTempBus]          temp_b4_5_18_i;
wire signed [`CalcTempBus]          temp_b4_5_19_r;
wire signed [`CalcTempBus]          temp_b4_5_19_i;
wire signed [`CalcTempBus]          temp_b4_5_20_r;
wire signed [`CalcTempBus]          temp_b4_5_20_i;
wire signed [`CalcTempBus]          temp_b4_5_21_r;
wire signed [`CalcTempBus]          temp_b4_5_21_i;
wire signed [`CalcTempBus]          temp_b4_5_22_r;
wire signed [`CalcTempBus]          temp_b4_5_22_i;
wire signed [`CalcTempBus]          temp_b4_5_23_r;
wire signed [`CalcTempBus]          temp_b4_5_23_i;
wire signed [`CalcTempBus]          temp_b4_5_24_r;
wire signed [`CalcTempBus]          temp_b4_5_24_i;
wire signed [`CalcTempBus]          temp_b4_5_25_r;
wire signed [`CalcTempBus]          temp_b4_5_25_i;
wire signed [`CalcTempBus]          temp_b4_5_26_r;
wire signed [`CalcTempBus]          temp_b4_5_26_i;
wire signed [`CalcTempBus]          temp_b4_5_27_r;
wire signed [`CalcTempBus]          temp_b4_5_27_i;
wire signed [`CalcTempBus]          temp_b4_5_28_r;
wire signed [`CalcTempBus]          temp_b4_5_28_i;
wire signed [`CalcTempBus]          temp_b4_5_29_r;
wire signed [`CalcTempBus]          temp_b4_5_29_i;
wire signed [`CalcTempBus]          temp_b4_5_30_r;
wire signed [`CalcTempBus]          temp_b4_5_30_i;
wire signed [`CalcTempBus]          temp_b4_5_31_r;
wire signed [`CalcTempBus]          temp_b4_5_31_i;
wire signed [`CalcTempBus]          temp_b4_5_32_r;
wire signed [`CalcTempBus]          temp_b4_5_32_i;
wire signed [`CalcTempBus]          temp_b4_6_1_r;
wire signed [`CalcTempBus]          temp_b4_6_1_i;
wire signed [`CalcTempBus]          temp_b4_6_2_r;
wire signed [`CalcTempBus]          temp_b4_6_2_i;
wire signed [`CalcTempBus]          temp_b4_6_3_r;
wire signed [`CalcTempBus]          temp_b4_6_3_i;
wire signed [`CalcTempBus]          temp_b4_6_4_r;
wire signed [`CalcTempBus]          temp_b4_6_4_i;
wire signed [`CalcTempBus]          temp_b4_6_5_r;
wire signed [`CalcTempBus]          temp_b4_6_5_i;
wire signed [`CalcTempBus]          temp_b4_6_6_r;
wire signed [`CalcTempBus]          temp_b4_6_6_i;
wire signed [`CalcTempBus]          temp_b4_6_7_r;
wire signed [`CalcTempBus]          temp_b4_6_7_i;
wire signed [`CalcTempBus]          temp_b4_6_8_r;
wire signed [`CalcTempBus]          temp_b4_6_8_i;
wire signed [`CalcTempBus]          temp_b4_6_9_r;
wire signed [`CalcTempBus]          temp_b4_6_9_i;
wire signed [`CalcTempBus]          temp_b4_6_10_r;
wire signed [`CalcTempBus]          temp_b4_6_10_i;
wire signed [`CalcTempBus]          temp_b4_6_11_r;
wire signed [`CalcTempBus]          temp_b4_6_11_i;
wire signed [`CalcTempBus]          temp_b4_6_12_r;
wire signed [`CalcTempBus]          temp_b4_6_12_i;
wire signed [`CalcTempBus]          temp_b4_6_13_r;
wire signed [`CalcTempBus]          temp_b4_6_13_i;
wire signed [`CalcTempBus]          temp_b4_6_14_r;
wire signed [`CalcTempBus]          temp_b4_6_14_i;
wire signed [`CalcTempBus]          temp_b4_6_15_r;
wire signed [`CalcTempBus]          temp_b4_6_15_i;
wire signed [`CalcTempBus]          temp_b4_6_16_r;
wire signed [`CalcTempBus]          temp_b4_6_16_i;
wire signed [`CalcTempBus]          temp_b4_6_17_r;
wire signed [`CalcTempBus]          temp_b4_6_17_i;
wire signed [`CalcTempBus]          temp_b4_6_18_r;
wire signed [`CalcTempBus]          temp_b4_6_18_i;
wire signed [`CalcTempBus]          temp_b4_6_19_r;
wire signed [`CalcTempBus]          temp_b4_6_19_i;
wire signed [`CalcTempBus]          temp_b4_6_20_r;
wire signed [`CalcTempBus]          temp_b4_6_20_i;
wire signed [`CalcTempBus]          temp_b4_6_21_r;
wire signed [`CalcTempBus]          temp_b4_6_21_i;
wire signed [`CalcTempBus]          temp_b4_6_22_r;
wire signed [`CalcTempBus]          temp_b4_6_22_i;
wire signed [`CalcTempBus]          temp_b4_6_23_r;
wire signed [`CalcTempBus]          temp_b4_6_23_i;
wire signed [`CalcTempBus]          temp_b4_6_24_r;
wire signed [`CalcTempBus]          temp_b4_6_24_i;
wire signed [`CalcTempBus]          temp_b4_6_25_r;
wire signed [`CalcTempBus]          temp_b4_6_25_i;
wire signed [`CalcTempBus]          temp_b4_6_26_r;
wire signed [`CalcTempBus]          temp_b4_6_26_i;
wire signed [`CalcTempBus]          temp_b4_6_27_r;
wire signed [`CalcTempBus]          temp_b4_6_27_i;
wire signed [`CalcTempBus]          temp_b4_6_28_r;
wire signed [`CalcTempBus]          temp_b4_6_28_i;
wire signed [`CalcTempBus]          temp_b4_6_29_r;
wire signed [`CalcTempBus]          temp_b4_6_29_i;
wire signed [`CalcTempBus]          temp_b4_6_30_r;
wire signed [`CalcTempBus]          temp_b4_6_30_i;
wire signed [`CalcTempBus]          temp_b4_6_31_r;
wire signed [`CalcTempBus]          temp_b4_6_31_i;
wire signed [`CalcTempBus]          temp_b4_6_32_r;
wire signed [`CalcTempBus]          temp_b4_6_32_i;
wire signed [`CalcTempBus]          temp_b4_7_1_r;
wire signed [`CalcTempBus]          temp_b4_7_1_i;
wire signed [`CalcTempBus]          temp_b4_7_2_r;
wire signed [`CalcTempBus]          temp_b4_7_2_i;
wire signed [`CalcTempBus]          temp_b4_7_3_r;
wire signed [`CalcTempBus]          temp_b4_7_3_i;
wire signed [`CalcTempBus]          temp_b4_7_4_r;
wire signed [`CalcTempBus]          temp_b4_7_4_i;
wire signed [`CalcTempBus]          temp_b4_7_5_r;
wire signed [`CalcTempBus]          temp_b4_7_5_i;
wire signed [`CalcTempBus]          temp_b4_7_6_r;
wire signed [`CalcTempBus]          temp_b4_7_6_i;
wire signed [`CalcTempBus]          temp_b4_7_7_r;
wire signed [`CalcTempBus]          temp_b4_7_7_i;
wire signed [`CalcTempBus]          temp_b4_7_8_r;
wire signed [`CalcTempBus]          temp_b4_7_8_i;
wire signed [`CalcTempBus]          temp_b4_7_9_r;
wire signed [`CalcTempBus]          temp_b4_7_9_i;
wire signed [`CalcTempBus]          temp_b4_7_10_r;
wire signed [`CalcTempBus]          temp_b4_7_10_i;
wire signed [`CalcTempBus]          temp_b4_7_11_r;
wire signed [`CalcTempBus]          temp_b4_7_11_i;
wire signed [`CalcTempBus]          temp_b4_7_12_r;
wire signed [`CalcTempBus]          temp_b4_7_12_i;
wire signed [`CalcTempBus]          temp_b4_7_13_r;
wire signed [`CalcTempBus]          temp_b4_7_13_i;
wire signed [`CalcTempBus]          temp_b4_7_14_r;
wire signed [`CalcTempBus]          temp_b4_7_14_i;
wire signed [`CalcTempBus]          temp_b4_7_15_r;
wire signed [`CalcTempBus]          temp_b4_7_15_i;
wire signed [`CalcTempBus]          temp_b4_7_16_r;
wire signed [`CalcTempBus]          temp_b4_7_16_i;
wire signed [`CalcTempBus]          temp_b4_7_17_r;
wire signed [`CalcTempBus]          temp_b4_7_17_i;
wire signed [`CalcTempBus]          temp_b4_7_18_r;
wire signed [`CalcTempBus]          temp_b4_7_18_i;
wire signed [`CalcTempBus]          temp_b4_7_19_r;
wire signed [`CalcTempBus]          temp_b4_7_19_i;
wire signed [`CalcTempBus]          temp_b4_7_20_r;
wire signed [`CalcTempBus]          temp_b4_7_20_i;
wire signed [`CalcTempBus]          temp_b4_7_21_r;
wire signed [`CalcTempBus]          temp_b4_7_21_i;
wire signed [`CalcTempBus]          temp_b4_7_22_r;
wire signed [`CalcTempBus]          temp_b4_7_22_i;
wire signed [`CalcTempBus]          temp_b4_7_23_r;
wire signed [`CalcTempBus]          temp_b4_7_23_i;
wire signed [`CalcTempBus]          temp_b4_7_24_r;
wire signed [`CalcTempBus]          temp_b4_7_24_i;
wire signed [`CalcTempBus]          temp_b4_7_25_r;
wire signed [`CalcTempBus]          temp_b4_7_25_i;
wire signed [`CalcTempBus]          temp_b4_7_26_r;
wire signed [`CalcTempBus]          temp_b4_7_26_i;
wire signed [`CalcTempBus]          temp_b4_7_27_r;
wire signed [`CalcTempBus]          temp_b4_7_27_i;
wire signed [`CalcTempBus]          temp_b4_7_28_r;
wire signed [`CalcTempBus]          temp_b4_7_28_i;
wire signed [`CalcTempBus]          temp_b4_7_29_r;
wire signed [`CalcTempBus]          temp_b4_7_29_i;
wire signed [`CalcTempBus]          temp_b4_7_30_r;
wire signed [`CalcTempBus]          temp_b4_7_30_i;
wire signed [`CalcTempBus]          temp_b4_7_31_r;
wire signed [`CalcTempBus]          temp_b4_7_31_i;
wire signed [`CalcTempBus]          temp_b4_7_32_r;
wire signed [`CalcTempBus]          temp_b4_7_32_i;
wire signed [`CalcTempBus]          temp_b4_8_1_r;
wire signed [`CalcTempBus]          temp_b4_8_1_i;
wire signed [`CalcTempBus]          temp_b4_8_2_r;
wire signed [`CalcTempBus]          temp_b4_8_2_i;
wire signed [`CalcTempBus]          temp_b4_8_3_r;
wire signed [`CalcTempBus]          temp_b4_8_3_i;
wire signed [`CalcTempBus]          temp_b4_8_4_r;
wire signed [`CalcTempBus]          temp_b4_8_4_i;
wire signed [`CalcTempBus]          temp_b4_8_5_r;
wire signed [`CalcTempBus]          temp_b4_8_5_i;
wire signed [`CalcTempBus]          temp_b4_8_6_r;
wire signed [`CalcTempBus]          temp_b4_8_6_i;
wire signed [`CalcTempBus]          temp_b4_8_7_r;
wire signed [`CalcTempBus]          temp_b4_8_7_i;
wire signed [`CalcTempBus]          temp_b4_8_8_r;
wire signed [`CalcTempBus]          temp_b4_8_8_i;
wire signed [`CalcTempBus]          temp_b4_8_9_r;
wire signed [`CalcTempBus]          temp_b4_8_9_i;
wire signed [`CalcTempBus]          temp_b4_8_10_r;
wire signed [`CalcTempBus]          temp_b4_8_10_i;
wire signed [`CalcTempBus]          temp_b4_8_11_r;
wire signed [`CalcTempBus]          temp_b4_8_11_i;
wire signed [`CalcTempBus]          temp_b4_8_12_r;
wire signed [`CalcTempBus]          temp_b4_8_12_i;
wire signed [`CalcTempBus]          temp_b4_8_13_r;
wire signed [`CalcTempBus]          temp_b4_8_13_i;
wire signed [`CalcTempBus]          temp_b4_8_14_r;
wire signed [`CalcTempBus]          temp_b4_8_14_i;
wire signed [`CalcTempBus]          temp_b4_8_15_r;
wire signed [`CalcTempBus]          temp_b4_8_15_i;
wire signed [`CalcTempBus]          temp_b4_8_16_r;
wire signed [`CalcTempBus]          temp_b4_8_16_i;
wire signed [`CalcTempBus]          temp_b4_8_17_r;
wire signed [`CalcTempBus]          temp_b4_8_17_i;
wire signed [`CalcTempBus]          temp_b4_8_18_r;
wire signed [`CalcTempBus]          temp_b4_8_18_i;
wire signed [`CalcTempBus]          temp_b4_8_19_r;
wire signed [`CalcTempBus]          temp_b4_8_19_i;
wire signed [`CalcTempBus]          temp_b4_8_20_r;
wire signed [`CalcTempBus]          temp_b4_8_20_i;
wire signed [`CalcTempBus]          temp_b4_8_21_r;
wire signed [`CalcTempBus]          temp_b4_8_21_i;
wire signed [`CalcTempBus]          temp_b4_8_22_r;
wire signed [`CalcTempBus]          temp_b4_8_22_i;
wire signed [`CalcTempBus]          temp_b4_8_23_r;
wire signed [`CalcTempBus]          temp_b4_8_23_i;
wire signed [`CalcTempBus]          temp_b4_8_24_r;
wire signed [`CalcTempBus]          temp_b4_8_24_i;
wire signed [`CalcTempBus]          temp_b4_8_25_r;
wire signed [`CalcTempBus]          temp_b4_8_25_i;
wire signed [`CalcTempBus]          temp_b4_8_26_r;
wire signed [`CalcTempBus]          temp_b4_8_26_i;
wire signed [`CalcTempBus]          temp_b4_8_27_r;
wire signed [`CalcTempBus]          temp_b4_8_27_i;
wire signed [`CalcTempBus]          temp_b4_8_28_r;
wire signed [`CalcTempBus]          temp_b4_8_28_i;
wire signed [`CalcTempBus]          temp_b4_8_29_r;
wire signed [`CalcTempBus]          temp_b4_8_29_i;
wire signed [`CalcTempBus]          temp_b4_8_30_r;
wire signed [`CalcTempBus]          temp_b4_8_30_i;
wire signed [`CalcTempBus]          temp_b4_8_31_r;
wire signed [`CalcTempBus]          temp_b4_8_31_i;
wire signed [`CalcTempBus]          temp_b4_8_32_r;
wire signed [`CalcTempBus]          temp_b4_8_32_i;
wire signed [`CalcTempBus]          temp_b4_9_1_r;
wire signed [`CalcTempBus]          temp_b4_9_1_i;
wire signed [`CalcTempBus]          temp_b4_9_2_r;
wire signed [`CalcTempBus]          temp_b4_9_2_i;
wire signed [`CalcTempBus]          temp_b4_9_3_r;
wire signed [`CalcTempBus]          temp_b4_9_3_i;
wire signed [`CalcTempBus]          temp_b4_9_4_r;
wire signed [`CalcTempBus]          temp_b4_9_4_i;
wire signed [`CalcTempBus]          temp_b4_9_5_r;
wire signed [`CalcTempBus]          temp_b4_9_5_i;
wire signed [`CalcTempBus]          temp_b4_9_6_r;
wire signed [`CalcTempBus]          temp_b4_9_6_i;
wire signed [`CalcTempBus]          temp_b4_9_7_r;
wire signed [`CalcTempBus]          temp_b4_9_7_i;
wire signed [`CalcTempBus]          temp_b4_9_8_r;
wire signed [`CalcTempBus]          temp_b4_9_8_i;
wire signed [`CalcTempBus]          temp_b4_9_9_r;
wire signed [`CalcTempBus]          temp_b4_9_9_i;
wire signed [`CalcTempBus]          temp_b4_9_10_r;
wire signed [`CalcTempBus]          temp_b4_9_10_i;
wire signed [`CalcTempBus]          temp_b4_9_11_r;
wire signed [`CalcTempBus]          temp_b4_9_11_i;
wire signed [`CalcTempBus]          temp_b4_9_12_r;
wire signed [`CalcTempBus]          temp_b4_9_12_i;
wire signed [`CalcTempBus]          temp_b4_9_13_r;
wire signed [`CalcTempBus]          temp_b4_9_13_i;
wire signed [`CalcTempBus]          temp_b4_9_14_r;
wire signed [`CalcTempBus]          temp_b4_9_14_i;
wire signed [`CalcTempBus]          temp_b4_9_15_r;
wire signed [`CalcTempBus]          temp_b4_9_15_i;
wire signed [`CalcTempBus]          temp_b4_9_16_r;
wire signed [`CalcTempBus]          temp_b4_9_16_i;
wire signed [`CalcTempBus]          temp_b4_9_17_r;
wire signed [`CalcTempBus]          temp_b4_9_17_i;
wire signed [`CalcTempBus]          temp_b4_9_18_r;
wire signed [`CalcTempBus]          temp_b4_9_18_i;
wire signed [`CalcTempBus]          temp_b4_9_19_r;
wire signed [`CalcTempBus]          temp_b4_9_19_i;
wire signed [`CalcTempBus]          temp_b4_9_20_r;
wire signed [`CalcTempBus]          temp_b4_9_20_i;
wire signed [`CalcTempBus]          temp_b4_9_21_r;
wire signed [`CalcTempBus]          temp_b4_9_21_i;
wire signed [`CalcTempBus]          temp_b4_9_22_r;
wire signed [`CalcTempBus]          temp_b4_9_22_i;
wire signed [`CalcTempBus]          temp_b4_9_23_r;
wire signed [`CalcTempBus]          temp_b4_9_23_i;
wire signed [`CalcTempBus]          temp_b4_9_24_r;
wire signed [`CalcTempBus]          temp_b4_9_24_i;
wire signed [`CalcTempBus]          temp_b4_9_25_r;
wire signed [`CalcTempBus]          temp_b4_9_25_i;
wire signed [`CalcTempBus]          temp_b4_9_26_r;
wire signed [`CalcTempBus]          temp_b4_9_26_i;
wire signed [`CalcTempBus]          temp_b4_9_27_r;
wire signed [`CalcTempBus]          temp_b4_9_27_i;
wire signed [`CalcTempBus]          temp_b4_9_28_r;
wire signed [`CalcTempBus]          temp_b4_9_28_i;
wire signed [`CalcTempBus]          temp_b4_9_29_r;
wire signed [`CalcTempBus]          temp_b4_9_29_i;
wire signed [`CalcTempBus]          temp_b4_9_30_r;
wire signed [`CalcTempBus]          temp_b4_9_30_i;
wire signed [`CalcTempBus]          temp_b4_9_31_r;
wire signed [`CalcTempBus]          temp_b4_9_31_i;
wire signed [`CalcTempBus]          temp_b4_9_32_r;
wire signed [`CalcTempBus]          temp_b4_9_32_i;
wire signed [`CalcTempBus]          temp_b4_10_1_r;
wire signed [`CalcTempBus]          temp_b4_10_1_i;
wire signed [`CalcTempBus]          temp_b4_10_2_r;
wire signed [`CalcTempBus]          temp_b4_10_2_i;
wire signed [`CalcTempBus]          temp_b4_10_3_r;
wire signed [`CalcTempBus]          temp_b4_10_3_i;
wire signed [`CalcTempBus]          temp_b4_10_4_r;
wire signed [`CalcTempBus]          temp_b4_10_4_i;
wire signed [`CalcTempBus]          temp_b4_10_5_r;
wire signed [`CalcTempBus]          temp_b4_10_5_i;
wire signed [`CalcTempBus]          temp_b4_10_6_r;
wire signed [`CalcTempBus]          temp_b4_10_6_i;
wire signed [`CalcTempBus]          temp_b4_10_7_r;
wire signed [`CalcTempBus]          temp_b4_10_7_i;
wire signed [`CalcTempBus]          temp_b4_10_8_r;
wire signed [`CalcTempBus]          temp_b4_10_8_i;
wire signed [`CalcTempBus]          temp_b4_10_9_r;
wire signed [`CalcTempBus]          temp_b4_10_9_i;
wire signed [`CalcTempBus]          temp_b4_10_10_r;
wire signed [`CalcTempBus]          temp_b4_10_10_i;
wire signed [`CalcTempBus]          temp_b4_10_11_r;
wire signed [`CalcTempBus]          temp_b4_10_11_i;
wire signed [`CalcTempBus]          temp_b4_10_12_r;
wire signed [`CalcTempBus]          temp_b4_10_12_i;
wire signed [`CalcTempBus]          temp_b4_10_13_r;
wire signed [`CalcTempBus]          temp_b4_10_13_i;
wire signed [`CalcTempBus]          temp_b4_10_14_r;
wire signed [`CalcTempBus]          temp_b4_10_14_i;
wire signed [`CalcTempBus]          temp_b4_10_15_r;
wire signed [`CalcTempBus]          temp_b4_10_15_i;
wire signed [`CalcTempBus]          temp_b4_10_16_r;
wire signed [`CalcTempBus]          temp_b4_10_16_i;
wire signed [`CalcTempBus]          temp_b4_10_17_r;
wire signed [`CalcTempBus]          temp_b4_10_17_i;
wire signed [`CalcTempBus]          temp_b4_10_18_r;
wire signed [`CalcTempBus]          temp_b4_10_18_i;
wire signed [`CalcTempBus]          temp_b4_10_19_r;
wire signed [`CalcTempBus]          temp_b4_10_19_i;
wire signed [`CalcTempBus]          temp_b4_10_20_r;
wire signed [`CalcTempBus]          temp_b4_10_20_i;
wire signed [`CalcTempBus]          temp_b4_10_21_r;
wire signed [`CalcTempBus]          temp_b4_10_21_i;
wire signed [`CalcTempBus]          temp_b4_10_22_r;
wire signed [`CalcTempBus]          temp_b4_10_22_i;
wire signed [`CalcTempBus]          temp_b4_10_23_r;
wire signed [`CalcTempBus]          temp_b4_10_23_i;
wire signed [`CalcTempBus]          temp_b4_10_24_r;
wire signed [`CalcTempBus]          temp_b4_10_24_i;
wire signed [`CalcTempBus]          temp_b4_10_25_r;
wire signed [`CalcTempBus]          temp_b4_10_25_i;
wire signed [`CalcTempBus]          temp_b4_10_26_r;
wire signed [`CalcTempBus]          temp_b4_10_26_i;
wire signed [`CalcTempBus]          temp_b4_10_27_r;
wire signed [`CalcTempBus]          temp_b4_10_27_i;
wire signed [`CalcTempBus]          temp_b4_10_28_r;
wire signed [`CalcTempBus]          temp_b4_10_28_i;
wire signed [`CalcTempBus]          temp_b4_10_29_r;
wire signed [`CalcTempBus]          temp_b4_10_29_i;
wire signed [`CalcTempBus]          temp_b4_10_30_r;
wire signed [`CalcTempBus]          temp_b4_10_30_i;
wire signed [`CalcTempBus]          temp_b4_10_31_r;
wire signed [`CalcTempBus]          temp_b4_10_31_i;
wire signed [`CalcTempBus]          temp_b4_10_32_r;
wire signed [`CalcTempBus]          temp_b4_10_32_i;
wire signed [`CalcTempBus]          temp_b4_11_1_r;
wire signed [`CalcTempBus]          temp_b4_11_1_i;
wire signed [`CalcTempBus]          temp_b4_11_2_r;
wire signed [`CalcTempBus]          temp_b4_11_2_i;
wire signed [`CalcTempBus]          temp_b4_11_3_r;
wire signed [`CalcTempBus]          temp_b4_11_3_i;
wire signed [`CalcTempBus]          temp_b4_11_4_r;
wire signed [`CalcTempBus]          temp_b4_11_4_i;
wire signed [`CalcTempBus]          temp_b4_11_5_r;
wire signed [`CalcTempBus]          temp_b4_11_5_i;
wire signed [`CalcTempBus]          temp_b4_11_6_r;
wire signed [`CalcTempBus]          temp_b4_11_6_i;
wire signed [`CalcTempBus]          temp_b4_11_7_r;
wire signed [`CalcTempBus]          temp_b4_11_7_i;
wire signed [`CalcTempBus]          temp_b4_11_8_r;
wire signed [`CalcTempBus]          temp_b4_11_8_i;
wire signed [`CalcTempBus]          temp_b4_11_9_r;
wire signed [`CalcTempBus]          temp_b4_11_9_i;
wire signed [`CalcTempBus]          temp_b4_11_10_r;
wire signed [`CalcTempBus]          temp_b4_11_10_i;
wire signed [`CalcTempBus]          temp_b4_11_11_r;
wire signed [`CalcTempBus]          temp_b4_11_11_i;
wire signed [`CalcTempBus]          temp_b4_11_12_r;
wire signed [`CalcTempBus]          temp_b4_11_12_i;
wire signed [`CalcTempBus]          temp_b4_11_13_r;
wire signed [`CalcTempBus]          temp_b4_11_13_i;
wire signed [`CalcTempBus]          temp_b4_11_14_r;
wire signed [`CalcTempBus]          temp_b4_11_14_i;
wire signed [`CalcTempBus]          temp_b4_11_15_r;
wire signed [`CalcTempBus]          temp_b4_11_15_i;
wire signed [`CalcTempBus]          temp_b4_11_16_r;
wire signed [`CalcTempBus]          temp_b4_11_16_i;
wire signed [`CalcTempBus]          temp_b4_11_17_r;
wire signed [`CalcTempBus]          temp_b4_11_17_i;
wire signed [`CalcTempBus]          temp_b4_11_18_r;
wire signed [`CalcTempBus]          temp_b4_11_18_i;
wire signed [`CalcTempBus]          temp_b4_11_19_r;
wire signed [`CalcTempBus]          temp_b4_11_19_i;
wire signed [`CalcTempBus]          temp_b4_11_20_r;
wire signed [`CalcTempBus]          temp_b4_11_20_i;
wire signed [`CalcTempBus]          temp_b4_11_21_r;
wire signed [`CalcTempBus]          temp_b4_11_21_i;
wire signed [`CalcTempBus]          temp_b4_11_22_r;
wire signed [`CalcTempBus]          temp_b4_11_22_i;
wire signed [`CalcTempBus]          temp_b4_11_23_r;
wire signed [`CalcTempBus]          temp_b4_11_23_i;
wire signed [`CalcTempBus]          temp_b4_11_24_r;
wire signed [`CalcTempBus]          temp_b4_11_24_i;
wire signed [`CalcTempBus]          temp_b4_11_25_r;
wire signed [`CalcTempBus]          temp_b4_11_25_i;
wire signed [`CalcTempBus]          temp_b4_11_26_r;
wire signed [`CalcTempBus]          temp_b4_11_26_i;
wire signed [`CalcTempBus]          temp_b4_11_27_r;
wire signed [`CalcTempBus]          temp_b4_11_27_i;
wire signed [`CalcTempBus]          temp_b4_11_28_r;
wire signed [`CalcTempBus]          temp_b4_11_28_i;
wire signed [`CalcTempBus]          temp_b4_11_29_r;
wire signed [`CalcTempBus]          temp_b4_11_29_i;
wire signed [`CalcTempBus]          temp_b4_11_30_r;
wire signed [`CalcTempBus]          temp_b4_11_30_i;
wire signed [`CalcTempBus]          temp_b4_11_31_r;
wire signed [`CalcTempBus]          temp_b4_11_31_i;
wire signed [`CalcTempBus]          temp_b4_11_32_r;
wire signed [`CalcTempBus]          temp_b4_11_32_i;
wire signed [`CalcTempBus]          temp_b4_12_1_r;
wire signed [`CalcTempBus]          temp_b4_12_1_i;
wire signed [`CalcTempBus]          temp_b4_12_2_r;
wire signed [`CalcTempBus]          temp_b4_12_2_i;
wire signed [`CalcTempBus]          temp_b4_12_3_r;
wire signed [`CalcTempBus]          temp_b4_12_3_i;
wire signed [`CalcTempBus]          temp_b4_12_4_r;
wire signed [`CalcTempBus]          temp_b4_12_4_i;
wire signed [`CalcTempBus]          temp_b4_12_5_r;
wire signed [`CalcTempBus]          temp_b4_12_5_i;
wire signed [`CalcTempBus]          temp_b4_12_6_r;
wire signed [`CalcTempBus]          temp_b4_12_6_i;
wire signed [`CalcTempBus]          temp_b4_12_7_r;
wire signed [`CalcTempBus]          temp_b4_12_7_i;
wire signed [`CalcTempBus]          temp_b4_12_8_r;
wire signed [`CalcTempBus]          temp_b4_12_8_i;
wire signed [`CalcTempBus]          temp_b4_12_9_r;
wire signed [`CalcTempBus]          temp_b4_12_9_i;
wire signed [`CalcTempBus]          temp_b4_12_10_r;
wire signed [`CalcTempBus]          temp_b4_12_10_i;
wire signed [`CalcTempBus]          temp_b4_12_11_r;
wire signed [`CalcTempBus]          temp_b4_12_11_i;
wire signed [`CalcTempBus]          temp_b4_12_12_r;
wire signed [`CalcTempBus]          temp_b4_12_12_i;
wire signed [`CalcTempBus]          temp_b4_12_13_r;
wire signed [`CalcTempBus]          temp_b4_12_13_i;
wire signed [`CalcTempBus]          temp_b4_12_14_r;
wire signed [`CalcTempBus]          temp_b4_12_14_i;
wire signed [`CalcTempBus]          temp_b4_12_15_r;
wire signed [`CalcTempBus]          temp_b4_12_15_i;
wire signed [`CalcTempBus]          temp_b4_12_16_r;
wire signed [`CalcTempBus]          temp_b4_12_16_i;
wire signed [`CalcTempBus]          temp_b4_12_17_r;
wire signed [`CalcTempBus]          temp_b4_12_17_i;
wire signed [`CalcTempBus]          temp_b4_12_18_r;
wire signed [`CalcTempBus]          temp_b4_12_18_i;
wire signed [`CalcTempBus]          temp_b4_12_19_r;
wire signed [`CalcTempBus]          temp_b4_12_19_i;
wire signed [`CalcTempBus]          temp_b4_12_20_r;
wire signed [`CalcTempBus]          temp_b4_12_20_i;
wire signed [`CalcTempBus]          temp_b4_12_21_r;
wire signed [`CalcTempBus]          temp_b4_12_21_i;
wire signed [`CalcTempBus]          temp_b4_12_22_r;
wire signed [`CalcTempBus]          temp_b4_12_22_i;
wire signed [`CalcTempBus]          temp_b4_12_23_r;
wire signed [`CalcTempBus]          temp_b4_12_23_i;
wire signed [`CalcTempBus]          temp_b4_12_24_r;
wire signed [`CalcTempBus]          temp_b4_12_24_i;
wire signed [`CalcTempBus]          temp_b4_12_25_r;
wire signed [`CalcTempBus]          temp_b4_12_25_i;
wire signed [`CalcTempBus]          temp_b4_12_26_r;
wire signed [`CalcTempBus]          temp_b4_12_26_i;
wire signed [`CalcTempBus]          temp_b4_12_27_r;
wire signed [`CalcTempBus]          temp_b4_12_27_i;
wire signed [`CalcTempBus]          temp_b4_12_28_r;
wire signed [`CalcTempBus]          temp_b4_12_28_i;
wire signed [`CalcTempBus]          temp_b4_12_29_r;
wire signed [`CalcTempBus]          temp_b4_12_29_i;
wire signed [`CalcTempBus]          temp_b4_12_30_r;
wire signed [`CalcTempBus]          temp_b4_12_30_i;
wire signed [`CalcTempBus]          temp_b4_12_31_r;
wire signed [`CalcTempBus]          temp_b4_12_31_i;
wire signed [`CalcTempBus]          temp_b4_12_32_r;
wire signed [`CalcTempBus]          temp_b4_12_32_i;
wire signed [`CalcTempBus]          temp_b4_13_1_r;
wire signed [`CalcTempBus]          temp_b4_13_1_i;
wire signed [`CalcTempBus]          temp_b4_13_2_r;
wire signed [`CalcTempBus]          temp_b4_13_2_i;
wire signed [`CalcTempBus]          temp_b4_13_3_r;
wire signed [`CalcTempBus]          temp_b4_13_3_i;
wire signed [`CalcTempBus]          temp_b4_13_4_r;
wire signed [`CalcTempBus]          temp_b4_13_4_i;
wire signed [`CalcTempBus]          temp_b4_13_5_r;
wire signed [`CalcTempBus]          temp_b4_13_5_i;
wire signed [`CalcTempBus]          temp_b4_13_6_r;
wire signed [`CalcTempBus]          temp_b4_13_6_i;
wire signed [`CalcTempBus]          temp_b4_13_7_r;
wire signed [`CalcTempBus]          temp_b4_13_7_i;
wire signed [`CalcTempBus]          temp_b4_13_8_r;
wire signed [`CalcTempBus]          temp_b4_13_8_i;
wire signed [`CalcTempBus]          temp_b4_13_9_r;
wire signed [`CalcTempBus]          temp_b4_13_9_i;
wire signed [`CalcTempBus]          temp_b4_13_10_r;
wire signed [`CalcTempBus]          temp_b4_13_10_i;
wire signed [`CalcTempBus]          temp_b4_13_11_r;
wire signed [`CalcTempBus]          temp_b4_13_11_i;
wire signed [`CalcTempBus]          temp_b4_13_12_r;
wire signed [`CalcTempBus]          temp_b4_13_12_i;
wire signed [`CalcTempBus]          temp_b4_13_13_r;
wire signed [`CalcTempBus]          temp_b4_13_13_i;
wire signed [`CalcTempBus]          temp_b4_13_14_r;
wire signed [`CalcTempBus]          temp_b4_13_14_i;
wire signed [`CalcTempBus]          temp_b4_13_15_r;
wire signed [`CalcTempBus]          temp_b4_13_15_i;
wire signed [`CalcTempBus]          temp_b4_13_16_r;
wire signed [`CalcTempBus]          temp_b4_13_16_i;
wire signed [`CalcTempBus]          temp_b4_13_17_r;
wire signed [`CalcTempBus]          temp_b4_13_17_i;
wire signed [`CalcTempBus]          temp_b4_13_18_r;
wire signed [`CalcTempBus]          temp_b4_13_18_i;
wire signed [`CalcTempBus]          temp_b4_13_19_r;
wire signed [`CalcTempBus]          temp_b4_13_19_i;
wire signed [`CalcTempBus]          temp_b4_13_20_r;
wire signed [`CalcTempBus]          temp_b4_13_20_i;
wire signed [`CalcTempBus]          temp_b4_13_21_r;
wire signed [`CalcTempBus]          temp_b4_13_21_i;
wire signed [`CalcTempBus]          temp_b4_13_22_r;
wire signed [`CalcTempBus]          temp_b4_13_22_i;
wire signed [`CalcTempBus]          temp_b4_13_23_r;
wire signed [`CalcTempBus]          temp_b4_13_23_i;
wire signed [`CalcTempBus]          temp_b4_13_24_r;
wire signed [`CalcTempBus]          temp_b4_13_24_i;
wire signed [`CalcTempBus]          temp_b4_13_25_r;
wire signed [`CalcTempBus]          temp_b4_13_25_i;
wire signed [`CalcTempBus]          temp_b4_13_26_r;
wire signed [`CalcTempBus]          temp_b4_13_26_i;
wire signed [`CalcTempBus]          temp_b4_13_27_r;
wire signed [`CalcTempBus]          temp_b4_13_27_i;
wire signed [`CalcTempBus]          temp_b4_13_28_r;
wire signed [`CalcTempBus]          temp_b4_13_28_i;
wire signed [`CalcTempBus]          temp_b4_13_29_r;
wire signed [`CalcTempBus]          temp_b4_13_29_i;
wire signed [`CalcTempBus]          temp_b4_13_30_r;
wire signed [`CalcTempBus]          temp_b4_13_30_i;
wire signed [`CalcTempBus]          temp_b4_13_31_r;
wire signed [`CalcTempBus]          temp_b4_13_31_i;
wire signed [`CalcTempBus]          temp_b4_13_32_r;
wire signed [`CalcTempBus]          temp_b4_13_32_i;
wire signed [`CalcTempBus]          temp_b4_14_1_r;
wire signed [`CalcTempBus]          temp_b4_14_1_i;
wire signed [`CalcTempBus]          temp_b4_14_2_r;
wire signed [`CalcTempBus]          temp_b4_14_2_i;
wire signed [`CalcTempBus]          temp_b4_14_3_r;
wire signed [`CalcTempBus]          temp_b4_14_3_i;
wire signed [`CalcTempBus]          temp_b4_14_4_r;
wire signed [`CalcTempBus]          temp_b4_14_4_i;
wire signed [`CalcTempBus]          temp_b4_14_5_r;
wire signed [`CalcTempBus]          temp_b4_14_5_i;
wire signed [`CalcTempBus]          temp_b4_14_6_r;
wire signed [`CalcTempBus]          temp_b4_14_6_i;
wire signed [`CalcTempBus]          temp_b4_14_7_r;
wire signed [`CalcTempBus]          temp_b4_14_7_i;
wire signed [`CalcTempBus]          temp_b4_14_8_r;
wire signed [`CalcTempBus]          temp_b4_14_8_i;
wire signed [`CalcTempBus]          temp_b4_14_9_r;
wire signed [`CalcTempBus]          temp_b4_14_9_i;
wire signed [`CalcTempBus]          temp_b4_14_10_r;
wire signed [`CalcTempBus]          temp_b4_14_10_i;
wire signed [`CalcTempBus]          temp_b4_14_11_r;
wire signed [`CalcTempBus]          temp_b4_14_11_i;
wire signed [`CalcTempBus]          temp_b4_14_12_r;
wire signed [`CalcTempBus]          temp_b4_14_12_i;
wire signed [`CalcTempBus]          temp_b4_14_13_r;
wire signed [`CalcTempBus]          temp_b4_14_13_i;
wire signed [`CalcTempBus]          temp_b4_14_14_r;
wire signed [`CalcTempBus]          temp_b4_14_14_i;
wire signed [`CalcTempBus]          temp_b4_14_15_r;
wire signed [`CalcTempBus]          temp_b4_14_15_i;
wire signed [`CalcTempBus]          temp_b4_14_16_r;
wire signed [`CalcTempBus]          temp_b4_14_16_i;
wire signed [`CalcTempBus]          temp_b4_14_17_r;
wire signed [`CalcTempBus]          temp_b4_14_17_i;
wire signed [`CalcTempBus]          temp_b4_14_18_r;
wire signed [`CalcTempBus]          temp_b4_14_18_i;
wire signed [`CalcTempBus]          temp_b4_14_19_r;
wire signed [`CalcTempBus]          temp_b4_14_19_i;
wire signed [`CalcTempBus]          temp_b4_14_20_r;
wire signed [`CalcTempBus]          temp_b4_14_20_i;
wire signed [`CalcTempBus]          temp_b4_14_21_r;
wire signed [`CalcTempBus]          temp_b4_14_21_i;
wire signed [`CalcTempBus]          temp_b4_14_22_r;
wire signed [`CalcTempBus]          temp_b4_14_22_i;
wire signed [`CalcTempBus]          temp_b4_14_23_r;
wire signed [`CalcTempBus]          temp_b4_14_23_i;
wire signed [`CalcTempBus]          temp_b4_14_24_r;
wire signed [`CalcTempBus]          temp_b4_14_24_i;
wire signed [`CalcTempBus]          temp_b4_14_25_r;
wire signed [`CalcTempBus]          temp_b4_14_25_i;
wire signed [`CalcTempBus]          temp_b4_14_26_r;
wire signed [`CalcTempBus]          temp_b4_14_26_i;
wire signed [`CalcTempBus]          temp_b4_14_27_r;
wire signed [`CalcTempBus]          temp_b4_14_27_i;
wire signed [`CalcTempBus]          temp_b4_14_28_r;
wire signed [`CalcTempBus]          temp_b4_14_28_i;
wire signed [`CalcTempBus]          temp_b4_14_29_r;
wire signed [`CalcTempBus]          temp_b4_14_29_i;
wire signed [`CalcTempBus]          temp_b4_14_30_r;
wire signed [`CalcTempBus]          temp_b4_14_30_i;
wire signed [`CalcTempBus]          temp_b4_14_31_r;
wire signed [`CalcTempBus]          temp_b4_14_31_i;
wire signed [`CalcTempBus]          temp_b4_14_32_r;
wire signed [`CalcTempBus]          temp_b4_14_32_i;
wire signed [`CalcTempBus]          temp_b4_15_1_r;
wire signed [`CalcTempBus]          temp_b4_15_1_i;
wire signed [`CalcTempBus]          temp_b4_15_2_r;
wire signed [`CalcTempBus]          temp_b4_15_2_i;
wire signed [`CalcTempBus]          temp_b4_15_3_r;
wire signed [`CalcTempBus]          temp_b4_15_3_i;
wire signed [`CalcTempBus]          temp_b4_15_4_r;
wire signed [`CalcTempBus]          temp_b4_15_4_i;
wire signed [`CalcTempBus]          temp_b4_15_5_r;
wire signed [`CalcTempBus]          temp_b4_15_5_i;
wire signed [`CalcTempBus]          temp_b4_15_6_r;
wire signed [`CalcTempBus]          temp_b4_15_6_i;
wire signed [`CalcTempBus]          temp_b4_15_7_r;
wire signed [`CalcTempBus]          temp_b4_15_7_i;
wire signed [`CalcTempBus]          temp_b4_15_8_r;
wire signed [`CalcTempBus]          temp_b4_15_8_i;
wire signed [`CalcTempBus]          temp_b4_15_9_r;
wire signed [`CalcTempBus]          temp_b4_15_9_i;
wire signed [`CalcTempBus]          temp_b4_15_10_r;
wire signed [`CalcTempBus]          temp_b4_15_10_i;
wire signed [`CalcTempBus]          temp_b4_15_11_r;
wire signed [`CalcTempBus]          temp_b4_15_11_i;
wire signed [`CalcTempBus]          temp_b4_15_12_r;
wire signed [`CalcTempBus]          temp_b4_15_12_i;
wire signed [`CalcTempBus]          temp_b4_15_13_r;
wire signed [`CalcTempBus]          temp_b4_15_13_i;
wire signed [`CalcTempBus]          temp_b4_15_14_r;
wire signed [`CalcTempBus]          temp_b4_15_14_i;
wire signed [`CalcTempBus]          temp_b4_15_15_r;
wire signed [`CalcTempBus]          temp_b4_15_15_i;
wire signed [`CalcTempBus]          temp_b4_15_16_r;
wire signed [`CalcTempBus]          temp_b4_15_16_i;
wire signed [`CalcTempBus]          temp_b4_15_17_r;
wire signed [`CalcTempBus]          temp_b4_15_17_i;
wire signed [`CalcTempBus]          temp_b4_15_18_r;
wire signed [`CalcTempBus]          temp_b4_15_18_i;
wire signed [`CalcTempBus]          temp_b4_15_19_r;
wire signed [`CalcTempBus]          temp_b4_15_19_i;
wire signed [`CalcTempBus]          temp_b4_15_20_r;
wire signed [`CalcTempBus]          temp_b4_15_20_i;
wire signed [`CalcTempBus]          temp_b4_15_21_r;
wire signed [`CalcTempBus]          temp_b4_15_21_i;
wire signed [`CalcTempBus]          temp_b4_15_22_r;
wire signed [`CalcTempBus]          temp_b4_15_22_i;
wire signed [`CalcTempBus]          temp_b4_15_23_r;
wire signed [`CalcTempBus]          temp_b4_15_23_i;
wire signed [`CalcTempBus]          temp_b4_15_24_r;
wire signed [`CalcTempBus]          temp_b4_15_24_i;
wire signed [`CalcTempBus]          temp_b4_15_25_r;
wire signed [`CalcTempBus]          temp_b4_15_25_i;
wire signed [`CalcTempBus]          temp_b4_15_26_r;
wire signed [`CalcTempBus]          temp_b4_15_26_i;
wire signed [`CalcTempBus]          temp_b4_15_27_r;
wire signed [`CalcTempBus]          temp_b4_15_27_i;
wire signed [`CalcTempBus]          temp_b4_15_28_r;
wire signed [`CalcTempBus]          temp_b4_15_28_i;
wire signed [`CalcTempBus]          temp_b4_15_29_r;
wire signed [`CalcTempBus]          temp_b4_15_29_i;
wire signed [`CalcTempBus]          temp_b4_15_30_r;
wire signed [`CalcTempBus]          temp_b4_15_30_i;
wire signed [`CalcTempBus]          temp_b4_15_31_r;
wire signed [`CalcTempBus]          temp_b4_15_31_i;
wire signed [`CalcTempBus]          temp_b4_15_32_r;
wire signed [`CalcTempBus]          temp_b4_15_32_i;
wire signed [`CalcTempBus]          temp_b4_16_1_r;
wire signed [`CalcTempBus]          temp_b4_16_1_i;
wire signed [`CalcTempBus]          temp_b4_16_2_r;
wire signed [`CalcTempBus]          temp_b4_16_2_i;
wire signed [`CalcTempBus]          temp_b4_16_3_r;
wire signed [`CalcTempBus]          temp_b4_16_3_i;
wire signed [`CalcTempBus]          temp_b4_16_4_r;
wire signed [`CalcTempBus]          temp_b4_16_4_i;
wire signed [`CalcTempBus]          temp_b4_16_5_r;
wire signed [`CalcTempBus]          temp_b4_16_5_i;
wire signed [`CalcTempBus]          temp_b4_16_6_r;
wire signed [`CalcTempBus]          temp_b4_16_6_i;
wire signed [`CalcTempBus]          temp_b4_16_7_r;
wire signed [`CalcTempBus]          temp_b4_16_7_i;
wire signed [`CalcTempBus]          temp_b4_16_8_r;
wire signed [`CalcTempBus]          temp_b4_16_8_i;
wire signed [`CalcTempBus]          temp_b4_16_9_r;
wire signed [`CalcTempBus]          temp_b4_16_9_i;
wire signed [`CalcTempBus]          temp_b4_16_10_r;
wire signed [`CalcTempBus]          temp_b4_16_10_i;
wire signed [`CalcTempBus]          temp_b4_16_11_r;
wire signed [`CalcTempBus]          temp_b4_16_11_i;
wire signed [`CalcTempBus]          temp_b4_16_12_r;
wire signed [`CalcTempBus]          temp_b4_16_12_i;
wire signed [`CalcTempBus]          temp_b4_16_13_r;
wire signed [`CalcTempBus]          temp_b4_16_13_i;
wire signed [`CalcTempBus]          temp_b4_16_14_r;
wire signed [`CalcTempBus]          temp_b4_16_14_i;
wire signed [`CalcTempBus]          temp_b4_16_15_r;
wire signed [`CalcTempBus]          temp_b4_16_15_i;
wire signed [`CalcTempBus]          temp_b4_16_16_r;
wire signed [`CalcTempBus]          temp_b4_16_16_i;
wire signed [`CalcTempBus]          temp_b4_16_17_r;
wire signed [`CalcTempBus]          temp_b4_16_17_i;
wire signed [`CalcTempBus]          temp_b4_16_18_r;
wire signed [`CalcTempBus]          temp_b4_16_18_i;
wire signed [`CalcTempBus]          temp_b4_16_19_r;
wire signed [`CalcTempBus]          temp_b4_16_19_i;
wire signed [`CalcTempBus]          temp_b4_16_20_r;
wire signed [`CalcTempBus]          temp_b4_16_20_i;
wire signed [`CalcTempBus]          temp_b4_16_21_r;
wire signed [`CalcTempBus]          temp_b4_16_21_i;
wire signed [`CalcTempBus]          temp_b4_16_22_r;
wire signed [`CalcTempBus]          temp_b4_16_22_i;
wire signed [`CalcTempBus]          temp_b4_16_23_r;
wire signed [`CalcTempBus]          temp_b4_16_23_i;
wire signed [`CalcTempBus]          temp_b4_16_24_r;
wire signed [`CalcTempBus]          temp_b4_16_24_i;
wire signed [`CalcTempBus]          temp_b4_16_25_r;
wire signed [`CalcTempBus]          temp_b4_16_25_i;
wire signed [`CalcTempBus]          temp_b4_16_26_r;
wire signed [`CalcTempBus]          temp_b4_16_26_i;
wire signed [`CalcTempBus]          temp_b4_16_27_r;
wire signed [`CalcTempBus]          temp_b4_16_27_i;
wire signed [`CalcTempBus]          temp_b4_16_28_r;
wire signed [`CalcTempBus]          temp_b4_16_28_i;
wire signed [`CalcTempBus]          temp_b4_16_29_r;
wire signed [`CalcTempBus]          temp_b4_16_29_i;
wire signed [`CalcTempBus]          temp_b4_16_30_r;
wire signed [`CalcTempBus]          temp_b4_16_30_i;
wire signed [`CalcTempBus]          temp_b4_16_31_r;
wire signed [`CalcTempBus]          temp_b4_16_31_i;
wire signed [`CalcTempBus]          temp_b4_16_32_r;
wire signed [`CalcTempBus]          temp_b4_16_32_i;
wire signed [`CalcTempBus]          temp_b4_17_1_r;
wire signed [`CalcTempBus]          temp_b4_17_1_i;
wire signed [`CalcTempBus]          temp_b4_17_2_r;
wire signed [`CalcTempBus]          temp_b4_17_2_i;
wire signed [`CalcTempBus]          temp_b4_17_3_r;
wire signed [`CalcTempBus]          temp_b4_17_3_i;
wire signed [`CalcTempBus]          temp_b4_17_4_r;
wire signed [`CalcTempBus]          temp_b4_17_4_i;
wire signed [`CalcTempBus]          temp_b4_17_5_r;
wire signed [`CalcTempBus]          temp_b4_17_5_i;
wire signed [`CalcTempBus]          temp_b4_17_6_r;
wire signed [`CalcTempBus]          temp_b4_17_6_i;
wire signed [`CalcTempBus]          temp_b4_17_7_r;
wire signed [`CalcTempBus]          temp_b4_17_7_i;
wire signed [`CalcTempBus]          temp_b4_17_8_r;
wire signed [`CalcTempBus]          temp_b4_17_8_i;
wire signed [`CalcTempBus]          temp_b4_17_9_r;
wire signed [`CalcTempBus]          temp_b4_17_9_i;
wire signed [`CalcTempBus]          temp_b4_17_10_r;
wire signed [`CalcTempBus]          temp_b4_17_10_i;
wire signed [`CalcTempBus]          temp_b4_17_11_r;
wire signed [`CalcTempBus]          temp_b4_17_11_i;
wire signed [`CalcTempBus]          temp_b4_17_12_r;
wire signed [`CalcTempBus]          temp_b4_17_12_i;
wire signed [`CalcTempBus]          temp_b4_17_13_r;
wire signed [`CalcTempBus]          temp_b4_17_13_i;
wire signed [`CalcTempBus]          temp_b4_17_14_r;
wire signed [`CalcTempBus]          temp_b4_17_14_i;
wire signed [`CalcTempBus]          temp_b4_17_15_r;
wire signed [`CalcTempBus]          temp_b4_17_15_i;
wire signed [`CalcTempBus]          temp_b4_17_16_r;
wire signed [`CalcTempBus]          temp_b4_17_16_i;
wire signed [`CalcTempBus]          temp_b4_17_17_r;
wire signed [`CalcTempBus]          temp_b4_17_17_i;
wire signed [`CalcTempBus]          temp_b4_17_18_r;
wire signed [`CalcTempBus]          temp_b4_17_18_i;
wire signed [`CalcTempBus]          temp_b4_17_19_r;
wire signed [`CalcTempBus]          temp_b4_17_19_i;
wire signed [`CalcTempBus]          temp_b4_17_20_r;
wire signed [`CalcTempBus]          temp_b4_17_20_i;
wire signed [`CalcTempBus]          temp_b4_17_21_r;
wire signed [`CalcTempBus]          temp_b4_17_21_i;
wire signed [`CalcTempBus]          temp_b4_17_22_r;
wire signed [`CalcTempBus]          temp_b4_17_22_i;
wire signed [`CalcTempBus]          temp_b4_17_23_r;
wire signed [`CalcTempBus]          temp_b4_17_23_i;
wire signed [`CalcTempBus]          temp_b4_17_24_r;
wire signed [`CalcTempBus]          temp_b4_17_24_i;
wire signed [`CalcTempBus]          temp_b4_17_25_r;
wire signed [`CalcTempBus]          temp_b4_17_25_i;
wire signed [`CalcTempBus]          temp_b4_17_26_r;
wire signed [`CalcTempBus]          temp_b4_17_26_i;
wire signed [`CalcTempBus]          temp_b4_17_27_r;
wire signed [`CalcTempBus]          temp_b4_17_27_i;
wire signed [`CalcTempBus]          temp_b4_17_28_r;
wire signed [`CalcTempBus]          temp_b4_17_28_i;
wire signed [`CalcTempBus]          temp_b4_17_29_r;
wire signed [`CalcTempBus]          temp_b4_17_29_i;
wire signed [`CalcTempBus]          temp_b4_17_30_r;
wire signed [`CalcTempBus]          temp_b4_17_30_i;
wire signed [`CalcTempBus]          temp_b4_17_31_r;
wire signed [`CalcTempBus]          temp_b4_17_31_i;
wire signed [`CalcTempBus]          temp_b4_17_32_r;
wire signed [`CalcTempBus]          temp_b4_17_32_i;
wire signed [`CalcTempBus]          temp_b4_18_1_r;
wire signed [`CalcTempBus]          temp_b4_18_1_i;
wire signed [`CalcTempBus]          temp_b4_18_2_r;
wire signed [`CalcTempBus]          temp_b4_18_2_i;
wire signed [`CalcTempBus]          temp_b4_18_3_r;
wire signed [`CalcTempBus]          temp_b4_18_3_i;
wire signed [`CalcTempBus]          temp_b4_18_4_r;
wire signed [`CalcTempBus]          temp_b4_18_4_i;
wire signed [`CalcTempBus]          temp_b4_18_5_r;
wire signed [`CalcTempBus]          temp_b4_18_5_i;
wire signed [`CalcTempBus]          temp_b4_18_6_r;
wire signed [`CalcTempBus]          temp_b4_18_6_i;
wire signed [`CalcTempBus]          temp_b4_18_7_r;
wire signed [`CalcTempBus]          temp_b4_18_7_i;
wire signed [`CalcTempBus]          temp_b4_18_8_r;
wire signed [`CalcTempBus]          temp_b4_18_8_i;
wire signed [`CalcTempBus]          temp_b4_18_9_r;
wire signed [`CalcTempBus]          temp_b4_18_9_i;
wire signed [`CalcTempBus]          temp_b4_18_10_r;
wire signed [`CalcTempBus]          temp_b4_18_10_i;
wire signed [`CalcTempBus]          temp_b4_18_11_r;
wire signed [`CalcTempBus]          temp_b4_18_11_i;
wire signed [`CalcTempBus]          temp_b4_18_12_r;
wire signed [`CalcTempBus]          temp_b4_18_12_i;
wire signed [`CalcTempBus]          temp_b4_18_13_r;
wire signed [`CalcTempBus]          temp_b4_18_13_i;
wire signed [`CalcTempBus]          temp_b4_18_14_r;
wire signed [`CalcTempBus]          temp_b4_18_14_i;
wire signed [`CalcTempBus]          temp_b4_18_15_r;
wire signed [`CalcTempBus]          temp_b4_18_15_i;
wire signed [`CalcTempBus]          temp_b4_18_16_r;
wire signed [`CalcTempBus]          temp_b4_18_16_i;
wire signed [`CalcTempBus]          temp_b4_18_17_r;
wire signed [`CalcTempBus]          temp_b4_18_17_i;
wire signed [`CalcTempBus]          temp_b4_18_18_r;
wire signed [`CalcTempBus]          temp_b4_18_18_i;
wire signed [`CalcTempBus]          temp_b4_18_19_r;
wire signed [`CalcTempBus]          temp_b4_18_19_i;
wire signed [`CalcTempBus]          temp_b4_18_20_r;
wire signed [`CalcTempBus]          temp_b4_18_20_i;
wire signed [`CalcTempBus]          temp_b4_18_21_r;
wire signed [`CalcTempBus]          temp_b4_18_21_i;
wire signed [`CalcTempBus]          temp_b4_18_22_r;
wire signed [`CalcTempBus]          temp_b4_18_22_i;
wire signed [`CalcTempBus]          temp_b4_18_23_r;
wire signed [`CalcTempBus]          temp_b4_18_23_i;
wire signed [`CalcTempBus]          temp_b4_18_24_r;
wire signed [`CalcTempBus]          temp_b4_18_24_i;
wire signed [`CalcTempBus]          temp_b4_18_25_r;
wire signed [`CalcTempBus]          temp_b4_18_25_i;
wire signed [`CalcTempBus]          temp_b4_18_26_r;
wire signed [`CalcTempBus]          temp_b4_18_26_i;
wire signed [`CalcTempBus]          temp_b4_18_27_r;
wire signed [`CalcTempBus]          temp_b4_18_27_i;
wire signed [`CalcTempBus]          temp_b4_18_28_r;
wire signed [`CalcTempBus]          temp_b4_18_28_i;
wire signed [`CalcTempBus]          temp_b4_18_29_r;
wire signed [`CalcTempBus]          temp_b4_18_29_i;
wire signed [`CalcTempBus]          temp_b4_18_30_r;
wire signed [`CalcTempBus]          temp_b4_18_30_i;
wire signed [`CalcTempBus]          temp_b4_18_31_r;
wire signed [`CalcTempBus]          temp_b4_18_31_i;
wire signed [`CalcTempBus]          temp_b4_18_32_r;
wire signed [`CalcTempBus]          temp_b4_18_32_i;
wire signed [`CalcTempBus]          temp_b4_19_1_r;
wire signed [`CalcTempBus]          temp_b4_19_1_i;
wire signed [`CalcTempBus]          temp_b4_19_2_r;
wire signed [`CalcTempBus]          temp_b4_19_2_i;
wire signed [`CalcTempBus]          temp_b4_19_3_r;
wire signed [`CalcTempBus]          temp_b4_19_3_i;
wire signed [`CalcTempBus]          temp_b4_19_4_r;
wire signed [`CalcTempBus]          temp_b4_19_4_i;
wire signed [`CalcTempBus]          temp_b4_19_5_r;
wire signed [`CalcTempBus]          temp_b4_19_5_i;
wire signed [`CalcTempBus]          temp_b4_19_6_r;
wire signed [`CalcTempBus]          temp_b4_19_6_i;
wire signed [`CalcTempBus]          temp_b4_19_7_r;
wire signed [`CalcTempBus]          temp_b4_19_7_i;
wire signed [`CalcTempBus]          temp_b4_19_8_r;
wire signed [`CalcTempBus]          temp_b4_19_8_i;
wire signed [`CalcTempBus]          temp_b4_19_9_r;
wire signed [`CalcTempBus]          temp_b4_19_9_i;
wire signed [`CalcTempBus]          temp_b4_19_10_r;
wire signed [`CalcTempBus]          temp_b4_19_10_i;
wire signed [`CalcTempBus]          temp_b4_19_11_r;
wire signed [`CalcTempBus]          temp_b4_19_11_i;
wire signed [`CalcTempBus]          temp_b4_19_12_r;
wire signed [`CalcTempBus]          temp_b4_19_12_i;
wire signed [`CalcTempBus]          temp_b4_19_13_r;
wire signed [`CalcTempBus]          temp_b4_19_13_i;
wire signed [`CalcTempBus]          temp_b4_19_14_r;
wire signed [`CalcTempBus]          temp_b4_19_14_i;
wire signed [`CalcTempBus]          temp_b4_19_15_r;
wire signed [`CalcTempBus]          temp_b4_19_15_i;
wire signed [`CalcTempBus]          temp_b4_19_16_r;
wire signed [`CalcTempBus]          temp_b4_19_16_i;
wire signed [`CalcTempBus]          temp_b4_19_17_r;
wire signed [`CalcTempBus]          temp_b4_19_17_i;
wire signed [`CalcTempBus]          temp_b4_19_18_r;
wire signed [`CalcTempBus]          temp_b4_19_18_i;
wire signed [`CalcTempBus]          temp_b4_19_19_r;
wire signed [`CalcTempBus]          temp_b4_19_19_i;
wire signed [`CalcTempBus]          temp_b4_19_20_r;
wire signed [`CalcTempBus]          temp_b4_19_20_i;
wire signed [`CalcTempBus]          temp_b4_19_21_r;
wire signed [`CalcTempBus]          temp_b4_19_21_i;
wire signed [`CalcTempBus]          temp_b4_19_22_r;
wire signed [`CalcTempBus]          temp_b4_19_22_i;
wire signed [`CalcTempBus]          temp_b4_19_23_r;
wire signed [`CalcTempBus]          temp_b4_19_23_i;
wire signed [`CalcTempBus]          temp_b4_19_24_r;
wire signed [`CalcTempBus]          temp_b4_19_24_i;
wire signed [`CalcTempBus]          temp_b4_19_25_r;
wire signed [`CalcTempBus]          temp_b4_19_25_i;
wire signed [`CalcTempBus]          temp_b4_19_26_r;
wire signed [`CalcTempBus]          temp_b4_19_26_i;
wire signed [`CalcTempBus]          temp_b4_19_27_r;
wire signed [`CalcTempBus]          temp_b4_19_27_i;
wire signed [`CalcTempBus]          temp_b4_19_28_r;
wire signed [`CalcTempBus]          temp_b4_19_28_i;
wire signed [`CalcTempBus]          temp_b4_19_29_r;
wire signed [`CalcTempBus]          temp_b4_19_29_i;
wire signed [`CalcTempBus]          temp_b4_19_30_r;
wire signed [`CalcTempBus]          temp_b4_19_30_i;
wire signed [`CalcTempBus]          temp_b4_19_31_r;
wire signed [`CalcTempBus]          temp_b4_19_31_i;
wire signed [`CalcTempBus]          temp_b4_19_32_r;
wire signed [`CalcTempBus]          temp_b4_19_32_i;
wire signed [`CalcTempBus]          temp_b4_20_1_r;
wire signed [`CalcTempBus]          temp_b4_20_1_i;
wire signed [`CalcTempBus]          temp_b4_20_2_r;
wire signed [`CalcTempBus]          temp_b4_20_2_i;
wire signed [`CalcTempBus]          temp_b4_20_3_r;
wire signed [`CalcTempBus]          temp_b4_20_3_i;
wire signed [`CalcTempBus]          temp_b4_20_4_r;
wire signed [`CalcTempBus]          temp_b4_20_4_i;
wire signed [`CalcTempBus]          temp_b4_20_5_r;
wire signed [`CalcTempBus]          temp_b4_20_5_i;
wire signed [`CalcTempBus]          temp_b4_20_6_r;
wire signed [`CalcTempBus]          temp_b4_20_6_i;
wire signed [`CalcTempBus]          temp_b4_20_7_r;
wire signed [`CalcTempBus]          temp_b4_20_7_i;
wire signed [`CalcTempBus]          temp_b4_20_8_r;
wire signed [`CalcTempBus]          temp_b4_20_8_i;
wire signed [`CalcTempBus]          temp_b4_20_9_r;
wire signed [`CalcTempBus]          temp_b4_20_9_i;
wire signed [`CalcTempBus]          temp_b4_20_10_r;
wire signed [`CalcTempBus]          temp_b4_20_10_i;
wire signed [`CalcTempBus]          temp_b4_20_11_r;
wire signed [`CalcTempBus]          temp_b4_20_11_i;
wire signed [`CalcTempBus]          temp_b4_20_12_r;
wire signed [`CalcTempBus]          temp_b4_20_12_i;
wire signed [`CalcTempBus]          temp_b4_20_13_r;
wire signed [`CalcTempBus]          temp_b4_20_13_i;
wire signed [`CalcTempBus]          temp_b4_20_14_r;
wire signed [`CalcTempBus]          temp_b4_20_14_i;
wire signed [`CalcTempBus]          temp_b4_20_15_r;
wire signed [`CalcTempBus]          temp_b4_20_15_i;
wire signed [`CalcTempBus]          temp_b4_20_16_r;
wire signed [`CalcTempBus]          temp_b4_20_16_i;
wire signed [`CalcTempBus]          temp_b4_20_17_r;
wire signed [`CalcTempBus]          temp_b4_20_17_i;
wire signed [`CalcTempBus]          temp_b4_20_18_r;
wire signed [`CalcTempBus]          temp_b4_20_18_i;
wire signed [`CalcTempBus]          temp_b4_20_19_r;
wire signed [`CalcTempBus]          temp_b4_20_19_i;
wire signed [`CalcTempBus]          temp_b4_20_20_r;
wire signed [`CalcTempBus]          temp_b4_20_20_i;
wire signed [`CalcTempBus]          temp_b4_20_21_r;
wire signed [`CalcTempBus]          temp_b4_20_21_i;
wire signed [`CalcTempBus]          temp_b4_20_22_r;
wire signed [`CalcTempBus]          temp_b4_20_22_i;
wire signed [`CalcTempBus]          temp_b4_20_23_r;
wire signed [`CalcTempBus]          temp_b4_20_23_i;
wire signed [`CalcTempBus]          temp_b4_20_24_r;
wire signed [`CalcTempBus]          temp_b4_20_24_i;
wire signed [`CalcTempBus]          temp_b4_20_25_r;
wire signed [`CalcTempBus]          temp_b4_20_25_i;
wire signed [`CalcTempBus]          temp_b4_20_26_r;
wire signed [`CalcTempBus]          temp_b4_20_26_i;
wire signed [`CalcTempBus]          temp_b4_20_27_r;
wire signed [`CalcTempBus]          temp_b4_20_27_i;
wire signed [`CalcTempBus]          temp_b4_20_28_r;
wire signed [`CalcTempBus]          temp_b4_20_28_i;
wire signed [`CalcTempBus]          temp_b4_20_29_r;
wire signed [`CalcTempBus]          temp_b4_20_29_i;
wire signed [`CalcTempBus]          temp_b4_20_30_r;
wire signed [`CalcTempBus]          temp_b4_20_30_i;
wire signed [`CalcTempBus]          temp_b4_20_31_r;
wire signed [`CalcTempBus]          temp_b4_20_31_i;
wire signed [`CalcTempBus]          temp_b4_20_32_r;
wire signed [`CalcTempBus]          temp_b4_20_32_i;
wire signed [`CalcTempBus]          temp_b4_21_1_r;
wire signed [`CalcTempBus]          temp_b4_21_1_i;
wire signed [`CalcTempBus]          temp_b4_21_2_r;
wire signed [`CalcTempBus]          temp_b4_21_2_i;
wire signed [`CalcTempBus]          temp_b4_21_3_r;
wire signed [`CalcTempBus]          temp_b4_21_3_i;
wire signed [`CalcTempBus]          temp_b4_21_4_r;
wire signed [`CalcTempBus]          temp_b4_21_4_i;
wire signed [`CalcTempBus]          temp_b4_21_5_r;
wire signed [`CalcTempBus]          temp_b4_21_5_i;
wire signed [`CalcTempBus]          temp_b4_21_6_r;
wire signed [`CalcTempBus]          temp_b4_21_6_i;
wire signed [`CalcTempBus]          temp_b4_21_7_r;
wire signed [`CalcTempBus]          temp_b4_21_7_i;
wire signed [`CalcTempBus]          temp_b4_21_8_r;
wire signed [`CalcTempBus]          temp_b4_21_8_i;
wire signed [`CalcTempBus]          temp_b4_21_9_r;
wire signed [`CalcTempBus]          temp_b4_21_9_i;
wire signed [`CalcTempBus]          temp_b4_21_10_r;
wire signed [`CalcTempBus]          temp_b4_21_10_i;
wire signed [`CalcTempBus]          temp_b4_21_11_r;
wire signed [`CalcTempBus]          temp_b4_21_11_i;
wire signed [`CalcTempBus]          temp_b4_21_12_r;
wire signed [`CalcTempBus]          temp_b4_21_12_i;
wire signed [`CalcTempBus]          temp_b4_21_13_r;
wire signed [`CalcTempBus]          temp_b4_21_13_i;
wire signed [`CalcTempBus]          temp_b4_21_14_r;
wire signed [`CalcTempBus]          temp_b4_21_14_i;
wire signed [`CalcTempBus]          temp_b4_21_15_r;
wire signed [`CalcTempBus]          temp_b4_21_15_i;
wire signed [`CalcTempBus]          temp_b4_21_16_r;
wire signed [`CalcTempBus]          temp_b4_21_16_i;
wire signed [`CalcTempBus]          temp_b4_21_17_r;
wire signed [`CalcTempBus]          temp_b4_21_17_i;
wire signed [`CalcTempBus]          temp_b4_21_18_r;
wire signed [`CalcTempBus]          temp_b4_21_18_i;
wire signed [`CalcTempBus]          temp_b4_21_19_r;
wire signed [`CalcTempBus]          temp_b4_21_19_i;
wire signed [`CalcTempBus]          temp_b4_21_20_r;
wire signed [`CalcTempBus]          temp_b4_21_20_i;
wire signed [`CalcTempBus]          temp_b4_21_21_r;
wire signed [`CalcTempBus]          temp_b4_21_21_i;
wire signed [`CalcTempBus]          temp_b4_21_22_r;
wire signed [`CalcTempBus]          temp_b4_21_22_i;
wire signed [`CalcTempBus]          temp_b4_21_23_r;
wire signed [`CalcTempBus]          temp_b4_21_23_i;
wire signed [`CalcTempBus]          temp_b4_21_24_r;
wire signed [`CalcTempBus]          temp_b4_21_24_i;
wire signed [`CalcTempBus]          temp_b4_21_25_r;
wire signed [`CalcTempBus]          temp_b4_21_25_i;
wire signed [`CalcTempBus]          temp_b4_21_26_r;
wire signed [`CalcTempBus]          temp_b4_21_26_i;
wire signed [`CalcTempBus]          temp_b4_21_27_r;
wire signed [`CalcTempBus]          temp_b4_21_27_i;
wire signed [`CalcTempBus]          temp_b4_21_28_r;
wire signed [`CalcTempBus]          temp_b4_21_28_i;
wire signed [`CalcTempBus]          temp_b4_21_29_r;
wire signed [`CalcTempBus]          temp_b4_21_29_i;
wire signed [`CalcTempBus]          temp_b4_21_30_r;
wire signed [`CalcTempBus]          temp_b4_21_30_i;
wire signed [`CalcTempBus]          temp_b4_21_31_r;
wire signed [`CalcTempBus]          temp_b4_21_31_i;
wire signed [`CalcTempBus]          temp_b4_21_32_r;
wire signed [`CalcTempBus]          temp_b4_21_32_i;
wire signed [`CalcTempBus]          temp_b4_22_1_r;
wire signed [`CalcTempBus]          temp_b4_22_1_i;
wire signed [`CalcTempBus]          temp_b4_22_2_r;
wire signed [`CalcTempBus]          temp_b4_22_2_i;
wire signed [`CalcTempBus]          temp_b4_22_3_r;
wire signed [`CalcTempBus]          temp_b4_22_3_i;
wire signed [`CalcTempBus]          temp_b4_22_4_r;
wire signed [`CalcTempBus]          temp_b4_22_4_i;
wire signed [`CalcTempBus]          temp_b4_22_5_r;
wire signed [`CalcTempBus]          temp_b4_22_5_i;
wire signed [`CalcTempBus]          temp_b4_22_6_r;
wire signed [`CalcTempBus]          temp_b4_22_6_i;
wire signed [`CalcTempBus]          temp_b4_22_7_r;
wire signed [`CalcTempBus]          temp_b4_22_7_i;
wire signed [`CalcTempBus]          temp_b4_22_8_r;
wire signed [`CalcTempBus]          temp_b4_22_8_i;
wire signed [`CalcTempBus]          temp_b4_22_9_r;
wire signed [`CalcTempBus]          temp_b4_22_9_i;
wire signed [`CalcTempBus]          temp_b4_22_10_r;
wire signed [`CalcTempBus]          temp_b4_22_10_i;
wire signed [`CalcTempBus]          temp_b4_22_11_r;
wire signed [`CalcTempBus]          temp_b4_22_11_i;
wire signed [`CalcTempBus]          temp_b4_22_12_r;
wire signed [`CalcTempBus]          temp_b4_22_12_i;
wire signed [`CalcTempBus]          temp_b4_22_13_r;
wire signed [`CalcTempBus]          temp_b4_22_13_i;
wire signed [`CalcTempBus]          temp_b4_22_14_r;
wire signed [`CalcTempBus]          temp_b4_22_14_i;
wire signed [`CalcTempBus]          temp_b4_22_15_r;
wire signed [`CalcTempBus]          temp_b4_22_15_i;
wire signed [`CalcTempBus]          temp_b4_22_16_r;
wire signed [`CalcTempBus]          temp_b4_22_16_i;
wire signed [`CalcTempBus]          temp_b4_22_17_r;
wire signed [`CalcTempBus]          temp_b4_22_17_i;
wire signed [`CalcTempBus]          temp_b4_22_18_r;
wire signed [`CalcTempBus]          temp_b4_22_18_i;
wire signed [`CalcTempBus]          temp_b4_22_19_r;
wire signed [`CalcTempBus]          temp_b4_22_19_i;
wire signed [`CalcTempBus]          temp_b4_22_20_r;
wire signed [`CalcTempBus]          temp_b4_22_20_i;
wire signed [`CalcTempBus]          temp_b4_22_21_r;
wire signed [`CalcTempBus]          temp_b4_22_21_i;
wire signed [`CalcTempBus]          temp_b4_22_22_r;
wire signed [`CalcTempBus]          temp_b4_22_22_i;
wire signed [`CalcTempBus]          temp_b4_22_23_r;
wire signed [`CalcTempBus]          temp_b4_22_23_i;
wire signed [`CalcTempBus]          temp_b4_22_24_r;
wire signed [`CalcTempBus]          temp_b4_22_24_i;
wire signed [`CalcTempBus]          temp_b4_22_25_r;
wire signed [`CalcTempBus]          temp_b4_22_25_i;
wire signed [`CalcTempBus]          temp_b4_22_26_r;
wire signed [`CalcTempBus]          temp_b4_22_26_i;
wire signed [`CalcTempBus]          temp_b4_22_27_r;
wire signed [`CalcTempBus]          temp_b4_22_27_i;
wire signed [`CalcTempBus]          temp_b4_22_28_r;
wire signed [`CalcTempBus]          temp_b4_22_28_i;
wire signed [`CalcTempBus]          temp_b4_22_29_r;
wire signed [`CalcTempBus]          temp_b4_22_29_i;
wire signed [`CalcTempBus]          temp_b4_22_30_r;
wire signed [`CalcTempBus]          temp_b4_22_30_i;
wire signed [`CalcTempBus]          temp_b4_22_31_r;
wire signed [`CalcTempBus]          temp_b4_22_31_i;
wire signed [`CalcTempBus]          temp_b4_22_32_r;
wire signed [`CalcTempBus]          temp_b4_22_32_i;
wire signed [`CalcTempBus]          temp_b4_23_1_r;
wire signed [`CalcTempBus]          temp_b4_23_1_i;
wire signed [`CalcTempBus]          temp_b4_23_2_r;
wire signed [`CalcTempBus]          temp_b4_23_2_i;
wire signed [`CalcTempBus]          temp_b4_23_3_r;
wire signed [`CalcTempBus]          temp_b4_23_3_i;
wire signed [`CalcTempBus]          temp_b4_23_4_r;
wire signed [`CalcTempBus]          temp_b4_23_4_i;
wire signed [`CalcTempBus]          temp_b4_23_5_r;
wire signed [`CalcTempBus]          temp_b4_23_5_i;
wire signed [`CalcTempBus]          temp_b4_23_6_r;
wire signed [`CalcTempBus]          temp_b4_23_6_i;
wire signed [`CalcTempBus]          temp_b4_23_7_r;
wire signed [`CalcTempBus]          temp_b4_23_7_i;
wire signed [`CalcTempBus]          temp_b4_23_8_r;
wire signed [`CalcTempBus]          temp_b4_23_8_i;
wire signed [`CalcTempBus]          temp_b4_23_9_r;
wire signed [`CalcTempBus]          temp_b4_23_9_i;
wire signed [`CalcTempBus]          temp_b4_23_10_r;
wire signed [`CalcTempBus]          temp_b4_23_10_i;
wire signed [`CalcTempBus]          temp_b4_23_11_r;
wire signed [`CalcTempBus]          temp_b4_23_11_i;
wire signed [`CalcTempBus]          temp_b4_23_12_r;
wire signed [`CalcTempBus]          temp_b4_23_12_i;
wire signed [`CalcTempBus]          temp_b4_23_13_r;
wire signed [`CalcTempBus]          temp_b4_23_13_i;
wire signed [`CalcTempBus]          temp_b4_23_14_r;
wire signed [`CalcTempBus]          temp_b4_23_14_i;
wire signed [`CalcTempBus]          temp_b4_23_15_r;
wire signed [`CalcTempBus]          temp_b4_23_15_i;
wire signed [`CalcTempBus]          temp_b4_23_16_r;
wire signed [`CalcTempBus]          temp_b4_23_16_i;
wire signed [`CalcTempBus]          temp_b4_23_17_r;
wire signed [`CalcTempBus]          temp_b4_23_17_i;
wire signed [`CalcTempBus]          temp_b4_23_18_r;
wire signed [`CalcTempBus]          temp_b4_23_18_i;
wire signed [`CalcTempBus]          temp_b4_23_19_r;
wire signed [`CalcTempBus]          temp_b4_23_19_i;
wire signed [`CalcTempBus]          temp_b4_23_20_r;
wire signed [`CalcTempBus]          temp_b4_23_20_i;
wire signed [`CalcTempBus]          temp_b4_23_21_r;
wire signed [`CalcTempBus]          temp_b4_23_21_i;
wire signed [`CalcTempBus]          temp_b4_23_22_r;
wire signed [`CalcTempBus]          temp_b4_23_22_i;
wire signed [`CalcTempBus]          temp_b4_23_23_r;
wire signed [`CalcTempBus]          temp_b4_23_23_i;
wire signed [`CalcTempBus]          temp_b4_23_24_r;
wire signed [`CalcTempBus]          temp_b4_23_24_i;
wire signed [`CalcTempBus]          temp_b4_23_25_r;
wire signed [`CalcTempBus]          temp_b4_23_25_i;
wire signed [`CalcTempBus]          temp_b4_23_26_r;
wire signed [`CalcTempBus]          temp_b4_23_26_i;
wire signed [`CalcTempBus]          temp_b4_23_27_r;
wire signed [`CalcTempBus]          temp_b4_23_27_i;
wire signed [`CalcTempBus]          temp_b4_23_28_r;
wire signed [`CalcTempBus]          temp_b4_23_28_i;
wire signed [`CalcTempBus]          temp_b4_23_29_r;
wire signed [`CalcTempBus]          temp_b4_23_29_i;
wire signed [`CalcTempBus]          temp_b4_23_30_r;
wire signed [`CalcTempBus]          temp_b4_23_30_i;
wire signed [`CalcTempBus]          temp_b4_23_31_r;
wire signed [`CalcTempBus]          temp_b4_23_31_i;
wire signed [`CalcTempBus]          temp_b4_23_32_r;
wire signed [`CalcTempBus]          temp_b4_23_32_i;
wire signed [`CalcTempBus]          temp_b4_24_1_r;
wire signed [`CalcTempBus]          temp_b4_24_1_i;
wire signed [`CalcTempBus]          temp_b4_24_2_r;
wire signed [`CalcTempBus]          temp_b4_24_2_i;
wire signed [`CalcTempBus]          temp_b4_24_3_r;
wire signed [`CalcTempBus]          temp_b4_24_3_i;
wire signed [`CalcTempBus]          temp_b4_24_4_r;
wire signed [`CalcTempBus]          temp_b4_24_4_i;
wire signed [`CalcTempBus]          temp_b4_24_5_r;
wire signed [`CalcTempBus]          temp_b4_24_5_i;
wire signed [`CalcTempBus]          temp_b4_24_6_r;
wire signed [`CalcTempBus]          temp_b4_24_6_i;
wire signed [`CalcTempBus]          temp_b4_24_7_r;
wire signed [`CalcTempBus]          temp_b4_24_7_i;
wire signed [`CalcTempBus]          temp_b4_24_8_r;
wire signed [`CalcTempBus]          temp_b4_24_8_i;
wire signed [`CalcTempBus]          temp_b4_24_9_r;
wire signed [`CalcTempBus]          temp_b4_24_9_i;
wire signed [`CalcTempBus]          temp_b4_24_10_r;
wire signed [`CalcTempBus]          temp_b4_24_10_i;
wire signed [`CalcTempBus]          temp_b4_24_11_r;
wire signed [`CalcTempBus]          temp_b4_24_11_i;
wire signed [`CalcTempBus]          temp_b4_24_12_r;
wire signed [`CalcTempBus]          temp_b4_24_12_i;
wire signed [`CalcTempBus]          temp_b4_24_13_r;
wire signed [`CalcTempBus]          temp_b4_24_13_i;
wire signed [`CalcTempBus]          temp_b4_24_14_r;
wire signed [`CalcTempBus]          temp_b4_24_14_i;
wire signed [`CalcTempBus]          temp_b4_24_15_r;
wire signed [`CalcTempBus]          temp_b4_24_15_i;
wire signed [`CalcTempBus]          temp_b4_24_16_r;
wire signed [`CalcTempBus]          temp_b4_24_16_i;
wire signed [`CalcTempBus]          temp_b4_24_17_r;
wire signed [`CalcTempBus]          temp_b4_24_17_i;
wire signed [`CalcTempBus]          temp_b4_24_18_r;
wire signed [`CalcTempBus]          temp_b4_24_18_i;
wire signed [`CalcTempBus]          temp_b4_24_19_r;
wire signed [`CalcTempBus]          temp_b4_24_19_i;
wire signed [`CalcTempBus]          temp_b4_24_20_r;
wire signed [`CalcTempBus]          temp_b4_24_20_i;
wire signed [`CalcTempBus]          temp_b4_24_21_r;
wire signed [`CalcTempBus]          temp_b4_24_21_i;
wire signed [`CalcTempBus]          temp_b4_24_22_r;
wire signed [`CalcTempBus]          temp_b4_24_22_i;
wire signed [`CalcTempBus]          temp_b4_24_23_r;
wire signed [`CalcTempBus]          temp_b4_24_23_i;
wire signed [`CalcTempBus]          temp_b4_24_24_r;
wire signed [`CalcTempBus]          temp_b4_24_24_i;
wire signed [`CalcTempBus]          temp_b4_24_25_r;
wire signed [`CalcTempBus]          temp_b4_24_25_i;
wire signed [`CalcTempBus]          temp_b4_24_26_r;
wire signed [`CalcTempBus]          temp_b4_24_26_i;
wire signed [`CalcTempBus]          temp_b4_24_27_r;
wire signed [`CalcTempBus]          temp_b4_24_27_i;
wire signed [`CalcTempBus]          temp_b4_24_28_r;
wire signed [`CalcTempBus]          temp_b4_24_28_i;
wire signed [`CalcTempBus]          temp_b4_24_29_r;
wire signed [`CalcTempBus]          temp_b4_24_29_i;
wire signed [`CalcTempBus]          temp_b4_24_30_r;
wire signed [`CalcTempBus]          temp_b4_24_30_i;
wire signed [`CalcTempBus]          temp_b4_24_31_r;
wire signed [`CalcTempBus]          temp_b4_24_31_i;
wire signed [`CalcTempBus]          temp_b4_24_32_r;
wire signed [`CalcTempBus]          temp_b4_24_32_i;
wire signed [`CalcTempBus]          temp_b4_25_1_r;
wire signed [`CalcTempBus]          temp_b4_25_1_i;
wire signed [`CalcTempBus]          temp_b4_25_2_r;
wire signed [`CalcTempBus]          temp_b4_25_2_i;
wire signed [`CalcTempBus]          temp_b4_25_3_r;
wire signed [`CalcTempBus]          temp_b4_25_3_i;
wire signed [`CalcTempBus]          temp_b4_25_4_r;
wire signed [`CalcTempBus]          temp_b4_25_4_i;
wire signed [`CalcTempBus]          temp_b4_25_5_r;
wire signed [`CalcTempBus]          temp_b4_25_5_i;
wire signed [`CalcTempBus]          temp_b4_25_6_r;
wire signed [`CalcTempBus]          temp_b4_25_6_i;
wire signed [`CalcTempBus]          temp_b4_25_7_r;
wire signed [`CalcTempBus]          temp_b4_25_7_i;
wire signed [`CalcTempBus]          temp_b4_25_8_r;
wire signed [`CalcTempBus]          temp_b4_25_8_i;
wire signed [`CalcTempBus]          temp_b4_25_9_r;
wire signed [`CalcTempBus]          temp_b4_25_9_i;
wire signed [`CalcTempBus]          temp_b4_25_10_r;
wire signed [`CalcTempBus]          temp_b4_25_10_i;
wire signed [`CalcTempBus]          temp_b4_25_11_r;
wire signed [`CalcTempBus]          temp_b4_25_11_i;
wire signed [`CalcTempBus]          temp_b4_25_12_r;
wire signed [`CalcTempBus]          temp_b4_25_12_i;
wire signed [`CalcTempBus]          temp_b4_25_13_r;
wire signed [`CalcTempBus]          temp_b4_25_13_i;
wire signed [`CalcTempBus]          temp_b4_25_14_r;
wire signed [`CalcTempBus]          temp_b4_25_14_i;
wire signed [`CalcTempBus]          temp_b4_25_15_r;
wire signed [`CalcTempBus]          temp_b4_25_15_i;
wire signed [`CalcTempBus]          temp_b4_25_16_r;
wire signed [`CalcTempBus]          temp_b4_25_16_i;
wire signed [`CalcTempBus]          temp_b4_25_17_r;
wire signed [`CalcTempBus]          temp_b4_25_17_i;
wire signed [`CalcTempBus]          temp_b4_25_18_r;
wire signed [`CalcTempBus]          temp_b4_25_18_i;
wire signed [`CalcTempBus]          temp_b4_25_19_r;
wire signed [`CalcTempBus]          temp_b4_25_19_i;
wire signed [`CalcTempBus]          temp_b4_25_20_r;
wire signed [`CalcTempBus]          temp_b4_25_20_i;
wire signed [`CalcTempBus]          temp_b4_25_21_r;
wire signed [`CalcTempBus]          temp_b4_25_21_i;
wire signed [`CalcTempBus]          temp_b4_25_22_r;
wire signed [`CalcTempBus]          temp_b4_25_22_i;
wire signed [`CalcTempBus]          temp_b4_25_23_r;
wire signed [`CalcTempBus]          temp_b4_25_23_i;
wire signed [`CalcTempBus]          temp_b4_25_24_r;
wire signed [`CalcTempBus]          temp_b4_25_24_i;
wire signed [`CalcTempBus]          temp_b4_25_25_r;
wire signed [`CalcTempBus]          temp_b4_25_25_i;
wire signed [`CalcTempBus]          temp_b4_25_26_r;
wire signed [`CalcTempBus]          temp_b4_25_26_i;
wire signed [`CalcTempBus]          temp_b4_25_27_r;
wire signed [`CalcTempBus]          temp_b4_25_27_i;
wire signed [`CalcTempBus]          temp_b4_25_28_r;
wire signed [`CalcTempBus]          temp_b4_25_28_i;
wire signed [`CalcTempBus]          temp_b4_25_29_r;
wire signed [`CalcTempBus]          temp_b4_25_29_i;
wire signed [`CalcTempBus]          temp_b4_25_30_r;
wire signed [`CalcTempBus]          temp_b4_25_30_i;
wire signed [`CalcTempBus]          temp_b4_25_31_r;
wire signed [`CalcTempBus]          temp_b4_25_31_i;
wire signed [`CalcTempBus]          temp_b4_25_32_r;
wire signed [`CalcTempBus]          temp_b4_25_32_i;
wire signed [`CalcTempBus]          temp_b4_26_1_r;
wire signed [`CalcTempBus]          temp_b4_26_1_i;
wire signed [`CalcTempBus]          temp_b4_26_2_r;
wire signed [`CalcTempBus]          temp_b4_26_2_i;
wire signed [`CalcTempBus]          temp_b4_26_3_r;
wire signed [`CalcTempBus]          temp_b4_26_3_i;
wire signed [`CalcTempBus]          temp_b4_26_4_r;
wire signed [`CalcTempBus]          temp_b4_26_4_i;
wire signed [`CalcTempBus]          temp_b4_26_5_r;
wire signed [`CalcTempBus]          temp_b4_26_5_i;
wire signed [`CalcTempBus]          temp_b4_26_6_r;
wire signed [`CalcTempBus]          temp_b4_26_6_i;
wire signed [`CalcTempBus]          temp_b4_26_7_r;
wire signed [`CalcTempBus]          temp_b4_26_7_i;
wire signed [`CalcTempBus]          temp_b4_26_8_r;
wire signed [`CalcTempBus]          temp_b4_26_8_i;
wire signed [`CalcTempBus]          temp_b4_26_9_r;
wire signed [`CalcTempBus]          temp_b4_26_9_i;
wire signed [`CalcTempBus]          temp_b4_26_10_r;
wire signed [`CalcTempBus]          temp_b4_26_10_i;
wire signed [`CalcTempBus]          temp_b4_26_11_r;
wire signed [`CalcTempBus]          temp_b4_26_11_i;
wire signed [`CalcTempBus]          temp_b4_26_12_r;
wire signed [`CalcTempBus]          temp_b4_26_12_i;
wire signed [`CalcTempBus]          temp_b4_26_13_r;
wire signed [`CalcTempBus]          temp_b4_26_13_i;
wire signed [`CalcTempBus]          temp_b4_26_14_r;
wire signed [`CalcTempBus]          temp_b4_26_14_i;
wire signed [`CalcTempBus]          temp_b4_26_15_r;
wire signed [`CalcTempBus]          temp_b4_26_15_i;
wire signed [`CalcTempBus]          temp_b4_26_16_r;
wire signed [`CalcTempBus]          temp_b4_26_16_i;
wire signed [`CalcTempBus]          temp_b4_26_17_r;
wire signed [`CalcTempBus]          temp_b4_26_17_i;
wire signed [`CalcTempBus]          temp_b4_26_18_r;
wire signed [`CalcTempBus]          temp_b4_26_18_i;
wire signed [`CalcTempBus]          temp_b4_26_19_r;
wire signed [`CalcTempBus]          temp_b4_26_19_i;
wire signed [`CalcTempBus]          temp_b4_26_20_r;
wire signed [`CalcTempBus]          temp_b4_26_20_i;
wire signed [`CalcTempBus]          temp_b4_26_21_r;
wire signed [`CalcTempBus]          temp_b4_26_21_i;
wire signed [`CalcTempBus]          temp_b4_26_22_r;
wire signed [`CalcTempBus]          temp_b4_26_22_i;
wire signed [`CalcTempBus]          temp_b4_26_23_r;
wire signed [`CalcTempBus]          temp_b4_26_23_i;
wire signed [`CalcTempBus]          temp_b4_26_24_r;
wire signed [`CalcTempBus]          temp_b4_26_24_i;
wire signed [`CalcTempBus]          temp_b4_26_25_r;
wire signed [`CalcTempBus]          temp_b4_26_25_i;
wire signed [`CalcTempBus]          temp_b4_26_26_r;
wire signed [`CalcTempBus]          temp_b4_26_26_i;
wire signed [`CalcTempBus]          temp_b4_26_27_r;
wire signed [`CalcTempBus]          temp_b4_26_27_i;
wire signed [`CalcTempBus]          temp_b4_26_28_r;
wire signed [`CalcTempBus]          temp_b4_26_28_i;
wire signed [`CalcTempBus]          temp_b4_26_29_r;
wire signed [`CalcTempBus]          temp_b4_26_29_i;
wire signed [`CalcTempBus]          temp_b4_26_30_r;
wire signed [`CalcTempBus]          temp_b4_26_30_i;
wire signed [`CalcTempBus]          temp_b4_26_31_r;
wire signed [`CalcTempBus]          temp_b4_26_31_i;
wire signed [`CalcTempBus]          temp_b4_26_32_r;
wire signed [`CalcTempBus]          temp_b4_26_32_i;
wire signed [`CalcTempBus]          temp_b4_27_1_r;
wire signed [`CalcTempBus]          temp_b4_27_1_i;
wire signed [`CalcTempBus]          temp_b4_27_2_r;
wire signed [`CalcTempBus]          temp_b4_27_2_i;
wire signed [`CalcTempBus]          temp_b4_27_3_r;
wire signed [`CalcTempBus]          temp_b4_27_3_i;
wire signed [`CalcTempBus]          temp_b4_27_4_r;
wire signed [`CalcTempBus]          temp_b4_27_4_i;
wire signed [`CalcTempBus]          temp_b4_27_5_r;
wire signed [`CalcTempBus]          temp_b4_27_5_i;
wire signed [`CalcTempBus]          temp_b4_27_6_r;
wire signed [`CalcTempBus]          temp_b4_27_6_i;
wire signed [`CalcTempBus]          temp_b4_27_7_r;
wire signed [`CalcTempBus]          temp_b4_27_7_i;
wire signed [`CalcTempBus]          temp_b4_27_8_r;
wire signed [`CalcTempBus]          temp_b4_27_8_i;
wire signed [`CalcTempBus]          temp_b4_27_9_r;
wire signed [`CalcTempBus]          temp_b4_27_9_i;
wire signed [`CalcTempBus]          temp_b4_27_10_r;
wire signed [`CalcTempBus]          temp_b4_27_10_i;
wire signed [`CalcTempBus]          temp_b4_27_11_r;
wire signed [`CalcTempBus]          temp_b4_27_11_i;
wire signed [`CalcTempBus]          temp_b4_27_12_r;
wire signed [`CalcTempBus]          temp_b4_27_12_i;
wire signed [`CalcTempBus]          temp_b4_27_13_r;
wire signed [`CalcTempBus]          temp_b4_27_13_i;
wire signed [`CalcTempBus]          temp_b4_27_14_r;
wire signed [`CalcTempBus]          temp_b4_27_14_i;
wire signed [`CalcTempBus]          temp_b4_27_15_r;
wire signed [`CalcTempBus]          temp_b4_27_15_i;
wire signed [`CalcTempBus]          temp_b4_27_16_r;
wire signed [`CalcTempBus]          temp_b4_27_16_i;
wire signed [`CalcTempBus]          temp_b4_27_17_r;
wire signed [`CalcTempBus]          temp_b4_27_17_i;
wire signed [`CalcTempBus]          temp_b4_27_18_r;
wire signed [`CalcTempBus]          temp_b4_27_18_i;
wire signed [`CalcTempBus]          temp_b4_27_19_r;
wire signed [`CalcTempBus]          temp_b4_27_19_i;
wire signed [`CalcTempBus]          temp_b4_27_20_r;
wire signed [`CalcTempBus]          temp_b4_27_20_i;
wire signed [`CalcTempBus]          temp_b4_27_21_r;
wire signed [`CalcTempBus]          temp_b4_27_21_i;
wire signed [`CalcTempBus]          temp_b4_27_22_r;
wire signed [`CalcTempBus]          temp_b4_27_22_i;
wire signed [`CalcTempBus]          temp_b4_27_23_r;
wire signed [`CalcTempBus]          temp_b4_27_23_i;
wire signed [`CalcTempBus]          temp_b4_27_24_r;
wire signed [`CalcTempBus]          temp_b4_27_24_i;
wire signed [`CalcTempBus]          temp_b4_27_25_r;
wire signed [`CalcTempBus]          temp_b4_27_25_i;
wire signed [`CalcTempBus]          temp_b4_27_26_r;
wire signed [`CalcTempBus]          temp_b4_27_26_i;
wire signed [`CalcTempBus]          temp_b4_27_27_r;
wire signed [`CalcTempBus]          temp_b4_27_27_i;
wire signed [`CalcTempBus]          temp_b4_27_28_r;
wire signed [`CalcTempBus]          temp_b4_27_28_i;
wire signed [`CalcTempBus]          temp_b4_27_29_r;
wire signed [`CalcTempBus]          temp_b4_27_29_i;
wire signed [`CalcTempBus]          temp_b4_27_30_r;
wire signed [`CalcTempBus]          temp_b4_27_30_i;
wire signed [`CalcTempBus]          temp_b4_27_31_r;
wire signed [`CalcTempBus]          temp_b4_27_31_i;
wire signed [`CalcTempBus]          temp_b4_27_32_r;
wire signed [`CalcTempBus]          temp_b4_27_32_i;
wire signed [`CalcTempBus]          temp_b4_28_1_r;
wire signed [`CalcTempBus]          temp_b4_28_1_i;
wire signed [`CalcTempBus]          temp_b4_28_2_r;
wire signed [`CalcTempBus]          temp_b4_28_2_i;
wire signed [`CalcTempBus]          temp_b4_28_3_r;
wire signed [`CalcTempBus]          temp_b4_28_3_i;
wire signed [`CalcTempBus]          temp_b4_28_4_r;
wire signed [`CalcTempBus]          temp_b4_28_4_i;
wire signed [`CalcTempBus]          temp_b4_28_5_r;
wire signed [`CalcTempBus]          temp_b4_28_5_i;
wire signed [`CalcTempBus]          temp_b4_28_6_r;
wire signed [`CalcTempBus]          temp_b4_28_6_i;
wire signed [`CalcTempBus]          temp_b4_28_7_r;
wire signed [`CalcTempBus]          temp_b4_28_7_i;
wire signed [`CalcTempBus]          temp_b4_28_8_r;
wire signed [`CalcTempBus]          temp_b4_28_8_i;
wire signed [`CalcTempBus]          temp_b4_28_9_r;
wire signed [`CalcTempBus]          temp_b4_28_9_i;
wire signed [`CalcTempBus]          temp_b4_28_10_r;
wire signed [`CalcTempBus]          temp_b4_28_10_i;
wire signed [`CalcTempBus]          temp_b4_28_11_r;
wire signed [`CalcTempBus]          temp_b4_28_11_i;
wire signed [`CalcTempBus]          temp_b4_28_12_r;
wire signed [`CalcTempBus]          temp_b4_28_12_i;
wire signed [`CalcTempBus]          temp_b4_28_13_r;
wire signed [`CalcTempBus]          temp_b4_28_13_i;
wire signed [`CalcTempBus]          temp_b4_28_14_r;
wire signed [`CalcTempBus]          temp_b4_28_14_i;
wire signed [`CalcTempBus]          temp_b4_28_15_r;
wire signed [`CalcTempBus]          temp_b4_28_15_i;
wire signed [`CalcTempBus]          temp_b4_28_16_r;
wire signed [`CalcTempBus]          temp_b4_28_16_i;
wire signed [`CalcTempBus]          temp_b4_28_17_r;
wire signed [`CalcTempBus]          temp_b4_28_17_i;
wire signed [`CalcTempBus]          temp_b4_28_18_r;
wire signed [`CalcTempBus]          temp_b4_28_18_i;
wire signed [`CalcTempBus]          temp_b4_28_19_r;
wire signed [`CalcTempBus]          temp_b4_28_19_i;
wire signed [`CalcTempBus]          temp_b4_28_20_r;
wire signed [`CalcTempBus]          temp_b4_28_20_i;
wire signed [`CalcTempBus]          temp_b4_28_21_r;
wire signed [`CalcTempBus]          temp_b4_28_21_i;
wire signed [`CalcTempBus]          temp_b4_28_22_r;
wire signed [`CalcTempBus]          temp_b4_28_22_i;
wire signed [`CalcTempBus]          temp_b4_28_23_r;
wire signed [`CalcTempBus]          temp_b4_28_23_i;
wire signed [`CalcTempBus]          temp_b4_28_24_r;
wire signed [`CalcTempBus]          temp_b4_28_24_i;
wire signed [`CalcTempBus]          temp_b4_28_25_r;
wire signed [`CalcTempBus]          temp_b4_28_25_i;
wire signed [`CalcTempBus]          temp_b4_28_26_r;
wire signed [`CalcTempBus]          temp_b4_28_26_i;
wire signed [`CalcTempBus]          temp_b4_28_27_r;
wire signed [`CalcTempBus]          temp_b4_28_27_i;
wire signed [`CalcTempBus]          temp_b4_28_28_r;
wire signed [`CalcTempBus]          temp_b4_28_28_i;
wire signed [`CalcTempBus]          temp_b4_28_29_r;
wire signed [`CalcTempBus]          temp_b4_28_29_i;
wire signed [`CalcTempBus]          temp_b4_28_30_r;
wire signed [`CalcTempBus]          temp_b4_28_30_i;
wire signed [`CalcTempBus]          temp_b4_28_31_r;
wire signed [`CalcTempBus]          temp_b4_28_31_i;
wire signed [`CalcTempBus]          temp_b4_28_32_r;
wire signed [`CalcTempBus]          temp_b4_28_32_i;
wire signed [`CalcTempBus]          temp_b4_29_1_r;
wire signed [`CalcTempBus]          temp_b4_29_1_i;
wire signed [`CalcTempBus]          temp_b4_29_2_r;
wire signed [`CalcTempBus]          temp_b4_29_2_i;
wire signed [`CalcTempBus]          temp_b4_29_3_r;
wire signed [`CalcTempBus]          temp_b4_29_3_i;
wire signed [`CalcTempBus]          temp_b4_29_4_r;
wire signed [`CalcTempBus]          temp_b4_29_4_i;
wire signed [`CalcTempBus]          temp_b4_29_5_r;
wire signed [`CalcTempBus]          temp_b4_29_5_i;
wire signed [`CalcTempBus]          temp_b4_29_6_r;
wire signed [`CalcTempBus]          temp_b4_29_6_i;
wire signed [`CalcTempBus]          temp_b4_29_7_r;
wire signed [`CalcTempBus]          temp_b4_29_7_i;
wire signed [`CalcTempBus]          temp_b4_29_8_r;
wire signed [`CalcTempBus]          temp_b4_29_8_i;
wire signed [`CalcTempBus]          temp_b4_29_9_r;
wire signed [`CalcTempBus]          temp_b4_29_9_i;
wire signed [`CalcTempBus]          temp_b4_29_10_r;
wire signed [`CalcTempBus]          temp_b4_29_10_i;
wire signed [`CalcTempBus]          temp_b4_29_11_r;
wire signed [`CalcTempBus]          temp_b4_29_11_i;
wire signed [`CalcTempBus]          temp_b4_29_12_r;
wire signed [`CalcTempBus]          temp_b4_29_12_i;
wire signed [`CalcTempBus]          temp_b4_29_13_r;
wire signed [`CalcTempBus]          temp_b4_29_13_i;
wire signed [`CalcTempBus]          temp_b4_29_14_r;
wire signed [`CalcTempBus]          temp_b4_29_14_i;
wire signed [`CalcTempBus]          temp_b4_29_15_r;
wire signed [`CalcTempBus]          temp_b4_29_15_i;
wire signed [`CalcTempBus]          temp_b4_29_16_r;
wire signed [`CalcTempBus]          temp_b4_29_16_i;
wire signed [`CalcTempBus]          temp_b4_29_17_r;
wire signed [`CalcTempBus]          temp_b4_29_17_i;
wire signed [`CalcTempBus]          temp_b4_29_18_r;
wire signed [`CalcTempBus]          temp_b4_29_18_i;
wire signed [`CalcTempBus]          temp_b4_29_19_r;
wire signed [`CalcTempBus]          temp_b4_29_19_i;
wire signed [`CalcTempBus]          temp_b4_29_20_r;
wire signed [`CalcTempBus]          temp_b4_29_20_i;
wire signed [`CalcTempBus]          temp_b4_29_21_r;
wire signed [`CalcTempBus]          temp_b4_29_21_i;
wire signed [`CalcTempBus]          temp_b4_29_22_r;
wire signed [`CalcTempBus]          temp_b4_29_22_i;
wire signed [`CalcTempBus]          temp_b4_29_23_r;
wire signed [`CalcTempBus]          temp_b4_29_23_i;
wire signed [`CalcTempBus]          temp_b4_29_24_r;
wire signed [`CalcTempBus]          temp_b4_29_24_i;
wire signed [`CalcTempBus]          temp_b4_29_25_r;
wire signed [`CalcTempBus]          temp_b4_29_25_i;
wire signed [`CalcTempBus]          temp_b4_29_26_r;
wire signed [`CalcTempBus]          temp_b4_29_26_i;
wire signed [`CalcTempBus]          temp_b4_29_27_r;
wire signed [`CalcTempBus]          temp_b4_29_27_i;
wire signed [`CalcTempBus]          temp_b4_29_28_r;
wire signed [`CalcTempBus]          temp_b4_29_28_i;
wire signed [`CalcTempBus]          temp_b4_29_29_r;
wire signed [`CalcTempBus]          temp_b4_29_29_i;
wire signed [`CalcTempBus]          temp_b4_29_30_r;
wire signed [`CalcTempBus]          temp_b4_29_30_i;
wire signed [`CalcTempBus]          temp_b4_29_31_r;
wire signed [`CalcTempBus]          temp_b4_29_31_i;
wire signed [`CalcTempBus]          temp_b4_29_32_r;
wire signed [`CalcTempBus]          temp_b4_29_32_i;
wire signed [`CalcTempBus]          temp_b4_30_1_r;
wire signed [`CalcTempBus]          temp_b4_30_1_i;
wire signed [`CalcTempBus]          temp_b4_30_2_r;
wire signed [`CalcTempBus]          temp_b4_30_2_i;
wire signed [`CalcTempBus]          temp_b4_30_3_r;
wire signed [`CalcTempBus]          temp_b4_30_3_i;
wire signed [`CalcTempBus]          temp_b4_30_4_r;
wire signed [`CalcTempBus]          temp_b4_30_4_i;
wire signed [`CalcTempBus]          temp_b4_30_5_r;
wire signed [`CalcTempBus]          temp_b4_30_5_i;
wire signed [`CalcTempBus]          temp_b4_30_6_r;
wire signed [`CalcTempBus]          temp_b4_30_6_i;
wire signed [`CalcTempBus]          temp_b4_30_7_r;
wire signed [`CalcTempBus]          temp_b4_30_7_i;
wire signed [`CalcTempBus]          temp_b4_30_8_r;
wire signed [`CalcTempBus]          temp_b4_30_8_i;
wire signed [`CalcTempBus]          temp_b4_30_9_r;
wire signed [`CalcTempBus]          temp_b4_30_9_i;
wire signed [`CalcTempBus]          temp_b4_30_10_r;
wire signed [`CalcTempBus]          temp_b4_30_10_i;
wire signed [`CalcTempBus]          temp_b4_30_11_r;
wire signed [`CalcTempBus]          temp_b4_30_11_i;
wire signed [`CalcTempBus]          temp_b4_30_12_r;
wire signed [`CalcTempBus]          temp_b4_30_12_i;
wire signed [`CalcTempBus]          temp_b4_30_13_r;
wire signed [`CalcTempBus]          temp_b4_30_13_i;
wire signed [`CalcTempBus]          temp_b4_30_14_r;
wire signed [`CalcTempBus]          temp_b4_30_14_i;
wire signed [`CalcTempBus]          temp_b4_30_15_r;
wire signed [`CalcTempBus]          temp_b4_30_15_i;
wire signed [`CalcTempBus]          temp_b4_30_16_r;
wire signed [`CalcTempBus]          temp_b4_30_16_i;
wire signed [`CalcTempBus]          temp_b4_30_17_r;
wire signed [`CalcTempBus]          temp_b4_30_17_i;
wire signed [`CalcTempBus]          temp_b4_30_18_r;
wire signed [`CalcTempBus]          temp_b4_30_18_i;
wire signed [`CalcTempBus]          temp_b4_30_19_r;
wire signed [`CalcTempBus]          temp_b4_30_19_i;
wire signed [`CalcTempBus]          temp_b4_30_20_r;
wire signed [`CalcTempBus]          temp_b4_30_20_i;
wire signed [`CalcTempBus]          temp_b4_30_21_r;
wire signed [`CalcTempBus]          temp_b4_30_21_i;
wire signed [`CalcTempBus]          temp_b4_30_22_r;
wire signed [`CalcTempBus]          temp_b4_30_22_i;
wire signed [`CalcTempBus]          temp_b4_30_23_r;
wire signed [`CalcTempBus]          temp_b4_30_23_i;
wire signed [`CalcTempBus]          temp_b4_30_24_r;
wire signed [`CalcTempBus]          temp_b4_30_24_i;
wire signed [`CalcTempBus]          temp_b4_30_25_r;
wire signed [`CalcTempBus]          temp_b4_30_25_i;
wire signed [`CalcTempBus]          temp_b4_30_26_r;
wire signed [`CalcTempBus]          temp_b4_30_26_i;
wire signed [`CalcTempBus]          temp_b4_30_27_r;
wire signed [`CalcTempBus]          temp_b4_30_27_i;
wire signed [`CalcTempBus]          temp_b4_30_28_r;
wire signed [`CalcTempBus]          temp_b4_30_28_i;
wire signed [`CalcTempBus]          temp_b4_30_29_r;
wire signed [`CalcTempBus]          temp_b4_30_29_i;
wire signed [`CalcTempBus]          temp_b4_30_30_r;
wire signed [`CalcTempBus]          temp_b4_30_30_i;
wire signed [`CalcTempBus]          temp_b4_30_31_r;
wire signed [`CalcTempBus]          temp_b4_30_31_i;
wire signed [`CalcTempBus]          temp_b4_30_32_r;
wire signed [`CalcTempBus]          temp_b4_30_32_i;
wire signed [`CalcTempBus]          temp_b4_31_1_r;
wire signed [`CalcTempBus]          temp_b4_31_1_i;
wire signed [`CalcTempBus]          temp_b4_31_2_r;
wire signed [`CalcTempBus]          temp_b4_31_2_i;
wire signed [`CalcTempBus]          temp_b4_31_3_r;
wire signed [`CalcTempBus]          temp_b4_31_3_i;
wire signed [`CalcTempBus]          temp_b4_31_4_r;
wire signed [`CalcTempBus]          temp_b4_31_4_i;
wire signed [`CalcTempBus]          temp_b4_31_5_r;
wire signed [`CalcTempBus]          temp_b4_31_5_i;
wire signed [`CalcTempBus]          temp_b4_31_6_r;
wire signed [`CalcTempBus]          temp_b4_31_6_i;
wire signed [`CalcTempBus]          temp_b4_31_7_r;
wire signed [`CalcTempBus]          temp_b4_31_7_i;
wire signed [`CalcTempBus]          temp_b4_31_8_r;
wire signed [`CalcTempBus]          temp_b4_31_8_i;
wire signed [`CalcTempBus]          temp_b4_31_9_r;
wire signed [`CalcTempBus]          temp_b4_31_9_i;
wire signed [`CalcTempBus]          temp_b4_31_10_r;
wire signed [`CalcTempBus]          temp_b4_31_10_i;
wire signed [`CalcTempBus]          temp_b4_31_11_r;
wire signed [`CalcTempBus]          temp_b4_31_11_i;
wire signed [`CalcTempBus]          temp_b4_31_12_r;
wire signed [`CalcTempBus]          temp_b4_31_12_i;
wire signed [`CalcTempBus]          temp_b4_31_13_r;
wire signed [`CalcTempBus]          temp_b4_31_13_i;
wire signed [`CalcTempBus]          temp_b4_31_14_r;
wire signed [`CalcTempBus]          temp_b4_31_14_i;
wire signed [`CalcTempBus]          temp_b4_31_15_r;
wire signed [`CalcTempBus]          temp_b4_31_15_i;
wire signed [`CalcTempBus]          temp_b4_31_16_r;
wire signed [`CalcTempBus]          temp_b4_31_16_i;
wire signed [`CalcTempBus]          temp_b4_31_17_r;
wire signed [`CalcTempBus]          temp_b4_31_17_i;
wire signed [`CalcTempBus]          temp_b4_31_18_r;
wire signed [`CalcTempBus]          temp_b4_31_18_i;
wire signed [`CalcTempBus]          temp_b4_31_19_r;
wire signed [`CalcTempBus]          temp_b4_31_19_i;
wire signed [`CalcTempBus]          temp_b4_31_20_r;
wire signed [`CalcTempBus]          temp_b4_31_20_i;
wire signed [`CalcTempBus]          temp_b4_31_21_r;
wire signed [`CalcTempBus]          temp_b4_31_21_i;
wire signed [`CalcTempBus]          temp_b4_31_22_r;
wire signed [`CalcTempBus]          temp_b4_31_22_i;
wire signed [`CalcTempBus]          temp_b4_31_23_r;
wire signed [`CalcTempBus]          temp_b4_31_23_i;
wire signed [`CalcTempBus]          temp_b4_31_24_r;
wire signed [`CalcTempBus]          temp_b4_31_24_i;
wire signed [`CalcTempBus]          temp_b4_31_25_r;
wire signed [`CalcTempBus]          temp_b4_31_25_i;
wire signed [`CalcTempBus]          temp_b4_31_26_r;
wire signed [`CalcTempBus]          temp_b4_31_26_i;
wire signed [`CalcTempBus]          temp_b4_31_27_r;
wire signed [`CalcTempBus]          temp_b4_31_27_i;
wire signed [`CalcTempBus]          temp_b4_31_28_r;
wire signed [`CalcTempBus]          temp_b4_31_28_i;
wire signed [`CalcTempBus]          temp_b4_31_29_r;
wire signed [`CalcTempBus]          temp_b4_31_29_i;
wire signed [`CalcTempBus]          temp_b4_31_30_r;
wire signed [`CalcTempBus]          temp_b4_31_30_i;
wire signed [`CalcTempBus]          temp_b4_31_31_r;
wire signed [`CalcTempBus]          temp_b4_31_31_i;
wire signed [`CalcTempBus]          temp_b4_31_32_r;
wire signed [`CalcTempBus]          temp_b4_31_32_i;
wire signed [`CalcTempBus]          temp_b4_32_1_r;
wire signed [`CalcTempBus]          temp_b4_32_1_i;
wire signed [`CalcTempBus]          temp_b4_32_2_r;
wire signed [`CalcTempBus]          temp_b4_32_2_i;
wire signed [`CalcTempBus]          temp_b4_32_3_r;
wire signed [`CalcTempBus]          temp_b4_32_3_i;
wire signed [`CalcTempBus]          temp_b4_32_4_r;
wire signed [`CalcTempBus]          temp_b4_32_4_i;
wire signed [`CalcTempBus]          temp_b4_32_5_r;
wire signed [`CalcTempBus]          temp_b4_32_5_i;
wire signed [`CalcTempBus]          temp_b4_32_6_r;
wire signed [`CalcTempBus]          temp_b4_32_6_i;
wire signed [`CalcTempBus]          temp_b4_32_7_r;
wire signed [`CalcTempBus]          temp_b4_32_7_i;
wire signed [`CalcTempBus]          temp_b4_32_8_r;
wire signed [`CalcTempBus]          temp_b4_32_8_i;
wire signed [`CalcTempBus]          temp_b4_32_9_r;
wire signed [`CalcTempBus]          temp_b4_32_9_i;
wire signed [`CalcTempBus]          temp_b4_32_10_r;
wire signed [`CalcTempBus]          temp_b4_32_10_i;
wire signed [`CalcTempBus]          temp_b4_32_11_r;
wire signed [`CalcTempBus]          temp_b4_32_11_i;
wire signed [`CalcTempBus]          temp_b4_32_12_r;
wire signed [`CalcTempBus]          temp_b4_32_12_i;
wire signed [`CalcTempBus]          temp_b4_32_13_r;
wire signed [`CalcTempBus]          temp_b4_32_13_i;
wire signed [`CalcTempBus]          temp_b4_32_14_r;
wire signed [`CalcTempBus]          temp_b4_32_14_i;
wire signed [`CalcTempBus]          temp_b4_32_15_r;
wire signed [`CalcTempBus]          temp_b4_32_15_i;
wire signed [`CalcTempBus]          temp_b4_32_16_r;
wire signed [`CalcTempBus]          temp_b4_32_16_i;
wire signed [`CalcTempBus]          temp_b4_32_17_r;
wire signed [`CalcTempBus]          temp_b4_32_17_i;
wire signed [`CalcTempBus]          temp_b4_32_18_r;
wire signed [`CalcTempBus]          temp_b4_32_18_i;
wire signed [`CalcTempBus]          temp_b4_32_19_r;
wire signed [`CalcTempBus]          temp_b4_32_19_i;
wire signed [`CalcTempBus]          temp_b4_32_20_r;
wire signed [`CalcTempBus]          temp_b4_32_20_i;
wire signed [`CalcTempBus]          temp_b4_32_21_r;
wire signed [`CalcTempBus]          temp_b4_32_21_i;
wire signed [`CalcTempBus]          temp_b4_32_22_r;
wire signed [`CalcTempBus]          temp_b4_32_22_i;
wire signed [`CalcTempBus]          temp_b4_32_23_r;
wire signed [`CalcTempBus]          temp_b4_32_23_i;
wire signed [`CalcTempBus]          temp_b4_32_24_r;
wire signed [`CalcTempBus]          temp_b4_32_24_i;
wire signed [`CalcTempBus]          temp_b4_32_25_r;
wire signed [`CalcTempBus]          temp_b4_32_25_i;
wire signed [`CalcTempBus]          temp_b4_32_26_r;
wire signed [`CalcTempBus]          temp_b4_32_26_i;
wire signed [`CalcTempBus]          temp_b4_32_27_r;
wire signed [`CalcTempBus]          temp_b4_32_27_i;
wire signed [`CalcTempBus]          temp_b4_32_28_r;
wire signed [`CalcTempBus]          temp_b4_32_28_i;
wire signed [`CalcTempBus]          temp_b4_32_29_r;
wire signed [`CalcTempBus]          temp_b4_32_29_i;
wire signed [`CalcTempBus]          temp_b4_32_30_r;
wire signed [`CalcTempBus]          temp_b4_32_30_i;
wire signed [`CalcTempBus]          temp_b4_32_31_r;
wire signed [`CalcTempBus]          temp_b4_32_31_i;
wire signed [`CalcTempBus]          temp_b4_32_32_r;
wire signed [`CalcTempBus]          temp_b4_32_32_i;
wire signed [`CalcTempBus]          temp_b5_1_1_r;
wire signed [`CalcTempBus]          temp_b5_1_1_i;
wire signed [`CalcTempBus]          temp_b5_1_2_r;
wire signed [`CalcTempBus]          temp_b5_1_2_i;
wire signed [`CalcTempBus]          temp_b5_1_3_r;
wire signed [`CalcTempBus]          temp_b5_1_3_i;
wire signed [`CalcTempBus]          temp_b5_1_4_r;
wire signed [`CalcTempBus]          temp_b5_1_4_i;
wire signed [`CalcTempBus]          temp_b5_1_5_r;
wire signed [`CalcTempBus]          temp_b5_1_5_i;
wire signed [`CalcTempBus]          temp_b5_1_6_r;
wire signed [`CalcTempBus]          temp_b5_1_6_i;
wire signed [`CalcTempBus]          temp_b5_1_7_r;
wire signed [`CalcTempBus]          temp_b5_1_7_i;
wire signed [`CalcTempBus]          temp_b5_1_8_r;
wire signed [`CalcTempBus]          temp_b5_1_8_i;
wire signed [`CalcTempBus]          temp_b5_1_9_r;
wire signed [`CalcTempBus]          temp_b5_1_9_i;
wire signed [`CalcTempBus]          temp_b5_1_10_r;
wire signed [`CalcTempBus]          temp_b5_1_10_i;
wire signed [`CalcTempBus]          temp_b5_1_11_r;
wire signed [`CalcTempBus]          temp_b5_1_11_i;
wire signed [`CalcTempBus]          temp_b5_1_12_r;
wire signed [`CalcTempBus]          temp_b5_1_12_i;
wire signed [`CalcTempBus]          temp_b5_1_13_r;
wire signed [`CalcTempBus]          temp_b5_1_13_i;
wire signed [`CalcTempBus]          temp_b5_1_14_r;
wire signed [`CalcTempBus]          temp_b5_1_14_i;
wire signed [`CalcTempBus]          temp_b5_1_15_r;
wire signed [`CalcTempBus]          temp_b5_1_15_i;
wire signed [`CalcTempBus]          temp_b5_1_16_r;
wire signed [`CalcTempBus]          temp_b5_1_16_i;
wire signed [`CalcTempBus]          temp_b5_1_17_r;
wire signed [`CalcTempBus]          temp_b5_1_17_i;
wire signed [`CalcTempBus]          temp_b5_1_18_r;
wire signed [`CalcTempBus]          temp_b5_1_18_i;
wire signed [`CalcTempBus]          temp_b5_1_19_r;
wire signed [`CalcTempBus]          temp_b5_1_19_i;
wire signed [`CalcTempBus]          temp_b5_1_20_r;
wire signed [`CalcTempBus]          temp_b5_1_20_i;
wire signed [`CalcTempBus]          temp_b5_1_21_r;
wire signed [`CalcTempBus]          temp_b5_1_21_i;
wire signed [`CalcTempBus]          temp_b5_1_22_r;
wire signed [`CalcTempBus]          temp_b5_1_22_i;
wire signed [`CalcTempBus]          temp_b5_1_23_r;
wire signed [`CalcTempBus]          temp_b5_1_23_i;
wire signed [`CalcTempBus]          temp_b5_1_24_r;
wire signed [`CalcTempBus]          temp_b5_1_24_i;
wire signed [`CalcTempBus]          temp_b5_1_25_r;
wire signed [`CalcTempBus]          temp_b5_1_25_i;
wire signed [`CalcTempBus]          temp_b5_1_26_r;
wire signed [`CalcTempBus]          temp_b5_1_26_i;
wire signed [`CalcTempBus]          temp_b5_1_27_r;
wire signed [`CalcTempBus]          temp_b5_1_27_i;
wire signed [`CalcTempBus]          temp_b5_1_28_r;
wire signed [`CalcTempBus]          temp_b5_1_28_i;
wire signed [`CalcTempBus]          temp_b5_1_29_r;
wire signed [`CalcTempBus]          temp_b5_1_29_i;
wire signed [`CalcTempBus]          temp_b5_1_30_r;
wire signed [`CalcTempBus]          temp_b5_1_30_i;
wire signed [`CalcTempBus]          temp_b5_1_31_r;
wire signed [`CalcTempBus]          temp_b5_1_31_i;
wire signed [`CalcTempBus]          temp_b5_1_32_r;
wire signed [`CalcTempBus]          temp_b5_1_32_i;
wire signed [`CalcTempBus]          temp_b5_2_1_r;
wire signed [`CalcTempBus]          temp_b5_2_1_i;
wire signed [`CalcTempBus]          temp_b5_2_2_r;
wire signed [`CalcTempBus]          temp_b5_2_2_i;
wire signed [`CalcTempBus]          temp_b5_2_3_r;
wire signed [`CalcTempBus]          temp_b5_2_3_i;
wire signed [`CalcTempBus]          temp_b5_2_4_r;
wire signed [`CalcTempBus]          temp_b5_2_4_i;
wire signed [`CalcTempBus]          temp_b5_2_5_r;
wire signed [`CalcTempBus]          temp_b5_2_5_i;
wire signed [`CalcTempBus]          temp_b5_2_6_r;
wire signed [`CalcTempBus]          temp_b5_2_6_i;
wire signed [`CalcTempBus]          temp_b5_2_7_r;
wire signed [`CalcTempBus]          temp_b5_2_7_i;
wire signed [`CalcTempBus]          temp_b5_2_8_r;
wire signed [`CalcTempBus]          temp_b5_2_8_i;
wire signed [`CalcTempBus]          temp_b5_2_9_r;
wire signed [`CalcTempBus]          temp_b5_2_9_i;
wire signed [`CalcTempBus]          temp_b5_2_10_r;
wire signed [`CalcTempBus]          temp_b5_2_10_i;
wire signed [`CalcTempBus]          temp_b5_2_11_r;
wire signed [`CalcTempBus]          temp_b5_2_11_i;
wire signed [`CalcTempBus]          temp_b5_2_12_r;
wire signed [`CalcTempBus]          temp_b5_2_12_i;
wire signed [`CalcTempBus]          temp_b5_2_13_r;
wire signed [`CalcTempBus]          temp_b5_2_13_i;
wire signed [`CalcTempBus]          temp_b5_2_14_r;
wire signed [`CalcTempBus]          temp_b5_2_14_i;
wire signed [`CalcTempBus]          temp_b5_2_15_r;
wire signed [`CalcTempBus]          temp_b5_2_15_i;
wire signed [`CalcTempBus]          temp_b5_2_16_r;
wire signed [`CalcTempBus]          temp_b5_2_16_i;
wire signed [`CalcTempBus]          temp_b5_2_17_r;
wire signed [`CalcTempBus]          temp_b5_2_17_i;
wire signed [`CalcTempBus]          temp_b5_2_18_r;
wire signed [`CalcTempBus]          temp_b5_2_18_i;
wire signed [`CalcTempBus]          temp_b5_2_19_r;
wire signed [`CalcTempBus]          temp_b5_2_19_i;
wire signed [`CalcTempBus]          temp_b5_2_20_r;
wire signed [`CalcTempBus]          temp_b5_2_20_i;
wire signed [`CalcTempBus]          temp_b5_2_21_r;
wire signed [`CalcTempBus]          temp_b5_2_21_i;
wire signed [`CalcTempBus]          temp_b5_2_22_r;
wire signed [`CalcTempBus]          temp_b5_2_22_i;
wire signed [`CalcTempBus]          temp_b5_2_23_r;
wire signed [`CalcTempBus]          temp_b5_2_23_i;
wire signed [`CalcTempBus]          temp_b5_2_24_r;
wire signed [`CalcTempBus]          temp_b5_2_24_i;
wire signed [`CalcTempBus]          temp_b5_2_25_r;
wire signed [`CalcTempBus]          temp_b5_2_25_i;
wire signed [`CalcTempBus]          temp_b5_2_26_r;
wire signed [`CalcTempBus]          temp_b5_2_26_i;
wire signed [`CalcTempBus]          temp_b5_2_27_r;
wire signed [`CalcTempBus]          temp_b5_2_27_i;
wire signed [`CalcTempBus]          temp_b5_2_28_r;
wire signed [`CalcTempBus]          temp_b5_2_28_i;
wire signed [`CalcTempBus]          temp_b5_2_29_r;
wire signed [`CalcTempBus]          temp_b5_2_29_i;
wire signed [`CalcTempBus]          temp_b5_2_30_r;
wire signed [`CalcTempBus]          temp_b5_2_30_i;
wire signed [`CalcTempBus]          temp_b5_2_31_r;
wire signed [`CalcTempBus]          temp_b5_2_31_i;
wire signed [`CalcTempBus]          temp_b5_2_32_r;
wire signed [`CalcTempBus]          temp_b5_2_32_i;
wire signed [`CalcTempBus]          temp_b5_3_1_r;
wire signed [`CalcTempBus]          temp_b5_3_1_i;
wire signed [`CalcTempBus]          temp_b5_3_2_r;
wire signed [`CalcTempBus]          temp_b5_3_2_i;
wire signed [`CalcTempBus]          temp_b5_3_3_r;
wire signed [`CalcTempBus]          temp_b5_3_3_i;
wire signed [`CalcTempBus]          temp_b5_3_4_r;
wire signed [`CalcTempBus]          temp_b5_3_4_i;
wire signed [`CalcTempBus]          temp_b5_3_5_r;
wire signed [`CalcTempBus]          temp_b5_3_5_i;
wire signed [`CalcTempBus]          temp_b5_3_6_r;
wire signed [`CalcTempBus]          temp_b5_3_6_i;
wire signed [`CalcTempBus]          temp_b5_3_7_r;
wire signed [`CalcTempBus]          temp_b5_3_7_i;
wire signed [`CalcTempBus]          temp_b5_3_8_r;
wire signed [`CalcTempBus]          temp_b5_3_8_i;
wire signed [`CalcTempBus]          temp_b5_3_9_r;
wire signed [`CalcTempBus]          temp_b5_3_9_i;
wire signed [`CalcTempBus]          temp_b5_3_10_r;
wire signed [`CalcTempBus]          temp_b5_3_10_i;
wire signed [`CalcTempBus]          temp_b5_3_11_r;
wire signed [`CalcTempBus]          temp_b5_3_11_i;
wire signed [`CalcTempBus]          temp_b5_3_12_r;
wire signed [`CalcTempBus]          temp_b5_3_12_i;
wire signed [`CalcTempBus]          temp_b5_3_13_r;
wire signed [`CalcTempBus]          temp_b5_3_13_i;
wire signed [`CalcTempBus]          temp_b5_3_14_r;
wire signed [`CalcTempBus]          temp_b5_3_14_i;
wire signed [`CalcTempBus]          temp_b5_3_15_r;
wire signed [`CalcTempBus]          temp_b5_3_15_i;
wire signed [`CalcTempBus]          temp_b5_3_16_r;
wire signed [`CalcTempBus]          temp_b5_3_16_i;
wire signed [`CalcTempBus]          temp_b5_3_17_r;
wire signed [`CalcTempBus]          temp_b5_3_17_i;
wire signed [`CalcTempBus]          temp_b5_3_18_r;
wire signed [`CalcTempBus]          temp_b5_3_18_i;
wire signed [`CalcTempBus]          temp_b5_3_19_r;
wire signed [`CalcTempBus]          temp_b5_3_19_i;
wire signed [`CalcTempBus]          temp_b5_3_20_r;
wire signed [`CalcTempBus]          temp_b5_3_20_i;
wire signed [`CalcTempBus]          temp_b5_3_21_r;
wire signed [`CalcTempBus]          temp_b5_3_21_i;
wire signed [`CalcTempBus]          temp_b5_3_22_r;
wire signed [`CalcTempBus]          temp_b5_3_22_i;
wire signed [`CalcTempBus]          temp_b5_3_23_r;
wire signed [`CalcTempBus]          temp_b5_3_23_i;
wire signed [`CalcTempBus]          temp_b5_3_24_r;
wire signed [`CalcTempBus]          temp_b5_3_24_i;
wire signed [`CalcTempBus]          temp_b5_3_25_r;
wire signed [`CalcTempBus]          temp_b5_3_25_i;
wire signed [`CalcTempBus]          temp_b5_3_26_r;
wire signed [`CalcTempBus]          temp_b5_3_26_i;
wire signed [`CalcTempBus]          temp_b5_3_27_r;
wire signed [`CalcTempBus]          temp_b5_3_27_i;
wire signed [`CalcTempBus]          temp_b5_3_28_r;
wire signed [`CalcTempBus]          temp_b5_3_28_i;
wire signed [`CalcTempBus]          temp_b5_3_29_r;
wire signed [`CalcTempBus]          temp_b5_3_29_i;
wire signed [`CalcTempBus]          temp_b5_3_30_r;
wire signed [`CalcTempBus]          temp_b5_3_30_i;
wire signed [`CalcTempBus]          temp_b5_3_31_r;
wire signed [`CalcTempBus]          temp_b5_3_31_i;
wire signed [`CalcTempBus]          temp_b5_3_32_r;
wire signed [`CalcTempBus]          temp_b5_3_32_i;
wire signed [`CalcTempBus]          temp_b5_4_1_r;
wire signed [`CalcTempBus]          temp_b5_4_1_i;
wire signed [`CalcTempBus]          temp_b5_4_2_r;
wire signed [`CalcTempBus]          temp_b5_4_2_i;
wire signed [`CalcTempBus]          temp_b5_4_3_r;
wire signed [`CalcTempBus]          temp_b5_4_3_i;
wire signed [`CalcTempBus]          temp_b5_4_4_r;
wire signed [`CalcTempBus]          temp_b5_4_4_i;
wire signed [`CalcTempBus]          temp_b5_4_5_r;
wire signed [`CalcTempBus]          temp_b5_4_5_i;
wire signed [`CalcTempBus]          temp_b5_4_6_r;
wire signed [`CalcTempBus]          temp_b5_4_6_i;
wire signed [`CalcTempBus]          temp_b5_4_7_r;
wire signed [`CalcTempBus]          temp_b5_4_7_i;
wire signed [`CalcTempBus]          temp_b5_4_8_r;
wire signed [`CalcTempBus]          temp_b5_4_8_i;
wire signed [`CalcTempBus]          temp_b5_4_9_r;
wire signed [`CalcTempBus]          temp_b5_4_9_i;
wire signed [`CalcTempBus]          temp_b5_4_10_r;
wire signed [`CalcTempBus]          temp_b5_4_10_i;
wire signed [`CalcTempBus]          temp_b5_4_11_r;
wire signed [`CalcTempBus]          temp_b5_4_11_i;
wire signed [`CalcTempBus]          temp_b5_4_12_r;
wire signed [`CalcTempBus]          temp_b5_4_12_i;
wire signed [`CalcTempBus]          temp_b5_4_13_r;
wire signed [`CalcTempBus]          temp_b5_4_13_i;
wire signed [`CalcTempBus]          temp_b5_4_14_r;
wire signed [`CalcTempBus]          temp_b5_4_14_i;
wire signed [`CalcTempBus]          temp_b5_4_15_r;
wire signed [`CalcTempBus]          temp_b5_4_15_i;
wire signed [`CalcTempBus]          temp_b5_4_16_r;
wire signed [`CalcTempBus]          temp_b5_4_16_i;
wire signed [`CalcTempBus]          temp_b5_4_17_r;
wire signed [`CalcTempBus]          temp_b5_4_17_i;
wire signed [`CalcTempBus]          temp_b5_4_18_r;
wire signed [`CalcTempBus]          temp_b5_4_18_i;
wire signed [`CalcTempBus]          temp_b5_4_19_r;
wire signed [`CalcTempBus]          temp_b5_4_19_i;
wire signed [`CalcTempBus]          temp_b5_4_20_r;
wire signed [`CalcTempBus]          temp_b5_4_20_i;
wire signed [`CalcTempBus]          temp_b5_4_21_r;
wire signed [`CalcTempBus]          temp_b5_4_21_i;
wire signed [`CalcTempBus]          temp_b5_4_22_r;
wire signed [`CalcTempBus]          temp_b5_4_22_i;
wire signed [`CalcTempBus]          temp_b5_4_23_r;
wire signed [`CalcTempBus]          temp_b5_4_23_i;
wire signed [`CalcTempBus]          temp_b5_4_24_r;
wire signed [`CalcTempBus]          temp_b5_4_24_i;
wire signed [`CalcTempBus]          temp_b5_4_25_r;
wire signed [`CalcTempBus]          temp_b5_4_25_i;
wire signed [`CalcTempBus]          temp_b5_4_26_r;
wire signed [`CalcTempBus]          temp_b5_4_26_i;
wire signed [`CalcTempBus]          temp_b5_4_27_r;
wire signed [`CalcTempBus]          temp_b5_4_27_i;
wire signed [`CalcTempBus]          temp_b5_4_28_r;
wire signed [`CalcTempBus]          temp_b5_4_28_i;
wire signed [`CalcTempBus]          temp_b5_4_29_r;
wire signed [`CalcTempBus]          temp_b5_4_29_i;
wire signed [`CalcTempBus]          temp_b5_4_30_r;
wire signed [`CalcTempBus]          temp_b5_4_30_i;
wire signed [`CalcTempBus]          temp_b5_4_31_r;
wire signed [`CalcTempBus]          temp_b5_4_31_i;
wire signed [`CalcTempBus]          temp_b5_4_32_r;
wire signed [`CalcTempBus]          temp_b5_4_32_i;
wire signed [`CalcTempBus]          temp_b5_5_1_r;
wire signed [`CalcTempBus]          temp_b5_5_1_i;
wire signed [`CalcTempBus]          temp_b5_5_2_r;
wire signed [`CalcTempBus]          temp_b5_5_2_i;
wire signed [`CalcTempBus]          temp_b5_5_3_r;
wire signed [`CalcTempBus]          temp_b5_5_3_i;
wire signed [`CalcTempBus]          temp_b5_5_4_r;
wire signed [`CalcTempBus]          temp_b5_5_4_i;
wire signed [`CalcTempBus]          temp_b5_5_5_r;
wire signed [`CalcTempBus]          temp_b5_5_5_i;
wire signed [`CalcTempBus]          temp_b5_5_6_r;
wire signed [`CalcTempBus]          temp_b5_5_6_i;
wire signed [`CalcTempBus]          temp_b5_5_7_r;
wire signed [`CalcTempBus]          temp_b5_5_7_i;
wire signed [`CalcTempBus]          temp_b5_5_8_r;
wire signed [`CalcTempBus]          temp_b5_5_8_i;
wire signed [`CalcTempBus]          temp_b5_5_9_r;
wire signed [`CalcTempBus]          temp_b5_5_9_i;
wire signed [`CalcTempBus]          temp_b5_5_10_r;
wire signed [`CalcTempBus]          temp_b5_5_10_i;
wire signed [`CalcTempBus]          temp_b5_5_11_r;
wire signed [`CalcTempBus]          temp_b5_5_11_i;
wire signed [`CalcTempBus]          temp_b5_5_12_r;
wire signed [`CalcTempBus]          temp_b5_5_12_i;
wire signed [`CalcTempBus]          temp_b5_5_13_r;
wire signed [`CalcTempBus]          temp_b5_5_13_i;
wire signed [`CalcTempBus]          temp_b5_5_14_r;
wire signed [`CalcTempBus]          temp_b5_5_14_i;
wire signed [`CalcTempBus]          temp_b5_5_15_r;
wire signed [`CalcTempBus]          temp_b5_5_15_i;
wire signed [`CalcTempBus]          temp_b5_5_16_r;
wire signed [`CalcTempBus]          temp_b5_5_16_i;
wire signed [`CalcTempBus]          temp_b5_5_17_r;
wire signed [`CalcTempBus]          temp_b5_5_17_i;
wire signed [`CalcTempBus]          temp_b5_5_18_r;
wire signed [`CalcTempBus]          temp_b5_5_18_i;
wire signed [`CalcTempBus]          temp_b5_5_19_r;
wire signed [`CalcTempBus]          temp_b5_5_19_i;
wire signed [`CalcTempBus]          temp_b5_5_20_r;
wire signed [`CalcTempBus]          temp_b5_5_20_i;
wire signed [`CalcTempBus]          temp_b5_5_21_r;
wire signed [`CalcTempBus]          temp_b5_5_21_i;
wire signed [`CalcTempBus]          temp_b5_5_22_r;
wire signed [`CalcTempBus]          temp_b5_5_22_i;
wire signed [`CalcTempBus]          temp_b5_5_23_r;
wire signed [`CalcTempBus]          temp_b5_5_23_i;
wire signed [`CalcTempBus]          temp_b5_5_24_r;
wire signed [`CalcTempBus]          temp_b5_5_24_i;
wire signed [`CalcTempBus]          temp_b5_5_25_r;
wire signed [`CalcTempBus]          temp_b5_5_25_i;
wire signed [`CalcTempBus]          temp_b5_5_26_r;
wire signed [`CalcTempBus]          temp_b5_5_26_i;
wire signed [`CalcTempBus]          temp_b5_5_27_r;
wire signed [`CalcTempBus]          temp_b5_5_27_i;
wire signed [`CalcTempBus]          temp_b5_5_28_r;
wire signed [`CalcTempBus]          temp_b5_5_28_i;
wire signed [`CalcTempBus]          temp_b5_5_29_r;
wire signed [`CalcTempBus]          temp_b5_5_29_i;
wire signed [`CalcTempBus]          temp_b5_5_30_r;
wire signed [`CalcTempBus]          temp_b5_5_30_i;
wire signed [`CalcTempBus]          temp_b5_5_31_r;
wire signed [`CalcTempBus]          temp_b5_5_31_i;
wire signed [`CalcTempBus]          temp_b5_5_32_r;
wire signed [`CalcTempBus]          temp_b5_5_32_i;
wire signed [`CalcTempBus]          temp_b5_6_1_r;
wire signed [`CalcTempBus]          temp_b5_6_1_i;
wire signed [`CalcTempBus]          temp_b5_6_2_r;
wire signed [`CalcTempBus]          temp_b5_6_2_i;
wire signed [`CalcTempBus]          temp_b5_6_3_r;
wire signed [`CalcTempBus]          temp_b5_6_3_i;
wire signed [`CalcTempBus]          temp_b5_6_4_r;
wire signed [`CalcTempBus]          temp_b5_6_4_i;
wire signed [`CalcTempBus]          temp_b5_6_5_r;
wire signed [`CalcTempBus]          temp_b5_6_5_i;
wire signed [`CalcTempBus]          temp_b5_6_6_r;
wire signed [`CalcTempBus]          temp_b5_6_6_i;
wire signed [`CalcTempBus]          temp_b5_6_7_r;
wire signed [`CalcTempBus]          temp_b5_6_7_i;
wire signed [`CalcTempBus]          temp_b5_6_8_r;
wire signed [`CalcTempBus]          temp_b5_6_8_i;
wire signed [`CalcTempBus]          temp_b5_6_9_r;
wire signed [`CalcTempBus]          temp_b5_6_9_i;
wire signed [`CalcTempBus]          temp_b5_6_10_r;
wire signed [`CalcTempBus]          temp_b5_6_10_i;
wire signed [`CalcTempBus]          temp_b5_6_11_r;
wire signed [`CalcTempBus]          temp_b5_6_11_i;
wire signed [`CalcTempBus]          temp_b5_6_12_r;
wire signed [`CalcTempBus]          temp_b5_6_12_i;
wire signed [`CalcTempBus]          temp_b5_6_13_r;
wire signed [`CalcTempBus]          temp_b5_6_13_i;
wire signed [`CalcTempBus]          temp_b5_6_14_r;
wire signed [`CalcTempBus]          temp_b5_6_14_i;
wire signed [`CalcTempBus]          temp_b5_6_15_r;
wire signed [`CalcTempBus]          temp_b5_6_15_i;
wire signed [`CalcTempBus]          temp_b5_6_16_r;
wire signed [`CalcTempBus]          temp_b5_6_16_i;
wire signed [`CalcTempBus]          temp_b5_6_17_r;
wire signed [`CalcTempBus]          temp_b5_6_17_i;
wire signed [`CalcTempBus]          temp_b5_6_18_r;
wire signed [`CalcTempBus]          temp_b5_6_18_i;
wire signed [`CalcTempBus]          temp_b5_6_19_r;
wire signed [`CalcTempBus]          temp_b5_6_19_i;
wire signed [`CalcTempBus]          temp_b5_6_20_r;
wire signed [`CalcTempBus]          temp_b5_6_20_i;
wire signed [`CalcTempBus]          temp_b5_6_21_r;
wire signed [`CalcTempBus]          temp_b5_6_21_i;
wire signed [`CalcTempBus]          temp_b5_6_22_r;
wire signed [`CalcTempBus]          temp_b5_6_22_i;
wire signed [`CalcTempBus]          temp_b5_6_23_r;
wire signed [`CalcTempBus]          temp_b5_6_23_i;
wire signed [`CalcTempBus]          temp_b5_6_24_r;
wire signed [`CalcTempBus]          temp_b5_6_24_i;
wire signed [`CalcTempBus]          temp_b5_6_25_r;
wire signed [`CalcTempBus]          temp_b5_6_25_i;
wire signed [`CalcTempBus]          temp_b5_6_26_r;
wire signed [`CalcTempBus]          temp_b5_6_26_i;
wire signed [`CalcTempBus]          temp_b5_6_27_r;
wire signed [`CalcTempBus]          temp_b5_6_27_i;
wire signed [`CalcTempBus]          temp_b5_6_28_r;
wire signed [`CalcTempBus]          temp_b5_6_28_i;
wire signed [`CalcTempBus]          temp_b5_6_29_r;
wire signed [`CalcTempBus]          temp_b5_6_29_i;
wire signed [`CalcTempBus]          temp_b5_6_30_r;
wire signed [`CalcTempBus]          temp_b5_6_30_i;
wire signed [`CalcTempBus]          temp_b5_6_31_r;
wire signed [`CalcTempBus]          temp_b5_6_31_i;
wire signed [`CalcTempBus]          temp_b5_6_32_r;
wire signed [`CalcTempBus]          temp_b5_6_32_i;
wire signed [`CalcTempBus]          temp_b5_7_1_r;
wire signed [`CalcTempBus]          temp_b5_7_1_i;
wire signed [`CalcTempBus]          temp_b5_7_2_r;
wire signed [`CalcTempBus]          temp_b5_7_2_i;
wire signed [`CalcTempBus]          temp_b5_7_3_r;
wire signed [`CalcTempBus]          temp_b5_7_3_i;
wire signed [`CalcTempBus]          temp_b5_7_4_r;
wire signed [`CalcTempBus]          temp_b5_7_4_i;
wire signed [`CalcTempBus]          temp_b5_7_5_r;
wire signed [`CalcTempBus]          temp_b5_7_5_i;
wire signed [`CalcTempBus]          temp_b5_7_6_r;
wire signed [`CalcTempBus]          temp_b5_7_6_i;
wire signed [`CalcTempBus]          temp_b5_7_7_r;
wire signed [`CalcTempBus]          temp_b5_7_7_i;
wire signed [`CalcTempBus]          temp_b5_7_8_r;
wire signed [`CalcTempBus]          temp_b5_7_8_i;
wire signed [`CalcTempBus]          temp_b5_7_9_r;
wire signed [`CalcTempBus]          temp_b5_7_9_i;
wire signed [`CalcTempBus]          temp_b5_7_10_r;
wire signed [`CalcTempBus]          temp_b5_7_10_i;
wire signed [`CalcTempBus]          temp_b5_7_11_r;
wire signed [`CalcTempBus]          temp_b5_7_11_i;
wire signed [`CalcTempBus]          temp_b5_7_12_r;
wire signed [`CalcTempBus]          temp_b5_7_12_i;
wire signed [`CalcTempBus]          temp_b5_7_13_r;
wire signed [`CalcTempBus]          temp_b5_7_13_i;
wire signed [`CalcTempBus]          temp_b5_7_14_r;
wire signed [`CalcTempBus]          temp_b5_7_14_i;
wire signed [`CalcTempBus]          temp_b5_7_15_r;
wire signed [`CalcTempBus]          temp_b5_7_15_i;
wire signed [`CalcTempBus]          temp_b5_7_16_r;
wire signed [`CalcTempBus]          temp_b5_7_16_i;
wire signed [`CalcTempBus]          temp_b5_7_17_r;
wire signed [`CalcTempBus]          temp_b5_7_17_i;
wire signed [`CalcTempBus]          temp_b5_7_18_r;
wire signed [`CalcTempBus]          temp_b5_7_18_i;
wire signed [`CalcTempBus]          temp_b5_7_19_r;
wire signed [`CalcTempBus]          temp_b5_7_19_i;
wire signed [`CalcTempBus]          temp_b5_7_20_r;
wire signed [`CalcTempBus]          temp_b5_7_20_i;
wire signed [`CalcTempBus]          temp_b5_7_21_r;
wire signed [`CalcTempBus]          temp_b5_7_21_i;
wire signed [`CalcTempBus]          temp_b5_7_22_r;
wire signed [`CalcTempBus]          temp_b5_7_22_i;
wire signed [`CalcTempBus]          temp_b5_7_23_r;
wire signed [`CalcTempBus]          temp_b5_7_23_i;
wire signed [`CalcTempBus]          temp_b5_7_24_r;
wire signed [`CalcTempBus]          temp_b5_7_24_i;
wire signed [`CalcTempBus]          temp_b5_7_25_r;
wire signed [`CalcTempBus]          temp_b5_7_25_i;
wire signed [`CalcTempBus]          temp_b5_7_26_r;
wire signed [`CalcTempBus]          temp_b5_7_26_i;
wire signed [`CalcTempBus]          temp_b5_7_27_r;
wire signed [`CalcTempBus]          temp_b5_7_27_i;
wire signed [`CalcTempBus]          temp_b5_7_28_r;
wire signed [`CalcTempBus]          temp_b5_7_28_i;
wire signed [`CalcTempBus]          temp_b5_7_29_r;
wire signed [`CalcTempBus]          temp_b5_7_29_i;
wire signed [`CalcTempBus]          temp_b5_7_30_r;
wire signed [`CalcTempBus]          temp_b5_7_30_i;
wire signed [`CalcTempBus]          temp_b5_7_31_r;
wire signed [`CalcTempBus]          temp_b5_7_31_i;
wire signed [`CalcTempBus]          temp_b5_7_32_r;
wire signed [`CalcTempBus]          temp_b5_7_32_i;
wire signed [`CalcTempBus]          temp_b5_8_1_r;
wire signed [`CalcTempBus]          temp_b5_8_1_i;
wire signed [`CalcTempBus]          temp_b5_8_2_r;
wire signed [`CalcTempBus]          temp_b5_8_2_i;
wire signed [`CalcTempBus]          temp_b5_8_3_r;
wire signed [`CalcTempBus]          temp_b5_8_3_i;
wire signed [`CalcTempBus]          temp_b5_8_4_r;
wire signed [`CalcTempBus]          temp_b5_8_4_i;
wire signed [`CalcTempBus]          temp_b5_8_5_r;
wire signed [`CalcTempBus]          temp_b5_8_5_i;
wire signed [`CalcTempBus]          temp_b5_8_6_r;
wire signed [`CalcTempBus]          temp_b5_8_6_i;
wire signed [`CalcTempBus]          temp_b5_8_7_r;
wire signed [`CalcTempBus]          temp_b5_8_7_i;
wire signed [`CalcTempBus]          temp_b5_8_8_r;
wire signed [`CalcTempBus]          temp_b5_8_8_i;
wire signed [`CalcTempBus]          temp_b5_8_9_r;
wire signed [`CalcTempBus]          temp_b5_8_9_i;
wire signed [`CalcTempBus]          temp_b5_8_10_r;
wire signed [`CalcTempBus]          temp_b5_8_10_i;
wire signed [`CalcTempBus]          temp_b5_8_11_r;
wire signed [`CalcTempBus]          temp_b5_8_11_i;
wire signed [`CalcTempBus]          temp_b5_8_12_r;
wire signed [`CalcTempBus]          temp_b5_8_12_i;
wire signed [`CalcTempBus]          temp_b5_8_13_r;
wire signed [`CalcTempBus]          temp_b5_8_13_i;
wire signed [`CalcTempBus]          temp_b5_8_14_r;
wire signed [`CalcTempBus]          temp_b5_8_14_i;
wire signed [`CalcTempBus]          temp_b5_8_15_r;
wire signed [`CalcTempBus]          temp_b5_8_15_i;
wire signed [`CalcTempBus]          temp_b5_8_16_r;
wire signed [`CalcTempBus]          temp_b5_8_16_i;
wire signed [`CalcTempBus]          temp_b5_8_17_r;
wire signed [`CalcTempBus]          temp_b5_8_17_i;
wire signed [`CalcTempBus]          temp_b5_8_18_r;
wire signed [`CalcTempBus]          temp_b5_8_18_i;
wire signed [`CalcTempBus]          temp_b5_8_19_r;
wire signed [`CalcTempBus]          temp_b5_8_19_i;
wire signed [`CalcTempBus]          temp_b5_8_20_r;
wire signed [`CalcTempBus]          temp_b5_8_20_i;
wire signed [`CalcTempBus]          temp_b5_8_21_r;
wire signed [`CalcTempBus]          temp_b5_8_21_i;
wire signed [`CalcTempBus]          temp_b5_8_22_r;
wire signed [`CalcTempBus]          temp_b5_8_22_i;
wire signed [`CalcTempBus]          temp_b5_8_23_r;
wire signed [`CalcTempBus]          temp_b5_8_23_i;
wire signed [`CalcTempBus]          temp_b5_8_24_r;
wire signed [`CalcTempBus]          temp_b5_8_24_i;
wire signed [`CalcTempBus]          temp_b5_8_25_r;
wire signed [`CalcTempBus]          temp_b5_8_25_i;
wire signed [`CalcTempBus]          temp_b5_8_26_r;
wire signed [`CalcTempBus]          temp_b5_8_26_i;
wire signed [`CalcTempBus]          temp_b5_8_27_r;
wire signed [`CalcTempBus]          temp_b5_8_27_i;
wire signed [`CalcTempBus]          temp_b5_8_28_r;
wire signed [`CalcTempBus]          temp_b5_8_28_i;
wire signed [`CalcTempBus]          temp_b5_8_29_r;
wire signed [`CalcTempBus]          temp_b5_8_29_i;
wire signed [`CalcTempBus]          temp_b5_8_30_r;
wire signed [`CalcTempBus]          temp_b5_8_30_i;
wire signed [`CalcTempBus]          temp_b5_8_31_r;
wire signed [`CalcTempBus]          temp_b5_8_31_i;
wire signed [`CalcTempBus]          temp_b5_8_32_r;
wire signed [`CalcTempBus]          temp_b5_8_32_i;
wire signed [`CalcTempBus]          temp_b5_9_1_r;
wire signed [`CalcTempBus]          temp_b5_9_1_i;
wire signed [`CalcTempBus]          temp_b5_9_2_r;
wire signed [`CalcTempBus]          temp_b5_9_2_i;
wire signed [`CalcTempBus]          temp_b5_9_3_r;
wire signed [`CalcTempBus]          temp_b5_9_3_i;
wire signed [`CalcTempBus]          temp_b5_9_4_r;
wire signed [`CalcTempBus]          temp_b5_9_4_i;
wire signed [`CalcTempBus]          temp_b5_9_5_r;
wire signed [`CalcTempBus]          temp_b5_9_5_i;
wire signed [`CalcTempBus]          temp_b5_9_6_r;
wire signed [`CalcTempBus]          temp_b5_9_6_i;
wire signed [`CalcTempBus]          temp_b5_9_7_r;
wire signed [`CalcTempBus]          temp_b5_9_7_i;
wire signed [`CalcTempBus]          temp_b5_9_8_r;
wire signed [`CalcTempBus]          temp_b5_9_8_i;
wire signed [`CalcTempBus]          temp_b5_9_9_r;
wire signed [`CalcTempBus]          temp_b5_9_9_i;
wire signed [`CalcTempBus]          temp_b5_9_10_r;
wire signed [`CalcTempBus]          temp_b5_9_10_i;
wire signed [`CalcTempBus]          temp_b5_9_11_r;
wire signed [`CalcTempBus]          temp_b5_9_11_i;
wire signed [`CalcTempBus]          temp_b5_9_12_r;
wire signed [`CalcTempBus]          temp_b5_9_12_i;
wire signed [`CalcTempBus]          temp_b5_9_13_r;
wire signed [`CalcTempBus]          temp_b5_9_13_i;
wire signed [`CalcTempBus]          temp_b5_9_14_r;
wire signed [`CalcTempBus]          temp_b5_9_14_i;
wire signed [`CalcTempBus]          temp_b5_9_15_r;
wire signed [`CalcTempBus]          temp_b5_9_15_i;
wire signed [`CalcTempBus]          temp_b5_9_16_r;
wire signed [`CalcTempBus]          temp_b5_9_16_i;
wire signed [`CalcTempBus]          temp_b5_9_17_r;
wire signed [`CalcTempBus]          temp_b5_9_17_i;
wire signed [`CalcTempBus]          temp_b5_9_18_r;
wire signed [`CalcTempBus]          temp_b5_9_18_i;
wire signed [`CalcTempBus]          temp_b5_9_19_r;
wire signed [`CalcTempBus]          temp_b5_9_19_i;
wire signed [`CalcTempBus]          temp_b5_9_20_r;
wire signed [`CalcTempBus]          temp_b5_9_20_i;
wire signed [`CalcTempBus]          temp_b5_9_21_r;
wire signed [`CalcTempBus]          temp_b5_9_21_i;
wire signed [`CalcTempBus]          temp_b5_9_22_r;
wire signed [`CalcTempBus]          temp_b5_9_22_i;
wire signed [`CalcTempBus]          temp_b5_9_23_r;
wire signed [`CalcTempBus]          temp_b5_9_23_i;
wire signed [`CalcTempBus]          temp_b5_9_24_r;
wire signed [`CalcTempBus]          temp_b5_9_24_i;
wire signed [`CalcTempBus]          temp_b5_9_25_r;
wire signed [`CalcTempBus]          temp_b5_9_25_i;
wire signed [`CalcTempBus]          temp_b5_9_26_r;
wire signed [`CalcTempBus]          temp_b5_9_26_i;
wire signed [`CalcTempBus]          temp_b5_9_27_r;
wire signed [`CalcTempBus]          temp_b5_9_27_i;
wire signed [`CalcTempBus]          temp_b5_9_28_r;
wire signed [`CalcTempBus]          temp_b5_9_28_i;
wire signed [`CalcTempBus]          temp_b5_9_29_r;
wire signed [`CalcTempBus]          temp_b5_9_29_i;
wire signed [`CalcTempBus]          temp_b5_9_30_r;
wire signed [`CalcTempBus]          temp_b5_9_30_i;
wire signed [`CalcTempBus]          temp_b5_9_31_r;
wire signed [`CalcTempBus]          temp_b5_9_31_i;
wire signed [`CalcTempBus]          temp_b5_9_32_r;
wire signed [`CalcTempBus]          temp_b5_9_32_i;
wire signed [`CalcTempBus]          temp_b5_10_1_r;
wire signed [`CalcTempBus]          temp_b5_10_1_i;
wire signed [`CalcTempBus]          temp_b5_10_2_r;
wire signed [`CalcTempBus]          temp_b5_10_2_i;
wire signed [`CalcTempBus]          temp_b5_10_3_r;
wire signed [`CalcTempBus]          temp_b5_10_3_i;
wire signed [`CalcTempBus]          temp_b5_10_4_r;
wire signed [`CalcTempBus]          temp_b5_10_4_i;
wire signed [`CalcTempBus]          temp_b5_10_5_r;
wire signed [`CalcTempBus]          temp_b5_10_5_i;
wire signed [`CalcTempBus]          temp_b5_10_6_r;
wire signed [`CalcTempBus]          temp_b5_10_6_i;
wire signed [`CalcTempBus]          temp_b5_10_7_r;
wire signed [`CalcTempBus]          temp_b5_10_7_i;
wire signed [`CalcTempBus]          temp_b5_10_8_r;
wire signed [`CalcTempBus]          temp_b5_10_8_i;
wire signed [`CalcTempBus]          temp_b5_10_9_r;
wire signed [`CalcTempBus]          temp_b5_10_9_i;
wire signed [`CalcTempBus]          temp_b5_10_10_r;
wire signed [`CalcTempBus]          temp_b5_10_10_i;
wire signed [`CalcTempBus]          temp_b5_10_11_r;
wire signed [`CalcTempBus]          temp_b5_10_11_i;
wire signed [`CalcTempBus]          temp_b5_10_12_r;
wire signed [`CalcTempBus]          temp_b5_10_12_i;
wire signed [`CalcTempBus]          temp_b5_10_13_r;
wire signed [`CalcTempBus]          temp_b5_10_13_i;
wire signed [`CalcTempBus]          temp_b5_10_14_r;
wire signed [`CalcTempBus]          temp_b5_10_14_i;
wire signed [`CalcTempBus]          temp_b5_10_15_r;
wire signed [`CalcTempBus]          temp_b5_10_15_i;
wire signed [`CalcTempBus]          temp_b5_10_16_r;
wire signed [`CalcTempBus]          temp_b5_10_16_i;
wire signed [`CalcTempBus]          temp_b5_10_17_r;
wire signed [`CalcTempBus]          temp_b5_10_17_i;
wire signed [`CalcTempBus]          temp_b5_10_18_r;
wire signed [`CalcTempBus]          temp_b5_10_18_i;
wire signed [`CalcTempBus]          temp_b5_10_19_r;
wire signed [`CalcTempBus]          temp_b5_10_19_i;
wire signed [`CalcTempBus]          temp_b5_10_20_r;
wire signed [`CalcTempBus]          temp_b5_10_20_i;
wire signed [`CalcTempBus]          temp_b5_10_21_r;
wire signed [`CalcTempBus]          temp_b5_10_21_i;
wire signed [`CalcTempBus]          temp_b5_10_22_r;
wire signed [`CalcTempBus]          temp_b5_10_22_i;
wire signed [`CalcTempBus]          temp_b5_10_23_r;
wire signed [`CalcTempBus]          temp_b5_10_23_i;
wire signed [`CalcTempBus]          temp_b5_10_24_r;
wire signed [`CalcTempBus]          temp_b5_10_24_i;
wire signed [`CalcTempBus]          temp_b5_10_25_r;
wire signed [`CalcTempBus]          temp_b5_10_25_i;
wire signed [`CalcTempBus]          temp_b5_10_26_r;
wire signed [`CalcTempBus]          temp_b5_10_26_i;
wire signed [`CalcTempBus]          temp_b5_10_27_r;
wire signed [`CalcTempBus]          temp_b5_10_27_i;
wire signed [`CalcTempBus]          temp_b5_10_28_r;
wire signed [`CalcTempBus]          temp_b5_10_28_i;
wire signed [`CalcTempBus]          temp_b5_10_29_r;
wire signed [`CalcTempBus]          temp_b5_10_29_i;
wire signed [`CalcTempBus]          temp_b5_10_30_r;
wire signed [`CalcTempBus]          temp_b5_10_30_i;
wire signed [`CalcTempBus]          temp_b5_10_31_r;
wire signed [`CalcTempBus]          temp_b5_10_31_i;
wire signed [`CalcTempBus]          temp_b5_10_32_r;
wire signed [`CalcTempBus]          temp_b5_10_32_i;
wire signed [`CalcTempBus]          temp_b5_11_1_r;
wire signed [`CalcTempBus]          temp_b5_11_1_i;
wire signed [`CalcTempBus]          temp_b5_11_2_r;
wire signed [`CalcTempBus]          temp_b5_11_2_i;
wire signed [`CalcTempBus]          temp_b5_11_3_r;
wire signed [`CalcTempBus]          temp_b5_11_3_i;
wire signed [`CalcTempBus]          temp_b5_11_4_r;
wire signed [`CalcTempBus]          temp_b5_11_4_i;
wire signed [`CalcTempBus]          temp_b5_11_5_r;
wire signed [`CalcTempBus]          temp_b5_11_5_i;
wire signed [`CalcTempBus]          temp_b5_11_6_r;
wire signed [`CalcTempBus]          temp_b5_11_6_i;
wire signed [`CalcTempBus]          temp_b5_11_7_r;
wire signed [`CalcTempBus]          temp_b5_11_7_i;
wire signed [`CalcTempBus]          temp_b5_11_8_r;
wire signed [`CalcTempBus]          temp_b5_11_8_i;
wire signed [`CalcTempBus]          temp_b5_11_9_r;
wire signed [`CalcTempBus]          temp_b5_11_9_i;
wire signed [`CalcTempBus]          temp_b5_11_10_r;
wire signed [`CalcTempBus]          temp_b5_11_10_i;
wire signed [`CalcTempBus]          temp_b5_11_11_r;
wire signed [`CalcTempBus]          temp_b5_11_11_i;
wire signed [`CalcTempBus]          temp_b5_11_12_r;
wire signed [`CalcTempBus]          temp_b5_11_12_i;
wire signed [`CalcTempBus]          temp_b5_11_13_r;
wire signed [`CalcTempBus]          temp_b5_11_13_i;
wire signed [`CalcTempBus]          temp_b5_11_14_r;
wire signed [`CalcTempBus]          temp_b5_11_14_i;
wire signed [`CalcTempBus]          temp_b5_11_15_r;
wire signed [`CalcTempBus]          temp_b5_11_15_i;
wire signed [`CalcTempBus]          temp_b5_11_16_r;
wire signed [`CalcTempBus]          temp_b5_11_16_i;
wire signed [`CalcTempBus]          temp_b5_11_17_r;
wire signed [`CalcTempBus]          temp_b5_11_17_i;
wire signed [`CalcTempBus]          temp_b5_11_18_r;
wire signed [`CalcTempBus]          temp_b5_11_18_i;
wire signed [`CalcTempBus]          temp_b5_11_19_r;
wire signed [`CalcTempBus]          temp_b5_11_19_i;
wire signed [`CalcTempBus]          temp_b5_11_20_r;
wire signed [`CalcTempBus]          temp_b5_11_20_i;
wire signed [`CalcTempBus]          temp_b5_11_21_r;
wire signed [`CalcTempBus]          temp_b5_11_21_i;
wire signed [`CalcTempBus]          temp_b5_11_22_r;
wire signed [`CalcTempBus]          temp_b5_11_22_i;
wire signed [`CalcTempBus]          temp_b5_11_23_r;
wire signed [`CalcTempBus]          temp_b5_11_23_i;
wire signed [`CalcTempBus]          temp_b5_11_24_r;
wire signed [`CalcTempBus]          temp_b5_11_24_i;
wire signed [`CalcTempBus]          temp_b5_11_25_r;
wire signed [`CalcTempBus]          temp_b5_11_25_i;
wire signed [`CalcTempBus]          temp_b5_11_26_r;
wire signed [`CalcTempBus]          temp_b5_11_26_i;
wire signed [`CalcTempBus]          temp_b5_11_27_r;
wire signed [`CalcTempBus]          temp_b5_11_27_i;
wire signed [`CalcTempBus]          temp_b5_11_28_r;
wire signed [`CalcTempBus]          temp_b5_11_28_i;
wire signed [`CalcTempBus]          temp_b5_11_29_r;
wire signed [`CalcTempBus]          temp_b5_11_29_i;
wire signed [`CalcTempBus]          temp_b5_11_30_r;
wire signed [`CalcTempBus]          temp_b5_11_30_i;
wire signed [`CalcTempBus]          temp_b5_11_31_r;
wire signed [`CalcTempBus]          temp_b5_11_31_i;
wire signed [`CalcTempBus]          temp_b5_11_32_r;
wire signed [`CalcTempBus]          temp_b5_11_32_i;
wire signed [`CalcTempBus]          temp_b5_12_1_r;
wire signed [`CalcTempBus]          temp_b5_12_1_i;
wire signed [`CalcTempBus]          temp_b5_12_2_r;
wire signed [`CalcTempBus]          temp_b5_12_2_i;
wire signed [`CalcTempBus]          temp_b5_12_3_r;
wire signed [`CalcTempBus]          temp_b5_12_3_i;
wire signed [`CalcTempBus]          temp_b5_12_4_r;
wire signed [`CalcTempBus]          temp_b5_12_4_i;
wire signed [`CalcTempBus]          temp_b5_12_5_r;
wire signed [`CalcTempBus]          temp_b5_12_5_i;
wire signed [`CalcTempBus]          temp_b5_12_6_r;
wire signed [`CalcTempBus]          temp_b5_12_6_i;
wire signed [`CalcTempBus]          temp_b5_12_7_r;
wire signed [`CalcTempBus]          temp_b5_12_7_i;
wire signed [`CalcTempBus]          temp_b5_12_8_r;
wire signed [`CalcTempBus]          temp_b5_12_8_i;
wire signed [`CalcTempBus]          temp_b5_12_9_r;
wire signed [`CalcTempBus]          temp_b5_12_9_i;
wire signed [`CalcTempBus]          temp_b5_12_10_r;
wire signed [`CalcTempBus]          temp_b5_12_10_i;
wire signed [`CalcTempBus]          temp_b5_12_11_r;
wire signed [`CalcTempBus]          temp_b5_12_11_i;
wire signed [`CalcTempBus]          temp_b5_12_12_r;
wire signed [`CalcTempBus]          temp_b5_12_12_i;
wire signed [`CalcTempBus]          temp_b5_12_13_r;
wire signed [`CalcTempBus]          temp_b5_12_13_i;
wire signed [`CalcTempBus]          temp_b5_12_14_r;
wire signed [`CalcTempBus]          temp_b5_12_14_i;
wire signed [`CalcTempBus]          temp_b5_12_15_r;
wire signed [`CalcTempBus]          temp_b5_12_15_i;
wire signed [`CalcTempBus]          temp_b5_12_16_r;
wire signed [`CalcTempBus]          temp_b5_12_16_i;
wire signed [`CalcTempBus]          temp_b5_12_17_r;
wire signed [`CalcTempBus]          temp_b5_12_17_i;
wire signed [`CalcTempBus]          temp_b5_12_18_r;
wire signed [`CalcTempBus]          temp_b5_12_18_i;
wire signed [`CalcTempBus]          temp_b5_12_19_r;
wire signed [`CalcTempBus]          temp_b5_12_19_i;
wire signed [`CalcTempBus]          temp_b5_12_20_r;
wire signed [`CalcTempBus]          temp_b5_12_20_i;
wire signed [`CalcTempBus]          temp_b5_12_21_r;
wire signed [`CalcTempBus]          temp_b5_12_21_i;
wire signed [`CalcTempBus]          temp_b5_12_22_r;
wire signed [`CalcTempBus]          temp_b5_12_22_i;
wire signed [`CalcTempBus]          temp_b5_12_23_r;
wire signed [`CalcTempBus]          temp_b5_12_23_i;
wire signed [`CalcTempBus]          temp_b5_12_24_r;
wire signed [`CalcTempBus]          temp_b5_12_24_i;
wire signed [`CalcTempBus]          temp_b5_12_25_r;
wire signed [`CalcTempBus]          temp_b5_12_25_i;
wire signed [`CalcTempBus]          temp_b5_12_26_r;
wire signed [`CalcTempBus]          temp_b5_12_26_i;
wire signed [`CalcTempBus]          temp_b5_12_27_r;
wire signed [`CalcTempBus]          temp_b5_12_27_i;
wire signed [`CalcTempBus]          temp_b5_12_28_r;
wire signed [`CalcTempBus]          temp_b5_12_28_i;
wire signed [`CalcTempBus]          temp_b5_12_29_r;
wire signed [`CalcTempBus]          temp_b5_12_29_i;
wire signed [`CalcTempBus]          temp_b5_12_30_r;
wire signed [`CalcTempBus]          temp_b5_12_30_i;
wire signed [`CalcTempBus]          temp_b5_12_31_r;
wire signed [`CalcTempBus]          temp_b5_12_31_i;
wire signed [`CalcTempBus]          temp_b5_12_32_r;
wire signed [`CalcTempBus]          temp_b5_12_32_i;
wire signed [`CalcTempBus]          temp_b5_13_1_r;
wire signed [`CalcTempBus]          temp_b5_13_1_i;
wire signed [`CalcTempBus]          temp_b5_13_2_r;
wire signed [`CalcTempBus]          temp_b5_13_2_i;
wire signed [`CalcTempBus]          temp_b5_13_3_r;
wire signed [`CalcTempBus]          temp_b5_13_3_i;
wire signed [`CalcTempBus]          temp_b5_13_4_r;
wire signed [`CalcTempBus]          temp_b5_13_4_i;
wire signed [`CalcTempBus]          temp_b5_13_5_r;
wire signed [`CalcTempBus]          temp_b5_13_5_i;
wire signed [`CalcTempBus]          temp_b5_13_6_r;
wire signed [`CalcTempBus]          temp_b5_13_6_i;
wire signed [`CalcTempBus]          temp_b5_13_7_r;
wire signed [`CalcTempBus]          temp_b5_13_7_i;
wire signed [`CalcTempBus]          temp_b5_13_8_r;
wire signed [`CalcTempBus]          temp_b5_13_8_i;
wire signed [`CalcTempBus]          temp_b5_13_9_r;
wire signed [`CalcTempBus]          temp_b5_13_9_i;
wire signed [`CalcTempBus]          temp_b5_13_10_r;
wire signed [`CalcTempBus]          temp_b5_13_10_i;
wire signed [`CalcTempBus]          temp_b5_13_11_r;
wire signed [`CalcTempBus]          temp_b5_13_11_i;
wire signed [`CalcTempBus]          temp_b5_13_12_r;
wire signed [`CalcTempBus]          temp_b5_13_12_i;
wire signed [`CalcTempBus]          temp_b5_13_13_r;
wire signed [`CalcTempBus]          temp_b5_13_13_i;
wire signed [`CalcTempBus]          temp_b5_13_14_r;
wire signed [`CalcTempBus]          temp_b5_13_14_i;
wire signed [`CalcTempBus]          temp_b5_13_15_r;
wire signed [`CalcTempBus]          temp_b5_13_15_i;
wire signed [`CalcTempBus]          temp_b5_13_16_r;
wire signed [`CalcTempBus]          temp_b5_13_16_i;
wire signed [`CalcTempBus]          temp_b5_13_17_r;
wire signed [`CalcTempBus]          temp_b5_13_17_i;
wire signed [`CalcTempBus]          temp_b5_13_18_r;
wire signed [`CalcTempBus]          temp_b5_13_18_i;
wire signed [`CalcTempBus]          temp_b5_13_19_r;
wire signed [`CalcTempBus]          temp_b5_13_19_i;
wire signed [`CalcTempBus]          temp_b5_13_20_r;
wire signed [`CalcTempBus]          temp_b5_13_20_i;
wire signed [`CalcTempBus]          temp_b5_13_21_r;
wire signed [`CalcTempBus]          temp_b5_13_21_i;
wire signed [`CalcTempBus]          temp_b5_13_22_r;
wire signed [`CalcTempBus]          temp_b5_13_22_i;
wire signed [`CalcTempBus]          temp_b5_13_23_r;
wire signed [`CalcTempBus]          temp_b5_13_23_i;
wire signed [`CalcTempBus]          temp_b5_13_24_r;
wire signed [`CalcTempBus]          temp_b5_13_24_i;
wire signed [`CalcTempBus]          temp_b5_13_25_r;
wire signed [`CalcTempBus]          temp_b5_13_25_i;
wire signed [`CalcTempBus]          temp_b5_13_26_r;
wire signed [`CalcTempBus]          temp_b5_13_26_i;
wire signed [`CalcTempBus]          temp_b5_13_27_r;
wire signed [`CalcTempBus]          temp_b5_13_27_i;
wire signed [`CalcTempBus]          temp_b5_13_28_r;
wire signed [`CalcTempBus]          temp_b5_13_28_i;
wire signed [`CalcTempBus]          temp_b5_13_29_r;
wire signed [`CalcTempBus]          temp_b5_13_29_i;
wire signed [`CalcTempBus]          temp_b5_13_30_r;
wire signed [`CalcTempBus]          temp_b5_13_30_i;
wire signed [`CalcTempBus]          temp_b5_13_31_r;
wire signed [`CalcTempBus]          temp_b5_13_31_i;
wire signed [`CalcTempBus]          temp_b5_13_32_r;
wire signed [`CalcTempBus]          temp_b5_13_32_i;
wire signed [`CalcTempBus]          temp_b5_14_1_r;
wire signed [`CalcTempBus]          temp_b5_14_1_i;
wire signed [`CalcTempBus]          temp_b5_14_2_r;
wire signed [`CalcTempBus]          temp_b5_14_2_i;
wire signed [`CalcTempBus]          temp_b5_14_3_r;
wire signed [`CalcTempBus]          temp_b5_14_3_i;
wire signed [`CalcTempBus]          temp_b5_14_4_r;
wire signed [`CalcTempBus]          temp_b5_14_4_i;
wire signed [`CalcTempBus]          temp_b5_14_5_r;
wire signed [`CalcTempBus]          temp_b5_14_5_i;
wire signed [`CalcTempBus]          temp_b5_14_6_r;
wire signed [`CalcTempBus]          temp_b5_14_6_i;
wire signed [`CalcTempBus]          temp_b5_14_7_r;
wire signed [`CalcTempBus]          temp_b5_14_7_i;
wire signed [`CalcTempBus]          temp_b5_14_8_r;
wire signed [`CalcTempBus]          temp_b5_14_8_i;
wire signed [`CalcTempBus]          temp_b5_14_9_r;
wire signed [`CalcTempBus]          temp_b5_14_9_i;
wire signed [`CalcTempBus]          temp_b5_14_10_r;
wire signed [`CalcTempBus]          temp_b5_14_10_i;
wire signed [`CalcTempBus]          temp_b5_14_11_r;
wire signed [`CalcTempBus]          temp_b5_14_11_i;
wire signed [`CalcTempBus]          temp_b5_14_12_r;
wire signed [`CalcTempBus]          temp_b5_14_12_i;
wire signed [`CalcTempBus]          temp_b5_14_13_r;
wire signed [`CalcTempBus]          temp_b5_14_13_i;
wire signed [`CalcTempBus]          temp_b5_14_14_r;
wire signed [`CalcTempBus]          temp_b5_14_14_i;
wire signed [`CalcTempBus]          temp_b5_14_15_r;
wire signed [`CalcTempBus]          temp_b5_14_15_i;
wire signed [`CalcTempBus]          temp_b5_14_16_r;
wire signed [`CalcTempBus]          temp_b5_14_16_i;
wire signed [`CalcTempBus]          temp_b5_14_17_r;
wire signed [`CalcTempBus]          temp_b5_14_17_i;
wire signed [`CalcTempBus]          temp_b5_14_18_r;
wire signed [`CalcTempBus]          temp_b5_14_18_i;
wire signed [`CalcTempBus]          temp_b5_14_19_r;
wire signed [`CalcTempBus]          temp_b5_14_19_i;
wire signed [`CalcTempBus]          temp_b5_14_20_r;
wire signed [`CalcTempBus]          temp_b5_14_20_i;
wire signed [`CalcTempBus]          temp_b5_14_21_r;
wire signed [`CalcTempBus]          temp_b5_14_21_i;
wire signed [`CalcTempBus]          temp_b5_14_22_r;
wire signed [`CalcTempBus]          temp_b5_14_22_i;
wire signed [`CalcTempBus]          temp_b5_14_23_r;
wire signed [`CalcTempBus]          temp_b5_14_23_i;
wire signed [`CalcTempBus]          temp_b5_14_24_r;
wire signed [`CalcTempBus]          temp_b5_14_24_i;
wire signed [`CalcTempBus]          temp_b5_14_25_r;
wire signed [`CalcTempBus]          temp_b5_14_25_i;
wire signed [`CalcTempBus]          temp_b5_14_26_r;
wire signed [`CalcTempBus]          temp_b5_14_26_i;
wire signed [`CalcTempBus]          temp_b5_14_27_r;
wire signed [`CalcTempBus]          temp_b5_14_27_i;
wire signed [`CalcTempBus]          temp_b5_14_28_r;
wire signed [`CalcTempBus]          temp_b5_14_28_i;
wire signed [`CalcTempBus]          temp_b5_14_29_r;
wire signed [`CalcTempBus]          temp_b5_14_29_i;
wire signed [`CalcTempBus]          temp_b5_14_30_r;
wire signed [`CalcTempBus]          temp_b5_14_30_i;
wire signed [`CalcTempBus]          temp_b5_14_31_r;
wire signed [`CalcTempBus]          temp_b5_14_31_i;
wire signed [`CalcTempBus]          temp_b5_14_32_r;
wire signed [`CalcTempBus]          temp_b5_14_32_i;
wire signed [`CalcTempBus]          temp_b5_15_1_r;
wire signed [`CalcTempBus]          temp_b5_15_1_i;
wire signed [`CalcTempBus]          temp_b5_15_2_r;
wire signed [`CalcTempBus]          temp_b5_15_2_i;
wire signed [`CalcTempBus]          temp_b5_15_3_r;
wire signed [`CalcTempBus]          temp_b5_15_3_i;
wire signed [`CalcTempBus]          temp_b5_15_4_r;
wire signed [`CalcTempBus]          temp_b5_15_4_i;
wire signed [`CalcTempBus]          temp_b5_15_5_r;
wire signed [`CalcTempBus]          temp_b5_15_5_i;
wire signed [`CalcTempBus]          temp_b5_15_6_r;
wire signed [`CalcTempBus]          temp_b5_15_6_i;
wire signed [`CalcTempBus]          temp_b5_15_7_r;
wire signed [`CalcTempBus]          temp_b5_15_7_i;
wire signed [`CalcTempBus]          temp_b5_15_8_r;
wire signed [`CalcTempBus]          temp_b5_15_8_i;
wire signed [`CalcTempBus]          temp_b5_15_9_r;
wire signed [`CalcTempBus]          temp_b5_15_9_i;
wire signed [`CalcTempBus]          temp_b5_15_10_r;
wire signed [`CalcTempBus]          temp_b5_15_10_i;
wire signed [`CalcTempBus]          temp_b5_15_11_r;
wire signed [`CalcTempBus]          temp_b5_15_11_i;
wire signed [`CalcTempBus]          temp_b5_15_12_r;
wire signed [`CalcTempBus]          temp_b5_15_12_i;
wire signed [`CalcTempBus]          temp_b5_15_13_r;
wire signed [`CalcTempBus]          temp_b5_15_13_i;
wire signed [`CalcTempBus]          temp_b5_15_14_r;
wire signed [`CalcTempBus]          temp_b5_15_14_i;
wire signed [`CalcTempBus]          temp_b5_15_15_r;
wire signed [`CalcTempBus]          temp_b5_15_15_i;
wire signed [`CalcTempBus]          temp_b5_15_16_r;
wire signed [`CalcTempBus]          temp_b5_15_16_i;
wire signed [`CalcTempBus]          temp_b5_15_17_r;
wire signed [`CalcTempBus]          temp_b5_15_17_i;
wire signed [`CalcTempBus]          temp_b5_15_18_r;
wire signed [`CalcTempBus]          temp_b5_15_18_i;
wire signed [`CalcTempBus]          temp_b5_15_19_r;
wire signed [`CalcTempBus]          temp_b5_15_19_i;
wire signed [`CalcTempBus]          temp_b5_15_20_r;
wire signed [`CalcTempBus]          temp_b5_15_20_i;
wire signed [`CalcTempBus]          temp_b5_15_21_r;
wire signed [`CalcTempBus]          temp_b5_15_21_i;
wire signed [`CalcTempBus]          temp_b5_15_22_r;
wire signed [`CalcTempBus]          temp_b5_15_22_i;
wire signed [`CalcTempBus]          temp_b5_15_23_r;
wire signed [`CalcTempBus]          temp_b5_15_23_i;
wire signed [`CalcTempBus]          temp_b5_15_24_r;
wire signed [`CalcTempBus]          temp_b5_15_24_i;
wire signed [`CalcTempBus]          temp_b5_15_25_r;
wire signed [`CalcTempBus]          temp_b5_15_25_i;
wire signed [`CalcTempBus]          temp_b5_15_26_r;
wire signed [`CalcTempBus]          temp_b5_15_26_i;
wire signed [`CalcTempBus]          temp_b5_15_27_r;
wire signed [`CalcTempBus]          temp_b5_15_27_i;
wire signed [`CalcTempBus]          temp_b5_15_28_r;
wire signed [`CalcTempBus]          temp_b5_15_28_i;
wire signed [`CalcTempBus]          temp_b5_15_29_r;
wire signed [`CalcTempBus]          temp_b5_15_29_i;
wire signed [`CalcTempBus]          temp_b5_15_30_r;
wire signed [`CalcTempBus]          temp_b5_15_30_i;
wire signed [`CalcTempBus]          temp_b5_15_31_r;
wire signed [`CalcTempBus]          temp_b5_15_31_i;
wire signed [`CalcTempBus]          temp_b5_15_32_r;
wire signed [`CalcTempBus]          temp_b5_15_32_i;
wire signed [`CalcTempBus]          temp_b5_16_1_r;
wire signed [`CalcTempBus]          temp_b5_16_1_i;
wire signed [`CalcTempBus]          temp_b5_16_2_r;
wire signed [`CalcTempBus]          temp_b5_16_2_i;
wire signed [`CalcTempBus]          temp_b5_16_3_r;
wire signed [`CalcTempBus]          temp_b5_16_3_i;
wire signed [`CalcTempBus]          temp_b5_16_4_r;
wire signed [`CalcTempBus]          temp_b5_16_4_i;
wire signed [`CalcTempBus]          temp_b5_16_5_r;
wire signed [`CalcTempBus]          temp_b5_16_5_i;
wire signed [`CalcTempBus]          temp_b5_16_6_r;
wire signed [`CalcTempBus]          temp_b5_16_6_i;
wire signed [`CalcTempBus]          temp_b5_16_7_r;
wire signed [`CalcTempBus]          temp_b5_16_7_i;
wire signed [`CalcTempBus]          temp_b5_16_8_r;
wire signed [`CalcTempBus]          temp_b5_16_8_i;
wire signed [`CalcTempBus]          temp_b5_16_9_r;
wire signed [`CalcTempBus]          temp_b5_16_9_i;
wire signed [`CalcTempBus]          temp_b5_16_10_r;
wire signed [`CalcTempBus]          temp_b5_16_10_i;
wire signed [`CalcTempBus]          temp_b5_16_11_r;
wire signed [`CalcTempBus]          temp_b5_16_11_i;
wire signed [`CalcTempBus]          temp_b5_16_12_r;
wire signed [`CalcTempBus]          temp_b5_16_12_i;
wire signed [`CalcTempBus]          temp_b5_16_13_r;
wire signed [`CalcTempBus]          temp_b5_16_13_i;
wire signed [`CalcTempBus]          temp_b5_16_14_r;
wire signed [`CalcTempBus]          temp_b5_16_14_i;
wire signed [`CalcTempBus]          temp_b5_16_15_r;
wire signed [`CalcTempBus]          temp_b5_16_15_i;
wire signed [`CalcTempBus]          temp_b5_16_16_r;
wire signed [`CalcTempBus]          temp_b5_16_16_i;
wire signed [`CalcTempBus]          temp_b5_16_17_r;
wire signed [`CalcTempBus]          temp_b5_16_17_i;
wire signed [`CalcTempBus]          temp_b5_16_18_r;
wire signed [`CalcTempBus]          temp_b5_16_18_i;
wire signed [`CalcTempBus]          temp_b5_16_19_r;
wire signed [`CalcTempBus]          temp_b5_16_19_i;
wire signed [`CalcTempBus]          temp_b5_16_20_r;
wire signed [`CalcTempBus]          temp_b5_16_20_i;
wire signed [`CalcTempBus]          temp_b5_16_21_r;
wire signed [`CalcTempBus]          temp_b5_16_21_i;
wire signed [`CalcTempBus]          temp_b5_16_22_r;
wire signed [`CalcTempBus]          temp_b5_16_22_i;
wire signed [`CalcTempBus]          temp_b5_16_23_r;
wire signed [`CalcTempBus]          temp_b5_16_23_i;
wire signed [`CalcTempBus]          temp_b5_16_24_r;
wire signed [`CalcTempBus]          temp_b5_16_24_i;
wire signed [`CalcTempBus]          temp_b5_16_25_r;
wire signed [`CalcTempBus]          temp_b5_16_25_i;
wire signed [`CalcTempBus]          temp_b5_16_26_r;
wire signed [`CalcTempBus]          temp_b5_16_26_i;
wire signed [`CalcTempBus]          temp_b5_16_27_r;
wire signed [`CalcTempBus]          temp_b5_16_27_i;
wire signed [`CalcTempBus]          temp_b5_16_28_r;
wire signed [`CalcTempBus]          temp_b5_16_28_i;
wire signed [`CalcTempBus]          temp_b5_16_29_r;
wire signed [`CalcTempBus]          temp_b5_16_29_i;
wire signed [`CalcTempBus]          temp_b5_16_30_r;
wire signed [`CalcTempBus]          temp_b5_16_30_i;
wire signed [`CalcTempBus]          temp_b5_16_31_r;
wire signed [`CalcTempBus]          temp_b5_16_31_i;
wire signed [`CalcTempBus]          temp_b5_16_32_r;
wire signed [`CalcTempBus]          temp_b5_16_32_i;
wire signed [`CalcTempBus]          temp_b5_17_1_r;
wire signed [`CalcTempBus]          temp_b5_17_1_i;
wire signed [`CalcTempBus]          temp_b5_17_2_r;
wire signed [`CalcTempBus]          temp_b5_17_2_i;
wire signed [`CalcTempBus]          temp_b5_17_3_r;
wire signed [`CalcTempBus]          temp_b5_17_3_i;
wire signed [`CalcTempBus]          temp_b5_17_4_r;
wire signed [`CalcTempBus]          temp_b5_17_4_i;
wire signed [`CalcTempBus]          temp_b5_17_5_r;
wire signed [`CalcTempBus]          temp_b5_17_5_i;
wire signed [`CalcTempBus]          temp_b5_17_6_r;
wire signed [`CalcTempBus]          temp_b5_17_6_i;
wire signed [`CalcTempBus]          temp_b5_17_7_r;
wire signed [`CalcTempBus]          temp_b5_17_7_i;
wire signed [`CalcTempBus]          temp_b5_17_8_r;
wire signed [`CalcTempBus]          temp_b5_17_8_i;
wire signed [`CalcTempBus]          temp_b5_17_9_r;
wire signed [`CalcTempBus]          temp_b5_17_9_i;
wire signed [`CalcTempBus]          temp_b5_17_10_r;
wire signed [`CalcTempBus]          temp_b5_17_10_i;
wire signed [`CalcTempBus]          temp_b5_17_11_r;
wire signed [`CalcTempBus]          temp_b5_17_11_i;
wire signed [`CalcTempBus]          temp_b5_17_12_r;
wire signed [`CalcTempBus]          temp_b5_17_12_i;
wire signed [`CalcTempBus]          temp_b5_17_13_r;
wire signed [`CalcTempBus]          temp_b5_17_13_i;
wire signed [`CalcTempBus]          temp_b5_17_14_r;
wire signed [`CalcTempBus]          temp_b5_17_14_i;
wire signed [`CalcTempBus]          temp_b5_17_15_r;
wire signed [`CalcTempBus]          temp_b5_17_15_i;
wire signed [`CalcTempBus]          temp_b5_17_16_r;
wire signed [`CalcTempBus]          temp_b5_17_16_i;
wire signed [`CalcTempBus]          temp_b5_17_17_r;
wire signed [`CalcTempBus]          temp_b5_17_17_i;
wire signed [`CalcTempBus]          temp_b5_17_18_r;
wire signed [`CalcTempBus]          temp_b5_17_18_i;
wire signed [`CalcTempBus]          temp_b5_17_19_r;
wire signed [`CalcTempBus]          temp_b5_17_19_i;
wire signed [`CalcTempBus]          temp_b5_17_20_r;
wire signed [`CalcTempBus]          temp_b5_17_20_i;
wire signed [`CalcTempBus]          temp_b5_17_21_r;
wire signed [`CalcTempBus]          temp_b5_17_21_i;
wire signed [`CalcTempBus]          temp_b5_17_22_r;
wire signed [`CalcTempBus]          temp_b5_17_22_i;
wire signed [`CalcTempBus]          temp_b5_17_23_r;
wire signed [`CalcTempBus]          temp_b5_17_23_i;
wire signed [`CalcTempBus]          temp_b5_17_24_r;
wire signed [`CalcTempBus]          temp_b5_17_24_i;
wire signed [`CalcTempBus]          temp_b5_17_25_r;
wire signed [`CalcTempBus]          temp_b5_17_25_i;
wire signed [`CalcTempBus]          temp_b5_17_26_r;
wire signed [`CalcTempBus]          temp_b5_17_26_i;
wire signed [`CalcTempBus]          temp_b5_17_27_r;
wire signed [`CalcTempBus]          temp_b5_17_27_i;
wire signed [`CalcTempBus]          temp_b5_17_28_r;
wire signed [`CalcTempBus]          temp_b5_17_28_i;
wire signed [`CalcTempBus]          temp_b5_17_29_r;
wire signed [`CalcTempBus]          temp_b5_17_29_i;
wire signed [`CalcTempBus]          temp_b5_17_30_r;
wire signed [`CalcTempBus]          temp_b5_17_30_i;
wire signed [`CalcTempBus]          temp_b5_17_31_r;
wire signed [`CalcTempBus]          temp_b5_17_31_i;
wire signed [`CalcTempBus]          temp_b5_17_32_r;
wire signed [`CalcTempBus]          temp_b5_17_32_i;
wire signed [`CalcTempBus]          temp_b5_18_1_r;
wire signed [`CalcTempBus]          temp_b5_18_1_i;
wire signed [`CalcTempBus]          temp_b5_18_2_r;
wire signed [`CalcTempBus]          temp_b5_18_2_i;
wire signed [`CalcTempBus]          temp_b5_18_3_r;
wire signed [`CalcTempBus]          temp_b5_18_3_i;
wire signed [`CalcTempBus]          temp_b5_18_4_r;
wire signed [`CalcTempBus]          temp_b5_18_4_i;
wire signed [`CalcTempBus]          temp_b5_18_5_r;
wire signed [`CalcTempBus]          temp_b5_18_5_i;
wire signed [`CalcTempBus]          temp_b5_18_6_r;
wire signed [`CalcTempBus]          temp_b5_18_6_i;
wire signed [`CalcTempBus]          temp_b5_18_7_r;
wire signed [`CalcTempBus]          temp_b5_18_7_i;
wire signed [`CalcTempBus]          temp_b5_18_8_r;
wire signed [`CalcTempBus]          temp_b5_18_8_i;
wire signed [`CalcTempBus]          temp_b5_18_9_r;
wire signed [`CalcTempBus]          temp_b5_18_9_i;
wire signed [`CalcTempBus]          temp_b5_18_10_r;
wire signed [`CalcTempBus]          temp_b5_18_10_i;
wire signed [`CalcTempBus]          temp_b5_18_11_r;
wire signed [`CalcTempBus]          temp_b5_18_11_i;
wire signed [`CalcTempBus]          temp_b5_18_12_r;
wire signed [`CalcTempBus]          temp_b5_18_12_i;
wire signed [`CalcTempBus]          temp_b5_18_13_r;
wire signed [`CalcTempBus]          temp_b5_18_13_i;
wire signed [`CalcTempBus]          temp_b5_18_14_r;
wire signed [`CalcTempBus]          temp_b5_18_14_i;
wire signed [`CalcTempBus]          temp_b5_18_15_r;
wire signed [`CalcTempBus]          temp_b5_18_15_i;
wire signed [`CalcTempBus]          temp_b5_18_16_r;
wire signed [`CalcTempBus]          temp_b5_18_16_i;
wire signed [`CalcTempBus]          temp_b5_18_17_r;
wire signed [`CalcTempBus]          temp_b5_18_17_i;
wire signed [`CalcTempBus]          temp_b5_18_18_r;
wire signed [`CalcTempBus]          temp_b5_18_18_i;
wire signed [`CalcTempBus]          temp_b5_18_19_r;
wire signed [`CalcTempBus]          temp_b5_18_19_i;
wire signed [`CalcTempBus]          temp_b5_18_20_r;
wire signed [`CalcTempBus]          temp_b5_18_20_i;
wire signed [`CalcTempBus]          temp_b5_18_21_r;
wire signed [`CalcTempBus]          temp_b5_18_21_i;
wire signed [`CalcTempBus]          temp_b5_18_22_r;
wire signed [`CalcTempBus]          temp_b5_18_22_i;
wire signed [`CalcTempBus]          temp_b5_18_23_r;
wire signed [`CalcTempBus]          temp_b5_18_23_i;
wire signed [`CalcTempBus]          temp_b5_18_24_r;
wire signed [`CalcTempBus]          temp_b5_18_24_i;
wire signed [`CalcTempBus]          temp_b5_18_25_r;
wire signed [`CalcTempBus]          temp_b5_18_25_i;
wire signed [`CalcTempBus]          temp_b5_18_26_r;
wire signed [`CalcTempBus]          temp_b5_18_26_i;
wire signed [`CalcTempBus]          temp_b5_18_27_r;
wire signed [`CalcTempBus]          temp_b5_18_27_i;
wire signed [`CalcTempBus]          temp_b5_18_28_r;
wire signed [`CalcTempBus]          temp_b5_18_28_i;
wire signed [`CalcTempBus]          temp_b5_18_29_r;
wire signed [`CalcTempBus]          temp_b5_18_29_i;
wire signed [`CalcTempBus]          temp_b5_18_30_r;
wire signed [`CalcTempBus]          temp_b5_18_30_i;
wire signed [`CalcTempBus]          temp_b5_18_31_r;
wire signed [`CalcTempBus]          temp_b5_18_31_i;
wire signed [`CalcTempBus]          temp_b5_18_32_r;
wire signed [`CalcTempBus]          temp_b5_18_32_i;
wire signed [`CalcTempBus]          temp_b5_19_1_r;
wire signed [`CalcTempBus]          temp_b5_19_1_i;
wire signed [`CalcTempBus]          temp_b5_19_2_r;
wire signed [`CalcTempBus]          temp_b5_19_2_i;
wire signed [`CalcTempBus]          temp_b5_19_3_r;
wire signed [`CalcTempBus]          temp_b5_19_3_i;
wire signed [`CalcTempBus]          temp_b5_19_4_r;
wire signed [`CalcTempBus]          temp_b5_19_4_i;
wire signed [`CalcTempBus]          temp_b5_19_5_r;
wire signed [`CalcTempBus]          temp_b5_19_5_i;
wire signed [`CalcTempBus]          temp_b5_19_6_r;
wire signed [`CalcTempBus]          temp_b5_19_6_i;
wire signed [`CalcTempBus]          temp_b5_19_7_r;
wire signed [`CalcTempBus]          temp_b5_19_7_i;
wire signed [`CalcTempBus]          temp_b5_19_8_r;
wire signed [`CalcTempBus]          temp_b5_19_8_i;
wire signed [`CalcTempBus]          temp_b5_19_9_r;
wire signed [`CalcTempBus]          temp_b5_19_9_i;
wire signed [`CalcTempBus]          temp_b5_19_10_r;
wire signed [`CalcTempBus]          temp_b5_19_10_i;
wire signed [`CalcTempBus]          temp_b5_19_11_r;
wire signed [`CalcTempBus]          temp_b5_19_11_i;
wire signed [`CalcTempBus]          temp_b5_19_12_r;
wire signed [`CalcTempBus]          temp_b5_19_12_i;
wire signed [`CalcTempBus]          temp_b5_19_13_r;
wire signed [`CalcTempBus]          temp_b5_19_13_i;
wire signed [`CalcTempBus]          temp_b5_19_14_r;
wire signed [`CalcTempBus]          temp_b5_19_14_i;
wire signed [`CalcTempBus]          temp_b5_19_15_r;
wire signed [`CalcTempBus]          temp_b5_19_15_i;
wire signed [`CalcTempBus]          temp_b5_19_16_r;
wire signed [`CalcTempBus]          temp_b5_19_16_i;
wire signed [`CalcTempBus]          temp_b5_19_17_r;
wire signed [`CalcTempBus]          temp_b5_19_17_i;
wire signed [`CalcTempBus]          temp_b5_19_18_r;
wire signed [`CalcTempBus]          temp_b5_19_18_i;
wire signed [`CalcTempBus]          temp_b5_19_19_r;
wire signed [`CalcTempBus]          temp_b5_19_19_i;
wire signed [`CalcTempBus]          temp_b5_19_20_r;
wire signed [`CalcTempBus]          temp_b5_19_20_i;
wire signed [`CalcTempBus]          temp_b5_19_21_r;
wire signed [`CalcTempBus]          temp_b5_19_21_i;
wire signed [`CalcTempBus]          temp_b5_19_22_r;
wire signed [`CalcTempBus]          temp_b5_19_22_i;
wire signed [`CalcTempBus]          temp_b5_19_23_r;
wire signed [`CalcTempBus]          temp_b5_19_23_i;
wire signed [`CalcTempBus]          temp_b5_19_24_r;
wire signed [`CalcTempBus]          temp_b5_19_24_i;
wire signed [`CalcTempBus]          temp_b5_19_25_r;
wire signed [`CalcTempBus]          temp_b5_19_25_i;
wire signed [`CalcTempBus]          temp_b5_19_26_r;
wire signed [`CalcTempBus]          temp_b5_19_26_i;
wire signed [`CalcTempBus]          temp_b5_19_27_r;
wire signed [`CalcTempBus]          temp_b5_19_27_i;
wire signed [`CalcTempBus]          temp_b5_19_28_r;
wire signed [`CalcTempBus]          temp_b5_19_28_i;
wire signed [`CalcTempBus]          temp_b5_19_29_r;
wire signed [`CalcTempBus]          temp_b5_19_29_i;
wire signed [`CalcTempBus]          temp_b5_19_30_r;
wire signed [`CalcTempBus]          temp_b5_19_30_i;
wire signed [`CalcTempBus]          temp_b5_19_31_r;
wire signed [`CalcTempBus]          temp_b5_19_31_i;
wire signed [`CalcTempBus]          temp_b5_19_32_r;
wire signed [`CalcTempBus]          temp_b5_19_32_i;
wire signed [`CalcTempBus]          temp_b5_20_1_r;
wire signed [`CalcTempBus]          temp_b5_20_1_i;
wire signed [`CalcTempBus]          temp_b5_20_2_r;
wire signed [`CalcTempBus]          temp_b5_20_2_i;
wire signed [`CalcTempBus]          temp_b5_20_3_r;
wire signed [`CalcTempBus]          temp_b5_20_3_i;
wire signed [`CalcTempBus]          temp_b5_20_4_r;
wire signed [`CalcTempBus]          temp_b5_20_4_i;
wire signed [`CalcTempBus]          temp_b5_20_5_r;
wire signed [`CalcTempBus]          temp_b5_20_5_i;
wire signed [`CalcTempBus]          temp_b5_20_6_r;
wire signed [`CalcTempBus]          temp_b5_20_6_i;
wire signed [`CalcTempBus]          temp_b5_20_7_r;
wire signed [`CalcTempBus]          temp_b5_20_7_i;
wire signed [`CalcTempBus]          temp_b5_20_8_r;
wire signed [`CalcTempBus]          temp_b5_20_8_i;
wire signed [`CalcTempBus]          temp_b5_20_9_r;
wire signed [`CalcTempBus]          temp_b5_20_9_i;
wire signed [`CalcTempBus]          temp_b5_20_10_r;
wire signed [`CalcTempBus]          temp_b5_20_10_i;
wire signed [`CalcTempBus]          temp_b5_20_11_r;
wire signed [`CalcTempBus]          temp_b5_20_11_i;
wire signed [`CalcTempBus]          temp_b5_20_12_r;
wire signed [`CalcTempBus]          temp_b5_20_12_i;
wire signed [`CalcTempBus]          temp_b5_20_13_r;
wire signed [`CalcTempBus]          temp_b5_20_13_i;
wire signed [`CalcTempBus]          temp_b5_20_14_r;
wire signed [`CalcTempBus]          temp_b5_20_14_i;
wire signed [`CalcTempBus]          temp_b5_20_15_r;
wire signed [`CalcTempBus]          temp_b5_20_15_i;
wire signed [`CalcTempBus]          temp_b5_20_16_r;
wire signed [`CalcTempBus]          temp_b5_20_16_i;
wire signed [`CalcTempBus]          temp_b5_20_17_r;
wire signed [`CalcTempBus]          temp_b5_20_17_i;
wire signed [`CalcTempBus]          temp_b5_20_18_r;
wire signed [`CalcTempBus]          temp_b5_20_18_i;
wire signed [`CalcTempBus]          temp_b5_20_19_r;
wire signed [`CalcTempBus]          temp_b5_20_19_i;
wire signed [`CalcTempBus]          temp_b5_20_20_r;
wire signed [`CalcTempBus]          temp_b5_20_20_i;
wire signed [`CalcTempBus]          temp_b5_20_21_r;
wire signed [`CalcTempBus]          temp_b5_20_21_i;
wire signed [`CalcTempBus]          temp_b5_20_22_r;
wire signed [`CalcTempBus]          temp_b5_20_22_i;
wire signed [`CalcTempBus]          temp_b5_20_23_r;
wire signed [`CalcTempBus]          temp_b5_20_23_i;
wire signed [`CalcTempBus]          temp_b5_20_24_r;
wire signed [`CalcTempBus]          temp_b5_20_24_i;
wire signed [`CalcTempBus]          temp_b5_20_25_r;
wire signed [`CalcTempBus]          temp_b5_20_25_i;
wire signed [`CalcTempBus]          temp_b5_20_26_r;
wire signed [`CalcTempBus]          temp_b5_20_26_i;
wire signed [`CalcTempBus]          temp_b5_20_27_r;
wire signed [`CalcTempBus]          temp_b5_20_27_i;
wire signed [`CalcTempBus]          temp_b5_20_28_r;
wire signed [`CalcTempBus]          temp_b5_20_28_i;
wire signed [`CalcTempBus]          temp_b5_20_29_r;
wire signed [`CalcTempBus]          temp_b5_20_29_i;
wire signed [`CalcTempBus]          temp_b5_20_30_r;
wire signed [`CalcTempBus]          temp_b5_20_30_i;
wire signed [`CalcTempBus]          temp_b5_20_31_r;
wire signed [`CalcTempBus]          temp_b5_20_31_i;
wire signed [`CalcTempBus]          temp_b5_20_32_r;
wire signed [`CalcTempBus]          temp_b5_20_32_i;
wire signed [`CalcTempBus]          temp_b5_21_1_r;
wire signed [`CalcTempBus]          temp_b5_21_1_i;
wire signed [`CalcTempBus]          temp_b5_21_2_r;
wire signed [`CalcTempBus]          temp_b5_21_2_i;
wire signed [`CalcTempBus]          temp_b5_21_3_r;
wire signed [`CalcTempBus]          temp_b5_21_3_i;
wire signed [`CalcTempBus]          temp_b5_21_4_r;
wire signed [`CalcTempBus]          temp_b5_21_4_i;
wire signed [`CalcTempBus]          temp_b5_21_5_r;
wire signed [`CalcTempBus]          temp_b5_21_5_i;
wire signed [`CalcTempBus]          temp_b5_21_6_r;
wire signed [`CalcTempBus]          temp_b5_21_6_i;
wire signed [`CalcTempBus]          temp_b5_21_7_r;
wire signed [`CalcTempBus]          temp_b5_21_7_i;
wire signed [`CalcTempBus]          temp_b5_21_8_r;
wire signed [`CalcTempBus]          temp_b5_21_8_i;
wire signed [`CalcTempBus]          temp_b5_21_9_r;
wire signed [`CalcTempBus]          temp_b5_21_9_i;
wire signed [`CalcTempBus]          temp_b5_21_10_r;
wire signed [`CalcTempBus]          temp_b5_21_10_i;
wire signed [`CalcTempBus]          temp_b5_21_11_r;
wire signed [`CalcTempBus]          temp_b5_21_11_i;
wire signed [`CalcTempBus]          temp_b5_21_12_r;
wire signed [`CalcTempBus]          temp_b5_21_12_i;
wire signed [`CalcTempBus]          temp_b5_21_13_r;
wire signed [`CalcTempBus]          temp_b5_21_13_i;
wire signed [`CalcTempBus]          temp_b5_21_14_r;
wire signed [`CalcTempBus]          temp_b5_21_14_i;
wire signed [`CalcTempBus]          temp_b5_21_15_r;
wire signed [`CalcTempBus]          temp_b5_21_15_i;
wire signed [`CalcTempBus]          temp_b5_21_16_r;
wire signed [`CalcTempBus]          temp_b5_21_16_i;
wire signed [`CalcTempBus]          temp_b5_21_17_r;
wire signed [`CalcTempBus]          temp_b5_21_17_i;
wire signed [`CalcTempBus]          temp_b5_21_18_r;
wire signed [`CalcTempBus]          temp_b5_21_18_i;
wire signed [`CalcTempBus]          temp_b5_21_19_r;
wire signed [`CalcTempBus]          temp_b5_21_19_i;
wire signed [`CalcTempBus]          temp_b5_21_20_r;
wire signed [`CalcTempBus]          temp_b5_21_20_i;
wire signed [`CalcTempBus]          temp_b5_21_21_r;
wire signed [`CalcTempBus]          temp_b5_21_21_i;
wire signed [`CalcTempBus]          temp_b5_21_22_r;
wire signed [`CalcTempBus]          temp_b5_21_22_i;
wire signed [`CalcTempBus]          temp_b5_21_23_r;
wire signed [`CalcTempBus]          temp_b5_21_23_i;
wire signed [`CalcTempBus]          temp_b5_21_24_r;
wire signed [`CalcTempBus]          temp_b5_21_24_i;
wire signed [`CalcTempBus]          temp_b5_21_25_r;
wire signed [`CalcTempBus]          temp_b5_21_25_i;
wire signed [`CalcTempBus]          temp_b5_21_26_r;
wire signed [`CalcTempBus]          temp_b5_21_26_i;
wire signed [`CalcTempBus]          temp_b5_21_27_r;
wire signed [`CalcTempBus]          temp_b5_21_27_i;
wire signed [`CalcTempBus]          temp_b5_21_28_r;
wire signed [`CalcTempBus]          temp_b5_21_28_i;
wire signed [`CalcTempBus]          temp_b5_21_29_r;
wire signed [`CalcTempBus]          temp_b5_21_29_i;
wire signed [`CalcTempBus]          temp_b5_21_30_r;
wire signed [`CalcTempBus]          temp_b5_21_30_i;
wire signed [`CalcTempBus]          temp_b5_21_31_r;
wire signed [`CalcTempBus]          temp_b5_21_31_i;
wire signed [`CalcTempBus]          temp_b5_21_32_r;
wire signed [`CalcTempBus]          temp_b5_21_32_i;
wire signed [`CalcTempBus]          temp_b5_22_1_r;
wire signed [`CalcTempBus]          temp_b5_22_1_i;
wire signed [`CalcTempBus]          temp_b5_22_2_r;
wire signed [`CalcTempBus]          temp_b5_22_2_i;
wire signed [`CalcTempBus]          temp_b5_22_3_r;
wire signed [`CalcTempBus]          temp_b5_22_3_i;
wire signed [`CalcTempBus]          temp_b5_22_4_r;
wire signed [`CalcTempBus]          temp_b5_22_4_i;
wire signed [`CalcTempBus]          temp_b5_22_5_r;
wire signed [`CalcTempBus]          temp_b5_22_5_i;
wire signed [`CalcTempBus]          temp_b5_22_6_r;
wire signed [`CalcTempBus]          temp_b5_22_6_i;
wire signed [`CalcTempBus]          temp_b5_22_7_r;
wire signed [`CalcTempBus]          temp_b5_22_7_i;
wire signed [`CalcTempBus]          temp_b5_22_8_r;
wire signed [`CalcTempBus]          temp_b5_22_8_i;
wire signed [`CalcTempBus]          temp_b5_22_9_r;
wire signed [`CalcTempBus]          temp_b5_22_9_i;
wire signed [`CalcTempBus]          temp_b5_22_10_r;
wire signed [`CalcTempBus]          temp_b5_22_10_i;
wire signed [`CalcTempBus]          temp_b5_22_11_r;
wire signed [`CalcTempBus]          temp_b5_22_11_i;
wire signed [`CalcTempBus]          temp_b5_22_12_r;
wire signed [`CalcTempBus]          temp_b5_22_12_i;
wire signed [`CalcTempBus]          temp_b5_22_13_r;
wire signed [`CalcTempBus]          temp_b5_22_13_i;
wire signed [`CalcTempBus]          temp_b5_22_14_r;
wire signed [`CalcTempBus]          temp_b5_22_14_i;
wire signed [`CalcTempBus]          temp_b5_22_15_r;
wire signed [`CalcTempBus]          temp_b5_22_15_i;
wire signed [`CalcTempBus]          temp_b5_22_16_r;
wire signed [`CalcTempBus]          temp_b5_22_16_i;
wire signed [`CalcTempBus]          temp_b5_22_17_r;
wire signed [`CalcTempBus]          temp_b5_22_17_i;
wire signed [`CalcTempBus]          temp_b5_22_18_r;
wire signed [`CalcTempBus]          temp_b5_22_18_i;
wire signed [`CalcTempBus]          temp_b5_22_19_r;
wire signed [`CalcTempBus]          temp_b5_22_19_i;
wire signed [`CalcTempBus]          temp_b5_22_20_r;
wire signed [`CalcTempBus]          temp_b5_22_20_i;
wire signed [`CalcTempBus]          temp_b5_22_21_r;
wire signed [`CalcTempBus]          temp_b5_22_21_i;
wire signed [`CalcTempBus]          temp_b5_22_22_r;
wire signed [`CalcTempBus]          temp_b5_22_22_i;
wire signed [`CalcTempBus]          temp_b5_22_23_r;
wire signed [`CalcTempBus]          temp_b5_22_23_i;
wire signed [`CalcTempBus]          temp_b5_22_24_r;
wire signed [`CalcTempBus]          temp_b5_22_24_i;
wire signed [`CalcTempBus]          temp_b5_22_25_r;
wire signed [`CalcTempBus]          temp_b5_22_25_i;
wire signed [`CalcTempBus]          temp_b5_22_26_r;
wire signed [`CalcTempBus]          temp_b5_22_26_i;
wire signed [`CalcTempBus]          temp_b5_22_27_r;
wire signed [`CalcTempBus]          temp_b5_22_27_i;
wire signed [`CalcTempBus]          temp_b5_22_28_r;
wire signed [`CalcTempBus]          temp_b5_22_28_i;
wire signed [`CalcTempBus]          temp_b5_22_29_r;
wire signed [`CalcTempBus]          temp_b5_22_29_i;
wire signed [`CalcTempBus]          temp_b5_22_30_r;
wire signed [`CalcTempBus]          temp_b5_22_30_i;
wire signed [`CalcTempBus]          temp_b5_22_31_r;
wire signed [`CalcTempBus]          temp_b5_22_31_i;
wire signed [`CalcTempBus]          temp_b5_22_32_r;
wire signed [`CalcTempBus]          temp_b5_22_32_i;
wire signed [`CalcTempBus]          temp_b5_23_1_r;
wire signed [`CalcTempBus]          temp_b5_23_1_i;
wire signed [`CalcTempBus]          temp_b5_23_2_r;
wire signed [`CalcTempBus]          temp_b5_23_2_i;
wire signed [`CalcTempBus]          temp_b5_23_3_r;
wire signed [`CalcTempBus]          temp_b5_23_3_i;
wire signed [`CalcTempBus]          temp_b5_23_4_r;
wire signed [`CalcTempBus]          temp_b5_23_4_i;
wire signed [`CalcTempBus]          temp_b5_23_5_r;
wire signed [`CalcTempBus]          temp_b5_23_5_i;
wire signed [`CalcTempBus]          temp_b5_23_6_r;
wire signed [`CalcTempBus]          temp_b5_23_6_i;
wire signed [`CalcTempBus]          temp_b5_23_7_r;
wire signed [`CalcTempBus]          temp_b5_23_7_i;
wire signed [`CalcTempBus]          temp_b5_23_8_r;
wire signed [`CalcTempBus]          temp_b5_23_8_i;
wire signed [`CalcTempBus]          temp_b5_23_9_r;
wire signed [`CalcTempBus]          temp_b5_23_9_i;
wire signed [`CalcTempBus]          temp_b5_23_10_r;
wire signed [`CalcTempBus]          temp_b5_23_10_i;
wire signed [`CalcTempBus]          temp_b5_23_11_r;
wire signed [`CalcTempBus]          temp_b5_23_11_i;
wire signed [`CalcTempBus]          temp_b5_23_12_r;
wire signed [`CalcTempBus]          temp_b5_23_12_i;
wire signed [`CalcTempBus]          temp_b5_23_13_r;
wire signed [`CalcTempBus]          temp_b5_23_13_i;
wire signed [`CalcTempBus]          temp_b5_23_14_r;
wire signed [`CalcTempBus]          temp_b5_23_14_i;
wire signed [`CalcTempBus]          temp_b5_23_15_r;
wire signed [`CalcTempBus]          temp_b5_23_15_i;
wire signed [`CalcTempBus]          temp_b5_23_16_r;
wire signed [`CalcTempBus]          temp_b5_23_16_i;
wire signed [`CalcTempBus]          temp_b5_23_17_r;
wire signed [`CalcTempBus]          temp_b5_23_17_i;
wire signed [`CalcTempBus]          temp_b5_23_18_r;
wire signed [`CalcTempBus]          temp_b5_23_18_i;
wire signed [`CalcTempBus]          temp_b5_23_19_r;
wire signed [`CalcTempBus]          temp_b5_23_19_i;
wire signed [`CalcTempBus]          temp_b5_23_20_r;
wire signed [`CalcTempBus]          temp_b5_23_20_i;
wire signed [`CalcTempBus]          temp_b5_23_21_r;
wire signed [`CalcTempBus]          temp_b5_23_21_i;
wire signed [`CalcTempBus]          temp_b5_23_22_r;
wire signed [`CalcTempBus]          temp_b5_23_22_i;
wire signed [`CalcTempBus]          temp_b5_23_23_r;
wire signed [`CalcTempBus]          temp_b5_23_23_i;
wire signed [`CalcTempBus]          temp_b5_23_24_r;
wire signed [`CalcTempBus]          temp_b5_23_24_i;
wire signed [`CalcTempBus]          temp_b5_23_25_r;
wire signed [`CalcTempBus]          temp_b5_23_25_i;
wire signed [`CalcTempBus]          temp_b5_23_26_r;
wire signed [`CalcTempBus]          temp_b5_23_26_i;
wire signed [`CalcTempBus]          temp_b5_23_27_r;
wire signed [`CalcTempBus]          temp_b5_23_27_i;
wire signed [`CalcTempBus]          temp_b5_23_28_r;
wire signed [`CalcTempBus]          temp_b5_23_28_i;
wire signed [`CalcTempBus]          temp_b5_23_29_r;
wire signed [`CalcTempBus]          temp_b5_23_29_i;
wire signed [`CalcTempBus]          temp_b5_23_30_r;
wire signed [`CalcTempBus]          temp_b5_23_30_i;
wire signed [`CalcTempBus]          temp_b5_23_31_r;
wire signed [`CalcTempBus]          temp_b5_23_31_i;
wire signed [`CalcTempBus]          temp_b5_23_32_r;
wire signed [`CalcTempBus]          temp_b5_23_32_i;
wire signed [`CalcTempBus]          temp_b5_24_1_r;
wire signed [`CalcTempBus]          temp_b5_24_1_i;
wire signed [`CalcTempBus]          temp_b5_24_2_r;
wire signed [`CalcTempBus]          temp_b5_24_2_i;
wire signed [`CalcTempBus]          temp_b5_24_3_r;
wire signed [`CalcTempBus]          temp_b5_24_3_i;
wire signed [`CalcTempBus]          temp_b5_24_4_r;
wire signed [`CalcTempBus]          temp_b5_24_4_i;
wire signed [`CalcTempBus]          temp_b5_24_5_r;
wire signed [`CalcTempBus]          temp_b5_24_5_i;
wire signed [`CalcTempBus]          temp_b5_24_6_r;
wire signed [`CalcTempBus]          temp_b5_24_6_i;
wire signed [`CalcTempBus]          temp_b5_24_7_r;
wire signed [`CalcTempBus]          temp_b5_24_7_i;
wire signed [`CalcTempBus]          temp_b5_24_8_r;
wire signed [`CalcTempBus]          temp_b5_24_8_i;
wire signed [`CalcTempBus]          temp_b5_24_9_r;
wire signed [`CalcTempBus]          temp_b5_24_9_i;
wire signed [`CalcTempBus]          temp_b5_24_10_r;
wire signed [`CalcTempBus]          temp_b5_24_10_i;
wire signed [`CalcTempBus]          temp_b5_24_11_r;
wire signed [`CalcTempBus]          temp_b5_24_11_i;
wire signed [`CalcTempBus]          temp_b5_24_12_r;
wire signed [`CalcTempBus]          temp_b5_24_12_i;
wire signed [`CalcTempBus]          temp_b5_24_13_r;
wire signed [`CalcTempBus]          temp_b5_24_13_i;
wire signed [`CalcTempBus]          temp_b5_24_14_r;
wire signed [`CalcTempBus]          temp_b5_24_14_i;
wire signed [`CalcTempBus]          temp_b5_24_15_r;
wire signed [`CalcTempBus]          temp_b5_24_15_i;
wire signed [`CalcTempBus]          temp_b5_24_16_r;
wire signed [`CalcTempBus]          temp_b5_24_16_i;
wire signed [`CalcTempBus]          temp_b5_24_17_r;
wire signed [`CalcTempBus]          temp_b5_24_17_i;
wire signed [`CalcTempBus]          temp_b5_24_18_r;
wire signed [`CalcTempBus]          temp_b5_24_18_i;
wire signed [`CalcTempBus]          temp_b5_24_19_r;
wire signed [`CalcTempBus]          temp_b5_24_19_i;
wire signed [`CalcTempBus]          temp_b5_24_20_r;
wire signed [`CalcTempBus]          temp_b5_24_20_i;
wire signed [`CalcTempBus]          temp_b5_24_21_r;
wire signed [`CalcTempBus]          temp_b5_24_21_i;
wire signed [`CalcTempBus]          temp_b5_24_22_r;
wire signed [`CalcTempBus]          temp_b5_24_22_i;
wire signed [`CalcTempBus]          temp_b5_24_23_r;
wire signed [`CalcTempBus]          temp_b5_24_23_i;
wire signed [`CalcTempBus]          temp_b5_24_24_r;
wire signed [`CalcTempBus]          temp_b5_24_24_i;
wire signed [`CalcTempBus]          temp_b5_24_25_r;
wire signed [`CalcTempBus]          temp_b5_24_25_i;
wire signed [`CalcTempBus]          temp_b5_24_26_r;
wire signed [`CalcTempBus]          temp_b5_24_26_i;
wire signed [`CalcTempBus]          temp_b5_24_27_r;
wire signed [`CalcTempBus]          temp_b5_24_27_i;
wire signed [`CalcTempBus]          temp_b5_24_28_r;
wire signed [`CalcTempBus]          temp_b5_24_28_i;
wire signed [`CalcTempBus]          temp_b5_24_29_r;
wire signed [`CalcTempBus]          temp_b5_24_29_i;
wire signed [`CalcTempBus]          temp_b5_24_30_r;
wire signed [`CalcTempBus]          temp_b5_24_30_i;
wire signed [`CalcTempBus]          temp_b5_24_31_r;
wire signed [`CalcTempBus]          temp_b5_24_31_i;
wire signed [`CalcTempBus]          temp_b5_24_32_r;
wire signed [`CalcTempBus]          temp_b5_24_32_i;
wire signed [`CalcTempBus]          temp_b5_25_1_r;
wire signed [`CalcTempBus]          temp_b5_25_1_i;
wire signed [`CalcTempBus]          temp_b5_25_2_r;
wire signed [`CalcTempBus]          temp_b5_25_2_i;
wire signed [`CalcTempBus]          temp_b5_25_3_r;
wire signed [`CalcTempBus]          temp_b5_25_3_i;
wire signed [`CalcTempBus]          temp_b5_25_4_r;
wire signed [`CalcTempBus]          temp_b5_25_4_i;
wire signed [`CalcTempBus]          temp_b5_25_5_r;
wire signed [`CalcTempBus]          temp_b5_25_5_i;
wire signed [`CalcTempBus]          temp_b5_25_6_r;
wire signed [`CalcTempBus]          temp_b5_25_6_i;
wire signed [`CalcTempBus]          temp_b5_25_7_r;
wire signed [`CalcTempBus]          temp_b5_25_7_i;
wire signed [`CalcTempBus]          temp_b5_25_8_r;
wire signed [`CalcTempBus]          temp_b5_25_8_i;
wire signed [`CalcTempBus]          temp_b5_25_9_r;
wire signed [`CalcTempBus]          temp_b5_25_9_i;
wire signed [`CalcTempBus]          temp_b5_25_10_r;
wire signed [`CalcTempBus]          temp_b5_25_10_i;
wire signed [`CalcTempBus]          temp_b5_25_11_r;
wire signed [`CalcTempBus]          temp_b5_25_11_i;
wire signed [`CalcTempBus]          temp_b5_25_12_r;
wire signed [`CalcTempBus]          temp_b5_25_12_i;
wire signed [`CalcTempBus]          temp_b5_25_13_r;
wire signed [`CalcTempBus]          temp_b5_25_13_i;
wire signed [`CalcTempBus]          temp_b5_25_14_r;
wire signed [`CalcTempBus]          temp_b5_25_14_i;
wire signed [`CalcTempBus]          temp_b5_25_15_r;
wire signed [`CalcTempBus]          temp_b5_25_15_i;
wire signed [`CalcTempBus]          temp_b5_25_16_r;
wire signed [`CalcTempBus]          temp_b5_25_16_i;
wire signed [`CalcTempBus]          temp_b5_25_17_r;
wire signed [`CalcTempBus]          temp_b5_25_17_i;
wire signed [`CalcTempBus]          temp_b5_25_18_r;
wire signed [`CalcTempBus]          temp_b5_25_18_i;
wire signed [`CalcTempBus]          temp_b5_25_19_r;
wire signed [`CalcTempBus]          temp_b5_25_19_i;
wire signed [`CalcTempBus]          temp_b5_25_20_r;
wire signed [`CalcTempBus]          temp_b5_25_20_i;
wire signed [`CalcTempBus]          temp_b5_25_21_r;
wire signed [`CalcTempBus]          temp_b5_25_21_i;
wire signed [`CalcTempBus]          temp_b5_25_22_r;
wire signed [`CalcTempBus]          temp_b5_25_22_i;
wire signed [`CalcTempBus]          temp_b5_25_23_r;
wire signed [`CalcTempBus]          temp_b5_25_23_i;
wire signed [`CalcTempBus]          temp_b5_25_24_r;
wire signed [`CalcTempBus]          temp_b5_25_24_i;
wire signed [`CalcTempBus]          temp_b5_25_25_r;
wire signed [`CalcTempBus]          temp_b5_25_25_i;
wire signed [`CalcTempBus]          temp_b5_25_26_r;
wire signed [`CalcTempBus]          temp_b5_25_26_i;
wire signed [`CalcTempBus]          temp_b5_25_27_r;
wire signed [`CalcTempBus]          temp_b5_25_27_i;
wire signed [`CalcTempBus]          temp_b5_25_28_r;
wire signed [`CalcTempBus]          temp_b5_25_28_i;
wire signed [`CalcTempBus]          temp_b5_25_29_r;
wire signed [`CalcTempBus]          temp_b5_25_29_i;
wire signed [`CalcTempBus]          temp_b5_25_30_r;
wire signed [`CalcTempBus]          temp_b5_25_30_i;
wire signed [`CalcTempBus]          temp_b5_25_31_r;
wire signed [`CalcTempBus]          temp_b5_25_31_i;
wire signed [`CalcTempBus]          temp_b5_25_32_r;
wire signed [`CalcTempBus]          temp_b5_25_32_i;
wire signed [`CalcTempBus]          temp_b5_26_1_r;
wire signed [`CalcTempBus]          temp_b5_26_1_i;
wire signed [`CalcTempBus]          temp_b5_26_2_r;
wire signed [`CalcTempBus]          temp_b5_26_2_i;
wire signed [`CalcTempBus]          temp_b5_26_3_r;
wire signed [`CalcTempBus]          temp_b5_26_3_i;
wire signed [`CalcTempBus]          temp_b5_26_4_r;
wire signed [`CalcTempBus]          temp_b5_26_4_i;
wire signed [`CalcTempBus]          temp_b5_26_5_r;
wire signed [`CalcTempBus]          temp_b5_26_5_i;
wire signed [`CalcTempBus]          temp_b5_26_6_r;
wire signed [`CalcTempBus]          temp_b5_26_6_i;
wire signed [`CalcTempBus]          temp_b5_26_7_r;
wire signed [`CalcTempBus]          temp_b5_26_7_i;
wire signed [`CalcTempBus]          temp_b5_26_8_r;
wire signed [`CalcTempBus]          temp_b5_26_8_i;
wire signed [`CalcTempBus]          temp_b5_26_9_r;
wire signed [`CalcTempBus]          temp_b5_26_9_i;
wire signed [`CalcTempBus]          temp_b5_26_10_r;
wire signed [`CalcTempBus]          temp_b5_26_10_i;
wire signed [`CalcTempBus]          temp_b5_26_11_r;
wire signed [`CalcTempBus]          temp_b5_26_11_i;
wire signed [`CalcTempBus]          temp_b5_26_12_r;
wire signed [`CalcTempBus]          temp_b5_26_12_i;
wire signed [`CalcTempBus]          temp_b5_26_13_r;
wire signed [`CalcTempBus]          temp_b5_26_13_i;
wire signed [`CalcTempBus]          temp_b5_26_14_r;
wire signed [`CalcTempBus]          temp_b5_26_14_i;
wire signed [`CalcTempBus]          temp_b5_26_15_r;
wire signed [`CalcTempBus]          temp_b5_26_15_i;
wire signed [`CalcTempBus]          temp_b5_26_16_r;
wire signed [`CalcTempBus]          temp_b5_26_16_i;
wire signed [`CalcTempBus]          temp_b5_26_17_r;
wire signed [`CalcTempBus]          temp_b5_26_17_i;
wire signed [`CalcTempBus]          temp_b5_26_18_r;
wire signed [`CalcTempBus]          temp_b5_26_18_i;
wire signed [`CalcTempBus]          temp_b5_26_19_r;
wire signed [`CalcTempBus]          temp_b5_26_19_i;
wire signed [`CalcTempBus]          temp_b5_26_20_r;
wire signed [`CalcTempBus]          temp_b5_26_20_i;
wire signed [`CalcTempBus]          temp_b5_26_21_r;
wire signed [`CalcTempBus]          temp_b5_26_21_i;
wire signed [`CalcTempBus]          temp_b5_26_22_r;
wire signed [`CalcTempBus]          temp_b5_26_22_i;
wire signed [`CalcTempBus]          temp_b5_26_23_r;
wire signed [`CalcTempBus]          temp_b5_26_23_i;
wire signed [`CalcTempBus]          temp_b5_26_24_r;
wire signed [`CalcTempBus]          temp_b5_26_24_i;
wire signed [`CalcTempBus]          temp_b5_26_25_r;
wire signed [`CalcTempBus]          temp_b5_26_25_i;
wire signed [`CalcTempBus]          temp_b5_26_26_r;
wire signed [`CalcTempBus]          temp_b5_26_26_i;
wire signed [`CalcTempBus]          temp_b5_26_27_r;
wire signed [`CalcTempBus]          temp_b5_26_27_i;
wire signed [`CalcTempBus]          temp_b5_26_28_r;
wire signed [`CalcTempBus]          temp_b5_26_28_i;
wire signed [`CalcTempBus]          temp_b5_26_29_r;
wire signed [`CalcTempBus]          temp_b5_26_29_i;
wire signed [`CalcTempBus]          temp_b5_26_30_r;
wire signed [`CalcTempBus]          temp_b5_26_30_i;
wire signed [`CalcTempBus]          temp_b5_26_31_r;
wire signed [`CalcTempBus]          temp_b5_26_31_i;
wire signed [`CalcTempBus]          temp_b5_26_32_r;
wire signed [`CalcTempBus]          temp_b5_26_32_i;
wire signed [`CalcTempBus]          temp_b5_27_1_r;
wire signed [`CalcTempBus]          temp_b5_27_1_i;
wire signed [`CalcTempBus]          temp_b5_27_2_r;
wire signed [`CalcTempBus]          temp_b5_27_2_i;
wire signed [`CalcTempBus]          temp_b5_27_3_r;
wire signed [`CalcTempBus]          temp_b5_27_3_i;
wire signed [`CalcTempBus]          temp_b5_27_4_r;
wire signed [`CalcTempBus]          temp_b5_27_4_i;
wire signed [`CalcTempBus]          temp_b5_27_5_r;
wire signed [`CalcTempBus]          temp_b5_27_5_i;
wire signed [`CalcTempBus]          temp_b5_27_6_r;
wire signed [`CalcTempBus]          temp_b5_27_6_i;
wire signed [`CalcTempBus]          temp_b5_27_7_r;
wire signed [`CalcTempBus]          temp_b5_27_7_i;
wire signed [`CalcTempBus]          temp_b5_27_8_r;
wire signed [`CalcTempBus]          temp_b5_27_8_i;
wire signed [`CalcTempBus]          temp_b5_27_9_r;
wire signed [`CalcTempBus]          temp_b5_27_9_i;
wire signed [`CalcTempBus]          temp_b5_27_10_r;
wire signed [`CalcTempBus]          temp_b5_27_10_i;
wire signed [`CalcTempBus]          temp_b5_27_11_r;
wire signed [`CalcTempBus]          temp_b5_27_11_i;
wire signed [`CalcTempBus]          temp_b5_27_12_r;
wire signed [`CalcTempBus]          temp_b5_27_12_i;
wire signed [`CalcTempBus]          temp_b5_27_13_r;
wire signed [`CalcTempBus]          temp_b5_27_13_i;
wire signed [`CalcTempBus]          temp_b5_27_14_r;
wire signed [`CalcTempBus]          temp_b5_27_14_i;
wire signed [`CalcTempBus]          temp_b5_27_15_r;
wire signed [`CalcTempBus]          temp_b5_27_15_i;
wire signed [`CalcTempBus]          temp_b5_27_16_r;
wire signed [`CalcTempBus]          temp_b5_27_16_i;
wire signed [`CalcTempBus]          temp_b5_27_17_r;
wire signed [`CalcTempBus]          temp_b5_27_17_i;
wire signed [`CalcTempBus]          temp_b5_27_18_r;
wire signed [`CalcTempBus]          temp_b5_27_18_i;
wire signed [`CalcTempBus]          temp_b5_27_19_r;
wire signed [`CalcTempBus]          temp_b5_27_19_i;
wire signed [`CalcTempBus]          temp_b5_27_20_r;
wire signed [`CalcTempBus]          temp_b5_27_20_i;
wire signed [`CalcTempBus]          temp_b5_27_21_r;
wire signed [`CalcTempBus]          temp_b5_27_21_i;
wire signed [`CalcTempBus]          temp_b5_27_22_r;
wire signed [`CalcTempBus]          temp_b5_27_22_i;
wire signed [`CalcTempBus]          temp_b5_27_23_r;
wire signed [`CalcTempBus]          temp_b5_27_23_i;
wire signed [`CalcTempBus]          temp_b5_27_24_r;
wire signed [`CalcTempBus]          temp_b5_27_24_i;
wire signed [`CalcTempBus]          temp_b5_27_25_r;
wire signed [`CalcTempBus]          temp_b5_27_25_i;
wire signed [`CalcTempBus]          temp_b5_27_26_r;
wire signed [`CalcTempBus]          temp_b5_27_26_i;
wire signed [`CalcTempBus]          temp_b5_27_27_r;
wire signed [`CalcTempBus]          temp_b5_27_27_i;
wire signed [`CalcTempBus]          temp_b5_27_28_r;
wire signed [`CalcTempBus]          temp_b5_27_28_i;
wire signed [`CalcTempBus]          temp_b5_27_29_r;
wire signed [`CalcTempBus]          temp_b5_27_29_i;
wire signed [`CalcTempBus]          temp_b5_27_30_r;
wire signed [`CalcTempBus]          temp_b5_27_30_i;
wire signed [`CalcTempBus]          temp_b5_27_31_r;
wire signed [`CalcTempBus]          temp_b5_27_31_i;
wire signed [`CalcTempBus]          temp_b5_27_32_r;
wire signed [`CalcTempBus]          temp_b5_27_32_i;
wire signed [`CalcTempBus]          temp_b5_28_1_r;
wire signed [`CalcTempBus]          temp_b5_28_1_i;
wire signed [`CalcTempBus]          temp_b5_28_2_r;
wire signed [`CalcTempBus]          temp_b5_28_2_i;
wire signed [`CalcTempBus]          temp_b5_28_3_r;
wire signed [`CalcTempBus]          temp_b5_28_3_i;
wire signed [`CalcTempBus]          temp_b5_28_4_r;
wire signed [`CalcTempBus]          temp_b5_28_4_i;
wire signed [`CalcTempBus]          temp_b5_28_5_r;
wire signed [`CalcTempBus]          temp_b5_28_5_i;
wire signed [`CalcTempBus]          temp_b5_28_6_r;
wire signed [`CalcTempBus]          temp_b5_28_6_i;
wire signed [`CalcTempBus]          temp_b5_28_7_r;
wire signed [`CalcTempBus]          temp_b5_28_7_i;
wire signed [`CalcTempBus]          temp_b5_28_8_r;
wire signed [`CalcTempBus]          temp_b5_28_8_i;
wire signed [`CalcTempBus]          temp_b5_28_9_r;
wire signed [`CalcTempBus]          temp_b5_28_9_i;
wire signed [`CalcTempBus]          temp_b5_28_10_r;
wire signed [`CalcTempBus]          temp_b5_28_10_i;
wire signed [`CalcTempBus]          temp_b5_28_11_r;
wire signed [`CalcTempBus]          temp_b5_28_11_i;
wire signed [`CalcTempBus]          temp_b5_28_12_r;
wire signed [`CalcTempBus]          temp_b5_28_12_i;
wire signed [`CalcTempBus]          temp_b5_28_13_r;
wire signed [`CalcTempBus]          temp_b5_28_13_i;
wire signed [`CalcTempBus]          temp_b5_28_14_r;
wire signed [`CalcTempBus]          temp_b5_28_14_i;
wire signed [`CalcTempBus]          temp_b5_28_15_r;
wire signed [`CalcTempBus]          temp_b5_28_15_i;
wire signed [`CalcTempBus]          temp_b5_28_16_r;
wire signed [`CalcTempBus]          temp_b5_28_16_i;
wire signed [`CalcTempBus]          temp_b5_28_17_r;
wire signed [`CalcTempBus]          temp_b5_28_17_i;
wire signed [`CalcTempBus]          temp_b5_28_18_r;
wire signed [`CalcTempBus]          temp_b5_28_18_i;
wire signed [`CalcTempBus]          temp_b5_28_19_r;
wire signed [`CalcTempBus]          temp_b5_28_19_i;
wire signed [`CalcTempBus]          temp_b5_28_20_r;
wire signed [`CalcTempBus]          temp_b5_28_20_i;
wire signed [`CalcTempBus]          temp_b5_28_21_r;
wire signed [`CalcTempBus]          temp_b5_28_21_i;
wire signed [`CalcTempBus]          temp_b5_28_22_r;
wire signed [`CalcTempBus]          temp_b5_28_22_i;
wire signed [`CalcTempBus]          temp_b5_28_23_r;
wire signed [`CalcTempBus]          temp_b5_28_23_i;
wire signed [`CalcTempBus]          temp_b5_28_24_r;
wire signed [`CalcTempBus]          temp_b5_28_24_i;
wire signed [`CalcTempBus]          temp_b5_28_25_r;
wire signed [`CalcTempBus]          temp_b5_28_25_i;
wire signed [`CalcTempBus]          temp_b5_28_26_r;
wire signed [`CalcTempBus]          temp_b5_28_26_i;
wire signed [`CalcTempBus]          temp_b5_28_27_r;
wire signed [`CalcTempBus]          temp_b5_28_27_i;
wire signed [`CalcTempBus]          temp_b5_28_28_r;
wire signed [`CalcTempBus]          temp_b5_28_28_i;
wire signed [`CalcTempBus]          temp_b5_28_29_r;
wire signed [`CalcTempBus]          temp_b5_28_29_i;
wire signed [`CalcTempBus]          temp_b5_28_30_r;
wire signed [`CalcTempBus]          temp_b5_28_30_i;
wire signed [`CalcTempBus]          temp_b5_28_31_r;
wire signed [`CalcTempBus]          temp_b5_28_31_i;
wire signed [`CalcTempBus]          temp_b5_28_32_r;
wire signed [`CalcTempBus]          temp_b5_28_32_i;
wire signed [`CalcTempBus]          temp_b5_29_1_r;
wire signed [`CalcTempBus]          temp_b5_29_1_i;
wire signed [`CalcTempBus]          temp_b5_29_2_r;
wire signed [`CalcTempBus]          temp_b5_29_2_i;
wire signed [`CalcTempBus]          temp_b5_29_3_r;
wire signed [`CalcTempBus]          temp_b5_29_3_i;
wire signed [`CalcTempBus]          temp_b5_29_4_r;
wire signed [`CalcTempBus]          temp_b5_29_4_i;
wire signed [`CalcTempBus]          temp_b5_29_5_r;
wire signed [`CalcTempBus]          temp_b5_29_5_i;
wire signed [`CalcTempBus]          temp_b5_29_6_r;
wire signed [`CalcTempBus]          temp_b5_29_6_i;
wire signed [`CalcTempBus]          temp_b5_29_7_r;
wire signed [`CalcTempBus]          temp_b5_29_7_i;
wire signed [`CalcTempBus]          temp_b5_29_8_r;
wire signed [`CalcTempBus]          temp_b5_29_8_i;
wire signed [`CalcTempBus]          temp_b5_29_9_r;
wire signed [`CalcTempBus]          temp_b5_29_9_i;
wire signed [`CalcTempBus]          temp_b5_29_10_r;
wire signed [`CalcTempBus]          temp_b5_29_10_i;
wire signed [`CalcTempBus]          temp_b5_29_11_r;
wire signed [`CalcTempBus]          temp_b5_29_11_i;
wire signed [`CalcTempBus]          temp_b5_29_12_r;
wire signed [`CalcTempBus]          temp_b5_29_12_i;
wire signed [`CalcTempBus]          temp_b5_29_13_r;
wire signed [`CalcTempBus]          temp_b5_29_13_i;
wire signed [`CalcTempBus]          temp_b5_29_14_r;
wire signed [`CalcTempBus]          temp_b5_29_14_i;
wire signed [`CalcTempBus]          temp_b5_29_15_r;
wire signed [`CalcTempBus]          temp_b5_29_15_i;
wire signed [`CalcTempBus]          temp_b5_29_16_r;
wire signed [`CalcTempBus]          temp_b5_29_16_i;
wire signed [`CalcTempBus]          temp_b5_29_17_r;
wire signed [`CalcTempBus]          temp_b5_29_17_i;
wire signed [`CalcTempBus]          temp_b5_29_18_r;
wire signed [`CalcTempBus]          temp_b5_29_18_i;
wire signed [`CalcTempBus]          temp_b5_29_19_r;
wire signed [`CalcTempBus]          temp_b5_29_19_i;
wire signed [`CalcTempBus]          temp_b5_29_20_r;
wire signed [`CalcTempBus]          temp_b5_29_20_i;
wire signed [`CalcTempBus]          temp_b5_29_21_r;
wire signed [`CalcTempBus]          temp_b5_29_21_i;
wire signed [`CalcTempBus]          temp_b5_29_22_r;
wire signed [`CalcTempBus]          temp_b5_29_22_i;
wire signed [`CalcTempBus]          temp_b5_29_23_r;
wire signed [`CalcTempBus]          temp_b5_29_23_i;
wire signed [`CalcTempBus]          temp_b5_29_24_r;
wire signed [`CalcTempBus]          temp_b5_29_24_i;
wire signed [`CalcTempBus]          temp_b5_29_25_r;
wire signed [`CalcTempBus]          temp_b5_29_25_i;
wire signed [`CalcTempBus]          temp_b5_29_26_r;
wire signed [`CalcTempBus]          temp_b5_29_26_i;
wire signed [`CalcTempBus]          temp_b5_29_27_r;
wire signed [`CalcTempBus]          temp_b5_29_27_i;
wire signed [`CalcTempBus]          temp_b5_29_28_r;
wire signed [`CalcTempBus]          temp_b5_29_28_i;
wire signed [`CalcTempBus]          temp_b5_29_29_r;
wire signed [`CalcTempBus]          temp_b5_29_29_i;
wire signed [`CalcTempBus]          temp_b5_29_30_r;
wire signed [`CalcTempBus]          temp_b5_29_30_i;
wire signed [`CalcTempBus]          temp_b5_29_31_r;
wire signed [`CalcTempBus]          temp_b5_29_31_i;
wire signed [`CalcTempBus]          temp_b5_29_32_r;
wire signed [`CalcTempBus]          temp_b5_29_32_i;
wire signed [`CalcTempBus]          temp_b5_30_1_r;
wire signed [`CalcTempBus]          temp_b5_30_1_i;
wire signed [`CalcTempBus]          temp_b5_30_2_r;
wire signed [`CalcTempBus]          temp_b5_30_2_i;
wire signed [`CalcTempBus]          temp_b5_30_3_r;
wire signed [`CalcTempBus]          temp_b5_30_3_i;
wire signed [`CalcTempBus]          temp_b5_30_4_r;
wire signed [`CalcTempBus]          temp_b5_30_4_i;
wire signed [`CalcTempBus]          temp_b5_30_5_r;
wire signed [`CalcTempBus]          temp_b5_30_5_i;
wire signed [`CalcTempBus]          temp_b5_30_6_r;
wire signed [`CalcTempBus]          temp_b5_30_6_i;
wire signed [`CalcTempBus]          temp_b5_30_7_r;
wire signed [`CalcTempBus]          temp_b5_30_7_i;
wire signed [`CalcTempBus]          temp_b5_30_8_r;
wire signed [`CalcTempBus]          temp_b5_30_8_i;
wire signed [`CalcTempBus]          temp_b5_30_9_r;
wire signed [`CalcTempBus]          temp_b5_30_9_i;
wire signed [`CalcTempBus]          temp_b5_30_10_r;
wire signed [`CalcTempBus]          temp_b5_30_10_i;
wire signed [`CalcTempBus]          temp_b5_30_11_r;
wire signed [`CalcTempBus]          temp_b5_30_11_i;
wire signed [`CalcTempBus]          temp_b5_30_12_r;
wire signed [`CalcTempBus]          temp_b5_30_12_i;
wire signed [`CalcTempBus]          temp_b5_30_13_r;
wire signed [`CalcTempBus]          temp_b5_30_13_i;
wire signed [`CalcTempBus]          temp_b5_30_14_r;
wire signed [`CalcTempBus]          temp_b5_30_14_i;
wire signed [`CalcTempBus]          temp_b5_30_15_r;
wire signed [`CalcTempBus]          temp_b5_30_15_i;
wire signed [`CalcTempBus]          temp_b5_30_16_r;
wire signed [`CalcTempBus]          temp_b5_30_16_i;
wire signed [`CalcTempBus]          temp_b5_30_17_r;
wire signed [`CalcTempBus]          temp_b5_30_17_i;
wire signed [`CalcTempBus]          temp_b5_30_18_r;
wire signed [`CalcTempBus]          temp_b5_30_18_i;
wire signed [`CalcTempBus]          temp_b5_30_19_r;
wire signed [`CalcTempBus]          temp_b5_30_19_i;
wire signed [`CalcTempBus]          temp_b5_30_20_r;
wire signed [`CalcTempBus]          temp_b5_30_20_i;
wire signed [`CalcTempBus]          temp_b5_30_21_r;
wire signed [`CalcTempBus]          temp_b5_30_21_i;
wire signed [`CalcTempBus]          temp_b5_30_22_r;
wire signed [`CalcTempBus]          temp_b5_30_22_i;
wire signed [`CalcTempBus]          temp_b5_30_23_r;
wire signed [`CalcTempBus]          temp_b5_30_23_i;
wire signed [`CalcTempBus]          temp_b5_30_24_r;
wire signed [`CalcTempBus]          temp_b5_30_24_i;
wire signed [`CalcTempBus]          temp_b5_30_25_r;
wire signed [`CalcTempBus]          temp_b5_30_25_i;
wire signed [`CalcTempBus]          temp_b5_30_26_r;
wire signed [`CalcTempBus]          temp_b5_30_26_i;
wire signed [`CalcTempBus]          temp_b5_30_27_r;
wire signed [`CalcTempBus]          temp_b5_30_27_i;
wire signed [`CalcTempBus]          temp_b5_30_28_r;
wire signed [`CalcTempBus]          temp_b5_30_28_i;
wire signed [`CalcTempBus]          temp_b5_30_29_r;
wire signed [`CalcTempBus]          temp_b5_30_29_i;
wire signed [`CalcTempBus]          temp_b5_30_30_r;
wire signed [`CalcTempBus]          temp_b5_30_30_i;
wire signed [`CalcTempBus]          temp_b5_30_31_r;
wire signed [`CalcTempBus]          temp_b5_30_31_i;
wire signed [`CalcTempBus]          temp_b5_30_32_r;
wire signed [`CalcTempBus]          temp_b5_30_32_i;
wire signed [`CalcTempBus]          temp_b5_31_1_r;
wire signed [`CalcTempBus]          temp_b5_31_1_i;
wire signed [`CalcTempBus]          temp_b5_31_2_r;
wire signed [`CalcTempBus]          temp_b5_31_2_i;
wire signed [`CalcTempBus]          temp_b5_31_3_r;
wire signed [`CalcTempBus]          temp_b5_31_3_i;
wire signed [`CalcTempBus]          temp_b5_31_4_r;
wire signed [`CalcTempBus]          temp_b5_31_4_i;
wire signed [`CalcTempBus]          temp_b5_31_5_r;
wire signed [`CalcTempBus]          temp_b5_31_5_i;
wire signed [`CalcTempBus]          temp_b5_31_6_r;
wire signed [`CalcTempBus]          temp_b5_31_6_i;
wire signed [`CalcTempBus]          temp_b5_31_7_r;
wire signed [`CalcTempBus]          temp_b5_31_7_i;
wire signed [`CalcTempBus]          temp_b5_31_8_r;
wire signed [`CalcTempBus]          temp_b5_31_8_i;
wire signed [`CalcTempBus]          temp_b5_31_9_r;
wire signed [`CalcTempBus]          temp_b5_31_9_i;
wire signed [`CalcTempBus]          temp_b5_31_10_r;
wire signed [`CalcTempBus]          temp_b5_31_10_i;
wire signed [`CalcTempBus]          temp_b5_31_11_r;
wire signed [`CalcTempBus]          temp_b5_31_11_i;
wire signed [`CalcTempBus]          temp_b5_31_12_r;
wire signed [`CalcTempBus]          temp_b5_31_12_i;
wire signed [`CalcTempBus]          temp_b5_31_13_r;
wire signed [`CalcTempBus]          temp_b5_31_13_i;
wire signed [`CalcTempBus]          temp_b5_31_14_r;
wire signed [`CalcTempBus]          temp_b5_31_14_i;
wire signed [`CalcTempBus]          temp_b5_31_15_r;
wire signed [`CalcTempBus]          temp_b5_31_15_i;
wire signed [`CalcTempBus]          temp_b5_31_16_r;
wire signed [`CalcTempBus]          temp_b5_31_16_i;
wire signed [`CalcTempBus]          temp_b5_31_17_r;
wire signed [`CalcTempBus]          temp_b5_31_17_i;
wire signed [`CalcTempBus]          temp_b5_31_18_r;
wire signed [`CalcTempBus]          temp_b5_31_18_i;
wire signed [`CalcTempBus]          temp_b5_31_19_r;
wire signed [`CalcTempBus]          temp_b5_31_19_i;
wire signed [`CalcTempBus]          temp_b5_31_20_r;
wire signed [`CalcTempBus]          temp_b5_31_20_i;
wire signed [`CalcTempBus]          temp_b5_31_21_r;
wire signed [`CalcTempBus]          temp_b5_31_21_i;
wire signed [`CalcTempBus]          temp_b5_31_22_r;
wire signed [`CalcTempBus]          temp_b5_31_22_i;
wire signed [`CalcTempBus]          temp_b5_31_23_r;
wire signed [`CalcTempBus]          temp_b5_31_23_i;
wire signed [`CalcTempBus]          temp_b5_31_24_r;
wire signed [`CalcTempBus]          temp_b5_31_24_i;
wire signed [`CalcTempBus]          temp_b5_31_25_r;
wire signed [`CalcTempBus]          temp_b5_31_25_i;
wire signed [`CalcTempBus]          temp_b5_31_26_r;
wire signed [`CalcTempBus]          temp_b5_31_26_i;
wire signed [`CalcTempBus]          temp_b5_31_27_r;
wire signed [`CalcTempBus]          temp_b5_31_27_i;
wire signed [`CalcTempBus]          temp_b5_31_28_r;
wire signed [`CalcTempBus]          temp_b5_31_28_i;
wire signed [`CalcTempBus]          temp_b5_31_29_r;
wire signed [`CalcTempBus]          temp_b5_31_29_i;
wire signed [`CalcTempBus]          temp_b5_31_30_r;
wire signed [`CalcTempBus]          temp_b5_31_30_i;
wire signed [`CalcTempBus]          temp_b5_31_31_r;
wire signed [`CalcTempBus]          temp_b5_31_31_i;
wire signed [`CalcTempBus]          temp_b5_31_32_r;
wire signed [`CalcTempBus]          temp_b5_31_32_i;
wire signed [`CalcTempBus]          temp_b5_32_1_r;
wire signed [`CalcTempBus]          temp_b5_32_1_i;
wire signed [`CalcTempBus]          temp_b5_32_2_r;
wire signed [`CalcTempBus]          temp_b5_32_2_i;
wire signed [`CalcTempBus]          temp_b5_32_3_r;
wire signed [`CalcTempBus]          temp_b5_32_3_i;
wire signed [`CalcTempBus]          temp_b5_32_4_r;
wire signed [`CalcTempBus]          temp_b5_32_4_i;
wire signed [`CalcTempBus]          temp_b5_32_5_r;
wire signed [`CalcTempBus]          temp_b5_32_5_i;
wire signed [`CalcTempBus]          temp_b5_32_6_r;
wire signed [`CalcTempBus]          temp_b5_32_6_i;
wire signed [`CalcTempBus]          temp_b5_32_7_r;
wire signed [`CalcTempBus]          temp_b5_32_7_i;
wire signed [`CalcTempBus]          temp_b5_32_8_r;
wire signed [`CalcTempBus]          temp_b5_32_8_i;
wire signed [`CalcTempBus]          temp_b5_32_9_r;
wire signed [`CalcTempBus]          temp_b5_32_9_i;
wire signed [`CalcTempBus]          temp_b5_32_10_r;
wire signed [`CalcTempBus]          temp_b5_32_10_i;
wire signed [`CalcTempBus]          temp_b5_32_11_r;
wire signed [`CalcTempBus]          temp_b5_32_11_i;
wire signed [`CalcTempBus]          temp_b5_32_12_r;
wire signed [`CalcTempBus]          temp_b5_32_12_i;
wire signed [`CalcTempBus]          temp_b5_32_13_r;
wire signed [`CalcTempBus]          temp_b5_32_13_i;
wire signed [`CalcTempBus]          temp_b5_32_14_r;
wire signed [`CalcTempBus]          temp_b5_32_14_i;
wire signed [`CalcTempBus]          temp_b5_32_15_r;
wire signed [`CalcTempBus]          temp_b5_32_15_i;
wire signed [`CalcTempBus]          temp_b5_32_16_r;
wire signed [`CalcTempBus]          temp_b5_32_16_i;
wire signed [`CalcTempBus]          temp_b5_32_17_r;
wire signed [`CalcTempBus]          temp_b5_32_17_i;
wire signed [`CalcTempBus]          temp_b5_32_18_r;
wire signed [`CalcTempBus]          temp_b5_32_18_i;
wire signed [`CalcTempBus]          temp_b5_32_19_r;
wire signed [`CalcTempBus]          temp_b5_32_19_i;
wire signed [`CalcTempBus]          temp_b5_32_20_r;
wire signed [`CalcTempBus]          temp_b5_32_20_i;
wire signed [`CalcTempBus]          temp_b5_32_21_r;
wire signed [`CalcTempBus]          temp_b5_32_21_i;
wire signed [`CalcTempBus]          temp_b5_32_22_r;
wire signed [`CalcTempBus]          temp_b5_32_22_i;
wire signed [`CalcTempBus]          temp_b5_32_23_r;
wire signed [`CalcTempBus]          temp_b5_32_23_i;
wire signed [`CalcTempBus]          temp_b5_32_24_r;
wire signed [`CalcTempBus]          temp_b5_32_24_i;
wire signed [`CalcTempBus]          temp_b5_32_25_r;
wire signed [`CalcTempBus]          temp_b5_32_25_i;
wire signed [`CalcTempBus]          temp_b5_32_26_r;
wire signed [`CalcTempBus]          temp_b5_32_26_i;
wire signed [`CalcTempBus]          temp_b5_32_27_r;
wire signed [`CalcTempBus]          temp_b5_32_27_i;
wire signed [`CalcTempBus]          temp_b5_32_28_r;
wire signed [`CalcTempBus]          temp_b5_32_28_i;
wire signed [`CalcTempBus]          temp_b5_32_29_r;
wire signed [`CalcTempBus]          temp_b5_32_29_i;
wire signed [`CalcTempBus]          temp_b5_32_30_r;
wire signed [`CalcTempBus]          temp_b5_32_30_i;
wire signed [`CalcTempBus]          temp_b5_32_31_r;
wire signed [`CalcTempBus]          temp_b5_32_31_i;
wire signed [`CalcTempBus]          temp_b5_32_32_r;
wire signed [`CalcTempBus]          temp_b5_32_32_i;

/******************port map******************/
MULT MULT1 (clk,in_1_1_r,in_1_1_i,in_1_2_r,in_1_2_i,in_2_1_r,in_2_1_i,in_2_2_r,in_2_2_i,temp_m1_1_1_r,temp_m1_1_1_i,temp_m1_1_2_r,temp_m1_1_2_i,temp_m1_2_1_r,temp_m1_2_1_i,temp_m1_2_2_r,temp_m1_2_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly1 (clk,temp_m1_1_1_r,temp_m1_1_1_i,temp_m1_1_2_r,temp_m1_1_2_i,temp_m1_2_1_r,temp_m1_2_1_i,temp_m1_2_2_r,temp_m1_2_2_i,temp_b1_1_1_r,temp_b1_1_1_i,temp_b1_1_2_r,temp_b1_1_2_i,temp_b1_2_1_r,temp_b1_2_1_i,temp_b1_2_2_r,temp_b1_2_2_i);
MULT MULT2 (clk,in_1_3_r,in_1_3_i,in_1_4_r,in_1_4_i,in_2_3_r,in_2_3_i,in_2_4_r,in_2_4_i,temp_m1_1_3_r,temp_m1_1_3_i,temp_m1_1_4_r,temp_m1_1_4_i,temp_m1_2_3_r,temp_m1_2_3_i,temp_m1_2_4_r,temp_m1_2_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly2 (clk,temp_m1_1_3_r,temp_m1_1_3_i,temp_m1_1_4_r,temp_m1_1_4_i,temp_m1_2_3_r,temp_m1_2_3_i,temp_m1_2_4_r,temp_m1_2_4_i,temp_b1_1_3_r,temp_b1_1_3_i,temp_b1_1_4_r,temp_b1_1_4_i,temp_b1_2_3_r,temp_b1_2_3_i,temp_b1_2_4_r,temp_b1_2_4_i);
MULT MULT3 (clk,in_1_5_r,in_1_5_i,in_1_6_r,in_1_6_i,in_2_5_r,in_2_5_i,in_2_6_r,in_2_6_i,temp_m1_1_5_r,temp_m1_1_5_i,temp_m1_1_6_r,temp_m1_1_6_i,temp_m1_2_5_r,temp_m1_2_5_i,temp_m1_2_6_r,temp_m1_2_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly3 (clk,temp_m1_1_5_r,temp_m1_1_5_i,temp_m1_1_6_r,temp_m1_1_6_i,temp_m1_2_5_r,temp_m1_2_5_i,temp_m1_2_6_r,temp_m1_2_6_i,temp_b1_1_5_r,temp_b1_1_5_i,temp_b1_1_6_r,temp_b1_1_6_i,temp_b1_2_5_r,temp_b1_2_5_i,temp_b1_2_6_r,temp_b1_2_6_i);
MULT MULT4 (clk,in_1_7_r,in_1_7_i,in_1_8_r,in_1_8_i,in_2_7_r,in_2_7_i,in_2_8_r,in_2_8_i,temp_m1_1_7_r,temp_m1_1_7_i,temp_m1_1_8_r,temp_m1_1_8_i,temp_m1_2_7_r,temp_m1_2_7_i,temp_m1_2_8_r,temp_m1_2_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly4 (clk,temp_m1_1_7_r,temp_m1_1_7_i,temp_m1_1_8_r,temp_m1_1_8_i,temp_m1_2_7_r,temp_m1_2_7_i,temp_m1_2_8_r,temp_m1_2_8_i,temp_b1_1_7_r,temp_b1_1_7_i,temp_b1_1_8_r,temp_b1_1_8_i,temp_b1_2_7_r,temp_b1_2_7_i,temp_b1_2_8_r,temp_b1_2_8_i);
MULT MULT5 (clk,in_1_9_r,in_1_9_i,in_1_10_r,in_1_10_i,in_2_9_r,in_2_9_i,in_2_10_r,in_2_10_i,temp_m1_1_9_r,temp_m1_1_9_i,temp_m1_1_10_r,temp_m1_1_10_i,temp_m1_2_9_r,temp_m1_2_9_i,temp_m1_2_10_r,temp_m1_2_10_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly5 (clk,temp_m1_1_9_r,temp_m1_1_9_i,temp_m1_1_10_r,temp_m1_1_10_i,temp_m1_2_9_r,temp_m1_2_9_i,temp_m1_2_10_r,temp_m1_2_10_i,temp_b1_1_9_r,temp_b1_1_9_i,temp_b1_1_10_r,temp_b1_1_10_i,temp_b1_2_9_r,temp_b1_2_9_i,temp_b1_2_10_r,temp_b1_2_10_i);
MULT MULT6 (clk,in_1_11_r,in_1_11_i,in_1_12_r,in_1_12_i,in_2_11_r,in_2_11_i,in_2_12_r,in_2_12_i,temp_m1_1_11_r,temp_m1_1_11_i,temp_m1_1_12_r,temp_m1_1_12_i,temp_m1_2_11_r,temp_m1_2_11_i,temp_m1_2_12_r,temp_m1_2_12_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly6 (clk,temp_m1_1_11_r,temp_m1_1_11_i,temp_m1_1_12_r,temp_m1_1_12_i,temp_m1_2_11_r,temp_m1_2_11_i,temp_m1_2_12_r,temp_m1_2_12_i,temp_b1_1_11_r,temp_b1_1_11_i,temp_b1_1_12_r,temp_b1_1_12_i,temp_b1_2_11_r,temp_b1_2_11_i,temp_b1_2_12_r,temp_b1_2_12_i);
MULT MULT7 (clk,in_1_13_r,in_1_13_i,in_1_14_r,in_1_14_i,in_2_13_r,in_2_13_i,in_2_14_r,in_2_14_i,temp_m1_1_13_r,temp_m1_1_13_i,temp_m1_1_14_r,temp_m1_1_14_i,temp_m1_2_13_r,temp_m1_2_13_i,temp_m1_2_14_r,temp_m1_2_14_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly7 (clk,temp_m1_1_13_r,temp_m1_1_13_i,temp_m1_1_14_r,temp_m1_1_14_i,temp_m1_2_13_r,temp_m1_2_13_i,temp_m1_2_14_r,temp_m1_2_14_i,temp_b1_1_13_r,temp_b1_1_13_i,temp_b1_1_14_r,temp_b1_1_14_i,temp_b1_2_13_r,temp_b1_2_13_i,temp_b1_2_14_r,temp_b1_2_14_i);
MULT MULT8 (clk,in_1_15_r,in_1_15_i,in_1_16_r,in_1_16_i,in_2_15_r,in_2_15_i,in_2_16_r,in_2_16_i,temp_m1_1_15_r,temp_m1_1_15_i,temp_m1_1_16_r,temp_m1_1_16_i,temp_m1_2_15_r,temp_m1_2_15_i,temp_m1_2_16_r,temp_m1_2_16_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly8 (clk,temp_m1_1_15_r,temp_m1_1_15_i,temp_m1_1_16_r,temp_m1_1_16_i,temp_m1_2_15_r,temp_m1_2_15_i,temp_m1_2_16_r,temp_m1_2_16_i,temp_b1_1_15_r,temp_b1_1_15_i,temp_b1_1_16_r,temp_b1_1_16_i,temp_b1_2_15_r,temp_b1_2_15_i,temp_b1_2_16_r,temp_b1_2_16_i);
MULT MULT9 (clk,in_1_17_r,in_1_17_i,in_1_18_r,in_1_18_i,in_2_17_r,in_2_17_i,in_2_18_r,in_2_18_i,temp_m1_1_17_r,temp_m1_1_17_i,temp_m1_1_18_r,temp_m1_1_18_i,temp_m1_2_17_r,temp_m1_2_17_i,temp_m1_2_18_r,temp_m1_2_18_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly9 (clk,temp_m1_1_17_r,temp_m1_1_17_i,temp_m1_1_18_r,temp_m1_1_18_i,temp_m1_2_17_r,temp_m1_2_17_i,temp_m1_2_18_r,temp_m1_2_18_i,temp_b1_1_17_r,temp_b1_1_17_i,temp_b1_1_18_r,temp_b1_1_18_i,temp_b1_2_17_r,temp_b1_2_17_i,temp_b1_2_18_r,temp_b1_2_18_i);
MULT MULT10 (clk,in_1_19_r,in_1_19_i,in_1_20_r,in_1_20_i,in_2_19_r,in_2_19_i,in_2_20_r,in_2_20_i,temp_m1_1_19_r,temp_m1_1_19_i,temp_m1_1_20_r,temp_m1_1_20_i,temp_m1_2_19_r,temp_m1_2_19_i,temp_m1_2_20_r,temp_m1_2_20_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly10 (clk,temp_m1_1_19_r,temp_m1_1_19_i,temp_m1_1_20_r,temp_m1_1_20_i,temp_m1_2_19_r,temp_m1_2_19_i,temp_m1_2_20_r,temp_m1_2_20_i,temp_b1_1_19_r,temp_b1_1_19_i,temp_b1_1_20_r,temp_b1_1_20_i,temp_b1_2_19_r,temp_b1_2_19_i,temp_b1_2_20_r,temp_b1_2_20_i);
MULT MULT11 (clk,in_1_21_r,in_1_21_i,in_1_22_r,in_1_22_i,in_2_21_r,in_2_21_i,in_2_22_r,in_2_22_i,temp_m1_1_21_r,temp_m1_1_21_i,temp_m1_1_22_r,temp_m1_1_22_i,temp_m1_2_21_r,temp_m1_2_21_i,temp_m1_2_22_r,temp_m1_2_22_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly11 (clk,temp_m1_1_21_r,temp_m1_1_21_i,temp_m1_1_22_r,temp_m1_1_22_i,temp_m1_2_21_r,temp_m1_2_21_i,temp_m1_2_22_r,temp_m1_2_22_i,temp_b1_1_21_r,temp_b1_1_21_i,temp_b1_1_22_r,temp_b1_1_22_i,temp_b1_2_21_r,temp_b1_2_21_i,temp_b1_2_22_r,temp_b1_2_22_i);
MULT MULT12 (clk,in_1_23_r,in_1_23_i,in_1_24_r,in_1_24_i,in_2_23_r,in_2_23_i,in_2_24_r,in_2_24_i,temp_m1_1_23_r,temp_m1_1_23_i,temp_m1_1_24_r,temp_m1_1_24_i,temp_m1_2_23_r,temp_m1_2_23_i,temp_m1_2_24_r,temp_m1_2_24_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly12 (clk,temp_m1_1_23_r,temp_m1_1_23_i,temp_m1_1_24_r,temp_m1_1_24_i,temp_m1_2_23_r,temp_m1_2_23_i,temp_m1_2_24_r,temp_m1_2_24_i,temp_b1_1_23_r,temp_b1_1_23_i,temp_b1_1_24_r,temp_b1_1_24_i,temp_b1_2_23_r,temp_b1_2_23_i,temp_b1_2_24_r,temp_b1_2_24_i);
MULT MULT13 (clk,in_1_25_r,in_1_25_i,in_1_26_r,in_1_26_i,in_2_25_r,in_2_25_i,in_2_26_r,in_2_26_i,temp_m1_1_25_r,temp_m1_1_25_i,temp_m1_1_26_r,temp_m1_1_26_i,temp_m1_2_25_r,temp_m1_2_25_i,temp_m1_2_26_r,temp_m1_2_26_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly13 (clk,temp_m1_1_25_r,temp_m1_1_25_i,temp_m1_1_26_r,temp_m1_1_26_i,temp_m1_2_25_r,temp_m1_2_25_i,temp_m1_2_26_r,temp_m1_2_26_i,temp_b1_1_25_r,temp_b1_1_25_i,temp_b1_1_26_r,temp_b1_1_26_i,temp_b1_2_25_r,temp_b1_2_25_i,temp_b1_2_26_r,temp_b1_2_26_i);
MULT MULT14 (clk,in_1_27_r,in_1_27_i,in_1_28_r,in_1_28_i,in_2_27_r,in_2_27_i,in_2_28_r,in_2_28_i,temp_m1_1_27_r,temp_m1_1_27_i,temp_m1_1_28_r,temp_m1_1_28_i,temp_m1_2_27_r,temp_m1_2_27_i,temp_m1_2_28_r,temp_m1_2_28_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly14 (clk,temp_m1_1_27_r,temp_m1_1_27_i,temp_m1_1_28_r,temp_m1_1_28_i,temp_m1_2_27_r,temp_m1_2_27_i,temp_m1_2_28_r,temp_m1_2_28_i,temp_b1_1_27_r,temp_b1_1_27_i,temp_b1_1_28_r,temp_b1_1_28_i,temp_b1_2_27_r,temp_b1_2_27_i,temp_b1_2_28_r,temp_b1_2_28_i);
MULT MULT15 (clk,in_1_29_r,in_1_29_i,in_1_30_r,in_1_30_i,in_2_29_r,in_2_29_i,in_2_30_r,in_2_30_i,temp_m1_1_29_r,temp_m1_1_29_i,temp_m1_1_30_r,temp_m1_1_30_i,temp_m1_2_29_r,temp_m1_2_29_i,temp_m1_2_30_r,temp_m1_2_30_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly15 (clk,temp_m1_1_29_r,temp_m1_1_29_i,temp_m1_1_30_r,temp_m1_1_30_i,temp_m1_2_29_r,temp_m1_2_29_i,temp_m1_2_30_r,temp_m1_2_30_i,temp_b1_1_29_r,temp_b1_1_29_i,temp_b1_1_30_r,temp_b1_1_30_i,temp_b1_2_29_r,temp_b1_2_29_i,temp_b1_2_30_r,temp_b1_2_30_i);
MULT MULT16 (clk,in_1_31_r,in_1_31_i,in_1_32_r,in_1_32_i,in_2_31_r,in_2_31_i,in_2_32_r,in_2_32_i,temp_m1_1_31_r,temp_m1_1_31_i,temp_m1_1_32_r,temp_m1_1_32_i,temp_m1_2_31_r,temp_m1_2_31_i,temp_m1_2_32_r,temp_m1_2_32_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly16 (clk,temp_m1_1_31_r,temp_m1_1_31_i,temp_m1_1_32_r,temp_m1_1_32_i,temp_m1_2_31_r,temp_m1_2_31_i,temp_m1_2_32_r,temp_m1_2_32_i,temp_b1_1_31_r,temp_b1_1_31_i,temp_b1_1_32_r,temp_b1_1_32_i,temp_b1_2_31_r,temp_b1_2_31_i,temp_b1_2_32_r,temp_b1_2_32_i);
MULT MULT17 (clk,in_3_1_r,in_3_1_i,in_3_2_r,in_3_2_i,in_4_1_r,in_4_1_i,in_4_2_r,in_4_2_i,temp_m1_3_1_r,temp_m1_3_1_i,temp_m1_3_2_r,temp_m1_3_2_i,temp_m1_4_1_r,temp_m1_4_1_i,temp_m1_4_2_r,temp_m1_4_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly17 (clk,temp_m1_3_1_r,temp_m1_3_1_i,temp_m1_3_2_r,temp_m1_3_2_i,temp_m1_4_1_r,temp_m1_4_1_i,temp_m1_4_2_r,temp_m1_4_2_i,temp_b1_3_1_r,temp_b1_3_1_i,temp_b1_3_2_r,temp_b1_3_2_i,temp_b1_4_1_r,temp_b1_4_1_i,temp_b1_4_2_r,temp_b1_4_2_i);
MULT MULT18 (clk,in_3_3_r,in_3_3_i,in_3_4_r,in_3_4_i,in_4_3_r,in_4_3_i,in_4_4_r,in_4_4_i,temp_m1_3_3_r,temp_m1_3_3_i,temp_m1_3_4_r,temp_m1_3_4_i,temp_m1_4_3_r,temp_m1_4_3_i,temp_m1_4_4_r,temp_m1_4_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly18 (clk,temp_m1_3_3_r,temp_m1_3_3_i,temp_m1_3_4_r,temp_m1_3_4_i,temp_m1_4_3_r,temp_m1_4_3_i,temp_m1_4_4_r,temp_m1_4_4_i,temp_b1_3_3_r,temp_b1_3_3_i,temp_b1_3_4_r,temp_b1_3_4_i,temp_b1_4_3_r,temp_b1_4_3_i,temp_b1_4_4_r,temp_b1_4_4_i);
MULT MULT19 (clk,in_3_5_r,in_3_5_i,in_3_6_r,in_3_6_i,in_4_5_r,in_4_5_i,in_4_6_r,in_4_6_i,temp_m1_3_5_r,temp_m1_3_5_i,temp_m1_3_6_r,temp_m1_3_6_i,temp_m1_4_5_r,temp_m1_4_5_i,temp_m1_4_6_r,temp_m1_4_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly19 (clk,temp_m1_3_5_r,temp_m1_3_5_i,temp_m1_3_6_r,temp_m1_3_6_i,temp_m1_4_5_r,temp_m1_4_5_i,temp_m1_4_6_r,temp_m1_4_6_i,temp_b1_3_5_r,temp_b1_3_5_i,temp_b1_3_6_r,temp_b1_3_6_i,temp_b1_4_5_r,temp_b1_4_5_i,temp_b1_4_6_r,temp_b1_4_6_i);
MULT MULT20 (clk,in_3_7_r,in_3_7_i,in_3_8_r,in_3_8_i,in_4_7_r,in_4_7_i,in_4_8_r,in_4_8_i,temp_m1_3_7_r,temp_m1_3_7_i,temp_m1_3_8_r,temp_m1_3_8_i,temp_m1_4_7_r,temp_m1_4_7_i,temp_m1_4_8_r,temp_m1_4_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly20 (clk,temp_m1_3_7_r,temp_m1_3_7_i,temp_m1_3_8_r,temp_m1_3_8_i,temp_m1_4_7_r,temp_m1_4_7_i,temp_m1_4_8_r,temp_m1_4_8_i,temp_b1_3_7_r,temp_b1_3_7_i,temp_b1_3_8_r,temp_b1_3_8_i,temp_b1_4_7_r,temp_b1_4_7_i,temp_b1_4_8_r,temp_b1_4_8_i);
MULT MULT21 (clk,in_3_9_r,in_3_9_i,in_3_10_r,in_3_10_i,in_4_9_r,in_4_9_i,in_4_10_r,in_4_10_i,temp_m1_3_9_r,temp_m1_3_9_i,temp_m1_3_10_r,temp_m1_3_10_i,temp_m1_4_9_r,temp_m1_4_9_i,temp_m1_4_10_r,temp_m1_4_10_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly21 (clk,temp_m1_3_9_r,temp_m1_3_9_i,temp_m1_3_10_r,temp_m1_3_10_i,temp_m1_4_9_r,temp_m1_4_9_i,temp_m1_4_10_r,temp_m1_4_10_i,temp_b1_3_9_r,temp_b1_3_9_i,temp_b1_3_10_r,temp_b1_3_10_i,temp_b1_4_9_r,temp_b1_4_9_i,temp_b1_4_10_r,temp_b1_4_10_i);
MULT MULT22 (clk,in_3_11_r,in_3_11_i,in_3_12_r,in_3_12_i,in_4_11_r,in_4_11_i,in_4_12_r,in_4_12_i,temp_m1_3_11_r,temp_m1_3_11_i,temp_m1_3_12_r,temp_m1_3_12_i,temp_m1_4_11_r,temp_m1_4_11_i,temp_m1_4_12_r,temp_m1_4_12_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly22 (clk,temp_m1_3_11_r,temp_m1_3_11_i,temp_m1_3_12_r,temp_m1_3_12_i,temp_m1_4_11_r,temp_m1_4_11_i,temp_m1_4_12_r,temp_m1_4_12_i,temp_b1_3_11_r,temp_b1_3_11_i,temp_b1_3_12_r,temp_b1_3_12_i,temp_b1_4_11_r,temp_b1_4_11_i,temp_b1_4_12_r,temp_b1_4_12_i);
MULT MULT23 (clk,in_3_13_r,in_3_13_i,in_3_14_r,in_3_14_i,in_4_13_r,in_4_13_i,in_4_14_r,in_4_14_i,temp_m1_3_13_r,temp_m1_3_13_i,temp_m1_3_14_r,temp_m1_3_14_i,temp_m1_4_13_r,temp_m1_4_13_i,temp_m1_4_14_r,temp_m1_4_14_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly23 (clk,temp_m1_3_13_r,temp_m1_3_13_i,temp_m1_3_14_r,temp_m1_3_14_i,temp_m1_4_13_r,temp_m1_4_13_i,temp_m1_4_14_r,temp_m1_4_14_i,temp_b1_3_13_r,temp_b1_3_13_i,temp_b1_3_14_r,temp_b1_3_14_i,temp_b1_4_13_r,temp_b1_4_13_i,temp_b1_4_14_r,temp_b1_4_14_i);
MULT MULT24 (clk,in_3_15_r,in_3_15_i,in_3_16_r,in_3_16_i,in_4_15_r,in_4_15_i,in_4_16_r,in_4_16_i,temp_m1_3_15_r,temp_m1_3_15_i,temp_m1_3_16_r,temp_m1_3_16_i,temp_m1_4_15_r,temp_m1_4_15_i,temp_m1_4_16_r,temp_m1_4_16_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly24 (clk,temp_m1_3_15_r,temp_m1_3_15_i,temp_m1_3_16_r,temp_m1_3_16_i,temp_m1_4_15_r,temp_m1_4_15_i,temp_m1_4_16_r,temp_m1_4_16_i,temp_b1_3_15_r,temp_b1_3_15_i,temp_b1_3_16_r,temp_b1_3_16_i,temp_b1_4_15_r,temp_b1_4_15_i,temp_b1_4_16_r,temp_b1_4_16_i);
MULT MULT25 (clk,in_3_17_r,in_3_17_i,in_3_18_r,in_3_18_i,in_4_17_r,in_4_17_i,in_4_18_r,in_4_18_i,temp_m1_3_17_r,temp_m1_3_17_i,temp_m1_3_18_r,temp_m1_3_18_i,temp_m1_4_17_r,temp_m1_4_17_i,temp_m1_4_18_r,temp_m1_4_18_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly25 (clk,temp_m1_3_17_r,temp_m1_3_17_i,temp_m1_3_18_r,temp_m1_3_18_i,temp_m1_4_17_r,temp_m1_4_17_i,temp_m1_4_18_r,temp_m1_4_18_i,temp_b1_3_17_r,temp_b1_3_17_i,temp_b1_3_18_r,temp_b1_3_18_i,temp_b1_4_17_r,temp_b1_4_17_i,temp_b1_4_18_r,temp_b1_4_18_i);
MULT MULT26 (clk,in_3_19_r,in_3_19_i,in_3_20_r,in_3_20_i,in_4_19_r,in_4_19_i,in_4_20_r,in_4_20_i,temp_m1_3_19_r,temp_m1_3_19_i,temp_m1_3_20_r,temp_m1_3_20_i,temp_m1_4_19_r,temp_m1_4_19_i,temp_m1_4_20_r,temp_m1_4_20_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly26 (clk,temp_m1_3_19_r,temp_m1_3_19_i,temp_m1_3_20_r,temp_m1_3_20_i,temp_m1_4_19_r,temp_m1_4_19_i,temp_m1_4_20_r,temp_m1_4_20_i,temp_b1_3_19_r,temp_b1_3_19_i,temp_b1_3_20_r,temp_b1_3_20_i,temp_b1_4_19_r,temp_b1_4_19_i,temp_b1_4_20_r,temp_b1_4_20_i);
MULT MULT27 (clk,in_3_21_r,in_3_21_i,in_3_22_r,in_3_22_i,in_4_21_r,in_4_21_i,in_4_22_r,in_4_22_i,temp_m1_3_21_r,temp_m1_3_21_i,temp_m1_3_22_r,temp_m1_3_22_i,temp_m1_4_21_r,temp_m1_4_21_i,temp_m1_4_22_r,temp_m1_4_22_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly27 (clk,temp_m1_3_21_r,temp_m1_3_21_i,temp_m1_3_22_r,temp_m1_3_22_i,temp_m1_4_21_r,temp_m1_4_21_i,temp_m1_4_22_r,temp_m1_4_22_i,temp_b1_3_21_r,temp_b1_3_21_i,temp_b1_3_22_r,temp_b1_3_22_i,temp_b1_4_21_r,temp_b1_4_21_i,temp_b1_4_22_r,temp_b1_4_22_i);
MULT MULT28 (clk,in_3_23_r,in_3_23_i,in_3_24_r,in_3_24_i,in_4_23_r,in_4_23_i,in_4_24_r,in_4_24_i,temp_m1_3_23_r,temp_m1_3_23_i,temp_m1_3_24_r,temp_m1_3_24_i,temp_m1_4_23_r,temp_m1_4_23_i,temp_m1_4_24_r,temp_m1_4_24_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly28 (clk,temp_m1_3_23_r,temp_m1_3_23_i,temp_m1_3_24_r,temp_m1_3_24_i,temp_m1_4_23_r,temp_m1_4_23_i,temp_m1_4_24_r,temp_m1_4_24_i,temp_b1_3_23_r,temp_b1_3_23_i,temp_b1_3_24_r,temp_b1_3_24_i,temp_b1_4_23_r,temp_b1_4_23_i,temp_b1_4_24_r,temp_b1_4_24_i);
MULT MULT29 (clk,in_3_25_r,in_3_25_i,in_3_26_r,in_3_26_i,in_4_25_r,in_4_25_i,in_4_26_r,in_4_26_i,temp_m1_3_25_r,temp_m1_3_25_i,temp_m1_3_26_r,temp_m1_3_26_i,temp_m1_4_25_r,temp_m1_4_25_i,temp_m1_4_26_r,temp_m1_4_26_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly29 (clk,temp_m1_3_25_r,temp_m1_3_25_i,temp_m1_3_26_r,temp_m1_3_26_i,temp_m1_4_25_r,temp_m1_4_25_i,temp_m1_4_26_r,temp_m1_4_26_i,temp_b1_3_25_r,temp_b1_3_25_i,temp_b1_3_26_r,temp_b1_3_26_i,temp_b1_4_25_r,temp_b1_4_25_i,temp_b1_4_26_r,temp_b1_4_26_i);
MULT MULT30 (clk,in_3_27_r,in_3_27_i,in_3_28_r,in_3_28_i,in_4_27_r,in_4_27_i,in_4_28_r,in_4_28_i,temp_m1_3_27_r,temp_m1_3_27_i,temp_m1_3_28_r,temp_m1_3_28_i,temp_m1_4_27_r,temp_m1_4_27_i,temp_m1_4_28_r,temp_m1_4_28_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly30 (clk,temp_m1_3_27_r,temp_m1_3_27_i,temp_m1_3_28_r,temp_m1_3_28_i,temp_m1_4_27_r,temp_m1_4_27_i,temp_m1_4_28_r,temp_m1_4_28_i,temp_b1_3_27_r,temp_b1_3_27_i,temp_b1_3_28_r,temp_b1_3_28_i,temp_b1_4_27_r,temp_b1_4_27_i,temp_b1_4_28_r,temp_b1_4_28_i);
MULT MULT31 (clk,in_3_29_r,in_3_29_i,in_3_30_r,in_3_30_i,in_4_29_r,in_4_29_i,in_4_30_r,in_4_30_i,temp_m1_3_29_r,temp_m1_3_29_i,temp_m1_3_30_r,temp_m1_3_30_i,temp_m1_4_29_r,temp_m1_4_29_i,temp_m1_4_30_r,temp_m1_4_30_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly31 (clk,temp_m1_3_29_r,temp_m1_3_29_i,temp_m1_3_30_r,temp_m1_3_30_i,temp_m1_4_29_r,temp_m1_4_29_i,temp_m1_4_30_r,temp_m1_4_30_i,temp_b1_3_29_r,temp_b1_3_29_i,temp_b1_3_30_r,temp_b1_3_30_i,temp_b1_4_29_r,temp_b1_4_29_i,temp_b1_4_30_r,temp_b1_4_30_i);
MULT MULT32 (clk,in_3_31_r,in_3_31_i,in_3_32_r,in_3_32_i,in_4_31_r,in_4_31_i,in_4_32_r,in_4_32_i,temp_m1_3_31_r,temp_m1_3_31_i,temp_m1_3_32_r,temp_m1_3_32_i,temp_m1_4_31_r,temp_m1_4_31_i,temp_m1_4_32_r,temp_m1_4_32_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly32 (clk,temp_m1_3_31_r,temp_m1_3_31_i,temp_m1_3_32_r,temp_m1_3_32_i,temp_m1_4_31_r,temp_m1_4_31_i,temp_m1_4_32_r,temp_m1_4_32_i,temp_b1_3_31_r,temp_b1_3_31_i,temp_b1_3_32_r,temp_b1_3_32_i,temp_b1_4_31_r,temp_b1_4_31_i,temp_b1_4_32_r,temp_b1_4_32_i);
MULT MULT33 (clk,in_5_1_r,in_5_1_i,in_5_2_r,in_5_2_i,in_6_1_r,in_6_1_i,in_6_2_r,in_6_2_i,temp_m1_5_1_r,temp_m1_5_1_i,temp_m1_5_2_r,temp_m1_5_2_i,temp_m1_6_1_r,temp_m1_6_1_i,temp_m1_6_2_r,temp_m1_6_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly33 (clk,temp_m1_5_1_r,temp_m1_5_1_i,temp_m1_5_2_r,temp_m1_5_2_i,temp_m1_6_1_r,temp_m1_6_1_i,temp_m1_6_2_r,temp_m1_6_2_i,temp_b1_5_1_r,temp_b1_5_1_i,temp_b1_5_2_r,temp_b1_5_2_i,temp_b1_6_1_r,temp_b1_6_1_i,temp_b1_6_2_r,temp_b1_6_2_i);
MULT MULT34 (clk,in_5_3_r,in_5_3_i,in_5_4_r,in_5_4_i,in_6_3_r,in_6_3_i,in_6_4_r,in_6_4_i,temp_m1_5_3_r,temp_m1_5_3_i,temp_m1_5_4_r,temp_m1_5_4_i,temp_m1_6_3_r,temp_m1_6_3_i,temp_m1_6_4_r,temp_m1_6_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly34 (clk,temp_m1_5_3_r,temp_m1_5_3_i,temp_m1_5_4_r,temp_m1_5_4_i,temp_m1_6_3_r,temp_m1_6_3_i,temp_m1_6_4_r,temp_m1_6_4_i,temp_b1_5_3_r,temp_b1_5_3_i,temp_b1_5_4_r,temp_b1_5_4_i,temp_b1_6_3_r,temp_b1_6_3_i,temp_b1_6_4_r,temp_b1_6_4_i);
MULT MULT35 (clk,in_5_5_r,in_5_5_i,in_5_6_r,in_5_6_i,in_6_5_r,in_6_5_i,in_6_6_r,in_6_6_i,temp_m1_5_5_r,temp_m1_5_5_i,temp_m1_5_6_r,temp_m1_5_6_i,temp_m1_6_5_r,temp_m1_6_5_i,temp_m1_6_6_r,temp_m1_6_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly35 (clk,temp_m1_5_5_r,temp_m1_5_5_i,temp_m1_5_6_r,temp_m1_5_6_i,temp_m1_6_5_r,temp_m1_6_5_i,temp_m1_6_6_r,temp_m1_6_6_i,temp_b1_5_5_r,temp_b1_5_5_i,temp_b1_5_6_r,temp_b1_5_6_i,temp_b1_6_5_r,temp_b1_6_5_i,temp_b1_6_6_r,temp_b1_6_6_i);
MULT MULT36 (clk,in_5_7_r,in_5_7_i,in_5_8_r,in_5_8_i,in_6_7_r,in_6_7_i,in_6_8_r,in_6_8_i,temp_m1_5_7_r,temp_m1_5_7_i,temp_m1_5_8_r,temp_m1_5_8_i,temp_m1_6_7_r,temp_m1_6_7_i,temp_m1_6_8_r,temp_m1_6_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly36 (clk,temp_m1_5_7_r,temp_m1_5_7_i,temp_m1_5_8_r,temp_m1_5_8_i,temp_m1_6_7_r,temp_m1_6_7_i,temp_m1_6_8_r,temp_m1_6_8_i,temp_b1_5_7_r,temp_b1_5_7_i,temp_b1_5_8_r,temp_b1_5_8_i,temp_b1_6_7_r,temp_b1_6_7_i,temp_b1_6_8_r,temp_b1_6_8_i);
MULT MULT37 (clk,in_5_9_r,in_5_9_i,in_5_10_r,in_5_10_i,in_6_9_r,in_6_9_i,in_6_10_r,in_6_10_i,temp_m1_5_9_r,temp_m1_5_9_i,temp_m1_5_10_r,temp_m1_5_10_i,temp_m1_6_9_r,temp_m1_6_9_i,temp_m1_6_10_r,temp_m1_6_10_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly37 (clk,temp_m1_5_9_r,temp_m1_5_9_i,temp_m1_5_10_r,temp_m1_5_10_i,temp_m1_6_9_r,temp_m1_6_9_i,temp_m1_6_10_r,temp_m1_6_10_i,temp_b1_5_9_r,temp_b1_5_9_i,temp_b1_5_10_r,temp_b1_5_10_i,temp_b1_6_9_r,temp_b1_6_9_i,temp_b1_6_10_r,temp_b1_6_10_i);
MULT MULT38 (clk,in_5_11_r,in_5_11_i,in_5_12_r,in_5_12_i,in_6_11_r,in_6_11_i,in_6_12_r,in_6_12_i,temp_m1_5_11_r,temp_m1_5_11_i,temp_m1_5_12_r,temp_m1_5_12_i,temp_m1_6_11_r,temp_m1_6_11_i,temp_m1_6_12_r,temp_m1_6_12_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly38 (clk,temp_m1_5_11_r,temp_m1_5_11_i,temp_m1_5_12_r,temp_m1_5_12_i,temp_m1_6_11_r,temp_m1_6_11_i,temp_m1_6_12_r,temp_m1_6_12_i,temp_b1_5_11_r,temp_b1_5_11_i,temp_b1_5_12_r,temp_b1_5_12_i,temp_b1_6_11_r,temp_b1_6_11_i,temp_b1_6_12_r,temp_b1_6_12_i);
MULT MULT39 (clk,in_5_13_r,in_5_13_i,in_5_14_r,in_5_14_i,in_6_13_r,in_6_13_i,in_6_14_r,in_6_14_i,temp_m1_5_13_r,temp_m1_5_13_i,temp_m1_5_14_r,temp_m1_5_14_i,temp_m1_6_13_r,temp_m1_6_13_i,temp_m1_6_14_r,temp_m1_6_14_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly39 (clk,temp_m1_5_13_r,temp_m1_5_13_i,temp_m1_5_14_r,temp_m1_5_14_i,temp_m1_6_13_r,temp_m1_6_13_i,temp_m1_6_14_r,temp_m1_6_14_i,temp_b1_5_13_r,temp_b1_5_13_i,temp_b1_5_14_r,temp_b1_5_14_i,temp_b1_6_13_r,temp_b1_6_13_i,temp_b1_6_14_r,temp_b1_6_14_i);
MULT MULT40 (clk,in_5_15_r,in_5_15_i,in_5_16_r,in_5_16_i,in_6_15_r,in_6_15_i,in_6_16_r,in_6_16_i,temp_m1_5_15_r,temp_m1_5_15_i,temp_m1_5_16_r,temp_m1_5_16_i,temp_m1_6_15_r,temp_m1_6_15_i,temp_m1_6_16_r,temp_m1_6_16_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly40 (clk,temp_m1_5_15_r,temp_m1_5_15_i,temp_m1_5_16_r,temp_m1_5_16_i,temp_m1_6_15_r,temp_m1_6_15_i,temp_m1_6_16_r,temp_m1_6_16_i,temp_b1_5_15_r,temp_b1_5_15_i,temp_b1_5_16_r,temp_b1_5_16_i,temp_b1_6_15_r,temp_b1_6_15_i,temp_b1_6_16_r,temp_b1_6_16_i);
MULT MULT41 (clk,in_5_17_r,in_5_17_i,in_5_18_r,in_5_18_i,in_6_17_r,in_6_17_i,in_6_18_r,in_6_18_i,temp_m1_5_17_r,temp_m1_5_17_i,temp_m1_5_18_r,temp_m1_5_18_i,temp_m1_6_17_r,temp_m1_6_17_i,temp_m1_6_18_r,temp_m1_6_18_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly41 (clk,temp_m1_5_17_r,temp_m1_5_17_i,temp_m1_5_18_r,temp_m1_5_18_i,temp_m1_6_17_r,temp_m1_6_17_i,temp_m1_6_18_r,temp_m1_6_18_i,temp_b1_5_17_r,temp_b1_5_17_i,temp_b1_5_18_r,temp_b1_5_18_i,temp_b1_6_17_r,temp_b1_6_17_i,temp_b1_6_18_r,temp_b1_6_18_i);
MULT MULT42 (clk,in_5_19_r,in_5_19_i,in_5_20_r,in_5_20_i,in_6_19_r,in_6_19_i,in_6_20_r,in_6_20_i,temp_m1_5_19_r,temp_m1_5_19_i,temp_m1_5_20_r,temp_m1_5_20_i,temp_m1_6_19_r,temp_m1_6_19_i,temp_m1_6_20_r,temp_m1_6_20_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly42 (clk,temp_m1_5_19_r,temp_m1_5_19_i,temp_m1_5_20_r,temp_m1_5_20_i,temp_m1_6_19_r,temp_m1_6_19_i,temp_m1_6_20_r,temp_m1_6_20_i,temp_b1_5_19_r,temp_b1_5_19_i,temp_b1_5_20_r,temp_b1_5_20_i,temp_b1_6_19_r,temp_b1_6_19_i,temp_b1_6_20_r,temp_b1_6_20_i);
MULT MULT43 (clk,in_5_21_r,in_5_21_i,in_5_22_r,in_5_22_i,in_6_21_r,in_6_21_i,in_6_22_r,in_6_22_i,temp_m1_5_21_r,temp_m1_5_21_i,temp_m1_5_22_r,temp_m1_5_22_i,temp_m1_6_21_r,temp_m1_6_21_i,temp_m1_6_22_r,temp_m1_6_22_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly43 (clk,temp_m1_5_21_r,temp_m1_5_21_i,temp_m1_5_22_r,temp_m1_5_22_i,temp_m1_6_21_r,temp_m1_6_21_i,temp_m1_6_22_r,temp_m1_6_22_i,temp_b1_5_21_r,temp_b1_5_21_i,temp_b1_5_22_r,temp_b1_5_22_i,temp_b1_6_21_r,temp_b1_6_21_i,temp_b1_6_22_r,temp_b1_6_22_i);
MULT MULT44 (clk,in_5_23_r,in_5_23_i,in_5_24_r,in_5_24_i,in_6_23_r,in_6_23_i,in_6_24_r,in_6_24_i,temp_m1_5_23_r,temp_m1_5_23_i,temp_m1_5_24_r,temp_m1_5_24_i,temp_m1_6_23_r,temp_m1_6_23_i,temp_m1_6_24_r,temp_m1_6_24_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly44 (clk,temp_m1_5_23_r,temp_m1_5_23_i,temp_m1_5_24_r,temp_m1_5_24_i,temp_m1_6_23_r,temp_m1_6_23_i,temp_m1_6_24_r,temp_m1_6_24_i,temp_b1_5_23_r,temp_b1_5_23_i,temp_b1_5_24_r,temp_b1_5_24_i,temp_b1_6_23_r,temp_b1_6_23_i,temp_b1_6_24_r,temp_b1_6_24_i);
MULT MULT45 (clk,in_5_25_r,in_5_25_i,in_5_26_r,in_5_26_i,in_6_25_r,in_6_25_i,in_6_26_r,in_6_26_i,temp_m1_5_25_r,temp_m1_5_25_i,temp_m1_5_26_r,temp_m1_5_26_i,temp_m1_6_25_r,temp_m1_6_25_i,temp_m1_6_26_r,temp_m1_6_26_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly45 (clk,temp_m1_5_25_r,temp_m1_5_25_i,temp_m1_5_26_r,temp_m1_5_26_i,temp_m1_6_25_r,temp_m1_6_25_i,temp_m1_6_26_r,temp_m1_6_26_i,temp_b1_5_25_r,temp_b1_5_25_i,temp_b1_5_26_r,temp_b1_5_26_i,temp_b1_6_25_r,temp_b1_6_25_i,temp_b1_6_26_r,temp_b1_6_26_i);
MULT MULT46 (clk,in_5_27_r,in_5_27_i,in_5_28_r,in_5_28_i,in_6_27_r,in_6_27_i,in_6_28_r,in_6_28_i,temp_m1_5_27_r,temp_m1_5_27_i,temp_m1_5_28_r,temp_m1_5_28_i,temp_m1_6_27_r,temp_m1_6_27_i,temp_m1_6_28_r,temp_m1_6_28_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly46 (clk,temp_m1_5_27_r,temp_m1_5_27_i,temp_m1_5_28_r,temp_m1_5_28_i,temp_m1_6_27_r,temp_m1_6_27_i,temp_m1_6_28_r,temp_m1_6_28_i,temp_b1_5_27_r,temp_b1_5_27_i,temp_b1_5_28_r,temp_b1_5_28_i,temp_b1_6_27_r,temp_b1_6_27_i,temp_b1_6_28_r,temp_b1_6_28_i);
MULT MULT47 (clk,in_5_29_r,in_5_29_i,in_5_30_r,in_5_30_i,in_6_29_r,in_6_29_i,in_6_30_r,in_6_30_i,temp_m1_5_29_r,temp_m1_5_29_i,temp_m1_5_30_r,temp_m1_5_30_i,temp_m1_6_29_r,temp_m1_6_29_i,temp_m1_6_30_r,temp_m1_6_30_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly47 (clk,temp_m1_5_29_r,temp_m1_5_29_i,temp_m1_5_30_r,temp_m1_5_30_i,temp_m1_6_29_r,temp_m1_6_29_i,temp_m1_6_30_r,temp_m1_6_30_i,temp_b1_5_29_r,temp_b1_5_29_i,temp_b1_5_30_r,temp_b1_5_30_i,temp_b1_6_29_r,temp_b1_6_29_i,temp_b1_6_30_r,temp_b1_6_30_i);
MULT MULT48 (clk,in_5_31_r,in_5_31_i,in_5_32_r,in_5_32_i,in_6_31_r,in_6_31_i,in_6_32_r,in_6_32_i,temp_m1_5_31_r,temp_m1_5_31_i,temp_m1_5_32_r,temp_m1_5_32_i,temp_m1_6_31_r,temp_m1_6_31_i,temp_m1_6_32_r,temp_m1_6_32_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly48 (clk,temp_m1_5_31_r,temp_m1_5_31_i,temp_m1_5_32_r,temp_m1_5_32_i,temp_m1_6_31_r,temp_m1_6_31_i,temp_m1_6_32_r,temp_m1_6_32_i,temp_b1_5_31_r,temp_b1_5_31_i,temp_b1_5_32_r,temp_b1_5_32_i,temp_b1_6_31_r,temp_b1_6_31_i,temp_b1_6_32_r,temp_b1_6_32_i);
MULT MULT49 (clk,in_7_1_r,in_7_1_i,in_7_2_r,in_7_2_i,in_8_1_r,in_8_1_i,in_8_2_r,in_8_2_i,temp_m1_7_1_r,temp_m1_7_1_i,temp_m1_7_2_r,temp_m1_7_2_i,temp_m1_8_1_r,temp_m1_8_1_i,temp_m1_8_2_r,temp_m1_8_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly49 (clk,temp_m1_7_1_r,temp_m1_7_1_i,temp_m1_7_2_r,temp_m1_7_2_i,temp_m1_8_1_r,temp_m1_8_1_i,temp_m1_8_2_r,temp_m1_8_2_i,temp_b1_7_1_r,temp_b1_7_1_i,temp_b1_7_2_r,temp_b1_7_2_i,temp_b1_8_1_r,temp_b1_8_1_i,temp_b1_8_2_r,temp_b1_8_2_i);
MULT MULT50 (clk,in_7_3_r,in_7_3_i,in_7_4_r,in_7_4_i,in_8_3_r,in_8_3_i,in_8_4_r,in_8_4_i,temp_m1_7_3_r,temp_m1_7_3_i,temp_m1_7_4_r,temp_m1_7_4_i,temp_m1_8_3_r,temp_m1_8_3_i,temp_m1_8_4_r,temp_m1_8_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly50 (clk,temp_m1_7_3_r,temp_m1_7_3_i,temp_m1_7_4_r,temp_m1_7_4_i,temp_m1_8_3_r,temp_m1_8_3_i,temp_m1_8_4_r,temp_m1_8_4_i,temp_b1_7_3_r,temp_b1_7_3_i,temp_b1_7_4_r,temp_b1_7_4_i,temp_b1_8_3_r,temp_b1_8_3_i,temp_b1_8_4_r,temp_b1_8_4_i);
MULT MULT51 (clk,in_7_5_r,in_7_5_i,in_7_6_r,in_7_6_i,in_8_5_r,in_8_5_i,in_8_6_r,in_8_6_i,temp_m1_7_5_r,temp_m1_7_5_i,temp_m1_7_6_r,temp_m1_7_6_i,temp_m1_8_5_r,temp_m1_8_5_i,temp_m1_8_6_r,temp_m1_8_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly51 (clk,temp_m1_7_5_r,temp_m1_7_5_i,temp_m1_7_6_r,temp_m1_7_6_i,temp_m1_8_5_r,temp_m1_8_5_i,temp_m1_8_6_r,temp_m1_8_6_i,temp_b1_7_5_r,temp_b1_7_5_i,temp_b1_7_6_r,temp_b1_7_6_i,temp_b1_8_5_r,temp_b1_8_5_i,temp_b1_8_6_r,temp_b1_8_6_i);
MULT MULT52 (clk,in_7_7_r,in_7_7_i,in_7_8_r,in_7_8_i,in_8_7_r,in_8_7_i,in_8_8_r,in_8_8_i,temp_m1_7_7_r,temp_m1_7_7_i,temp_m1_7_8_r,temp_m1_7_8_i,temp_m1_8_7_r,temp_m1_8_7_i,temp_m1_8_8_r,temp_m1_8_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly52 (clk,temp_m1_7_7_r,temp_m1_7_7_i,temp_m1_7_8_r,temp_m1_7_8_i,temp_m1_8_7_r,temp_m1_8_7_i,temp_m1_8_8_r,temp_m1_8_8_i,temp_b1_7_7_r,temp_b1_7_7_i,temp_b1_7_8_r,temp_b1_7_8_i,temp_b1_8_7_r,temp_b1_8_7_i,temp_b1_8_8_r,temp_b1_8_8_i);
MULT MULT53 (clk,in_7_9_r,in_7_9_i,in_7_10_r,in_7_10_i,in_8_9_r,in_8_9_i,in_8_10_r,in_8_10_i,temp_m1_7_9_r,temp_m1_7_9_i,temp_m1_7_10_r,temp_m1_7_10_i,temp_m1_8_9_r,temp_m1_8_9_i,temp_m1_8_10_r,temp_m1_8_10_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly53 (clk,temp_m1_7_9_r,temp_m1_7_9_i,temp_m1_7_10_r,temp_m1_7_10_i,temp_m1_8_9_r,temp_m1_8_9_i,temp_m1_8_10_r,temp_m1_8_10_i,temp_b1_7_9_r,temp_b1_7_9_i,temp_b1_7_10_r,temp_b1_7_10_i,temp_b1_8_9_r,temp_b1_8_9_i,temp_b1_8_10_r,temp_b1_8_10_i);
MULT MULT54 (clk,in_7_11_r,in_7_11_i,in_7_12_r,in_7_12_i,in_8_11_r,in_8_11_i,in_8_12_r,in_8_12_i,temp_m1_7_11_r,temp_m1_7_11_i,temp_m1_7_12_r,temp_m1_7_12_i,temp_m1_8_11_r,temp_m1_8_11_i,temp_m1_8_12_r,temp_m1_8_12_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly54 (clk,temp_m1_7_11_r,temp_m1_7_11_i,temp_m1_7_12_r,temp_m1_7_12_i,temp_m1_8_11_r,temp_m1_8_11_i,temp_m1_8_12_r,temp_m1_8_12_i,temp_b1_7_11_r,temp_b1_7_11_i,temp_b1_7_12_r,temp_b1_7_12_i,temp_b1_8_11_r,temp_b1_8_11_i,temp_b1_8_12_r,temp_b1_8_12_i);
MULT MULT55 (clk,in_7_13_r,in_7_13_i,in_7_14_r,in_7_14_i,in_8_13_r,in_8_13_i,in_8_14_r,in_8_14_i,temp_m1_7_13_r,temp_m1_7_13_i,temp_m1_7_14_r,temp_m1_7_14_i,temp_m1_8_13_r,temp_m1_8_13_i,temp_m1_8_14_r,temp_m1_8_14_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly55 (clk,temp_m1_7_13_r,temp_m1_7_13_i,temp_m1_7_14_r,temp_m1_7_14_i,temp_m1_8_13_r,temp_m1_8_13_i,temp_m1_8_14_r,temp_m1_8_14_i,temp_b1_7_13_r,temp_b1_7_13_i,temp_b1_7_14_r,temp_b1_7_14_i,temp_b1_8_13_r,temp_b1_8_13_i,temp_b1_8_14_r,temp_b1_8_14_i);
MULT MULT56 (clk,in_7_15_r,in_7_15_i,in_7_16_r,in_7_16_i,in_8_15_r,in_8_15_i,in_8_16_r,in_8_16_i,temp_m1_7_15_r,temp_m1_7_15_i,temp_m1_7_16_r,temp_m1_7_16_i,temp_m1_8_15_r,temp_m1_8_15_i,temp_m1_8_16_r,temp_m1_8_16_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly56 (clk,temp_m1_7_15_r,temp_m1_7_15_i,temp_m1_7_16_r,temp_m1_7_16_i,temp_m1_8_15_r,temp_m1_8_15_i,temp_m1_8_16_r,temp_m1_8_16_i,temp_b1_7_15_r,temp_b1_7_15_i,temp_b1_7_16_r,temp_b1_7_16_i,temp_b1_8_15_r,temp_b1_8_15_i,temp_b1_8_16_r,temp_b1_8_16_i);
MULT MULT57 (clk,in_7_17_r,in_7_17_i,in_7_18_r,in_7_18_i,in_8_17_r,in_8_17_i,in_8_18_r,in_8_18_i,temp_m1_7_17_r,temp_m1_7_17_i,temp_m1_7_18_r,temp_m1_7_18_i,temp_m1_8_17_r,temp_m1_8_17_i,temp_m1_8_18_r,temp_m1_8_18_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly57 (clk,temp_m1_7_17_r,temp_m1_7_17_i,temp_m1_7_18_r,temp_m1_7_18_i,temp_m1_8_17_r,temp_m1_8_17_i,temp_m1_8_18_r,temp_m1_8_18_i,temp_b1_7_17_r,temp_b1_7_17_i,temp_b1_7_18_r,temp_b1_7_18_i,temp_b1_8_17_r,temp_b1_8_17_i,temp_b1_8_18_r,temp_b1_8_18_i);
MULT MULT58 (clk,in_7_19_r,in_7_19_i,in_7_20_r,in_7_20_i,in_8_19_r,in_8_19_i,in_8_20_r,in_8_20_i,temp_m1_7_19_r,temp_m1_7_19_i,temp_m1_7_20_r,temp_m1_7_20_i,temp_m1_8_19_r,temp_m1_8_19_i,temp_m1_8_20_r,temp_m1_8_20_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly58 (clk,temp_m1_7_19_r,temp_m1_7_19_i,temp_m1_7_20_r,temp_m1_7_20_i,temp_m1_8_19_r,temp_m1_8_19_i,temp_m1_8_20_r,temp_m1_8_20_i,temp_b1_7_19_r,temp_b1_7_19_i,temp_b1_7_20_r,temp_b1_7_20_i,temp_b1_8_19_r,temp_b1_8_19_i,temp_b1_8_20_r,temp_b1_8_20_i);
MULT MULT59 (clk,in_7_21_r,in_7_21_i,in_7_22_r,in_7_22_i,in_8_21_r,in_8_21_i,in_8_22_r,in_8_22_i,temp_m1_7_21_r,temp_m1_7_21_i,temp_m1_7_22_r,temp_m1_7_22_i,temp_m1_8_21_r,temp_m1_8_21_i,temp_m1_8_22_r,temp_m1_8_22_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly59 (clk,temp_m1_7_21_r,temp_m1_7_21_i,temp_m1_7_22_r,temp_m1_7_22_i,temp_m1_8_21_r,temp_m1_8_21_i,temp_m1_8_22_r,temp_m1_8_22_i,temp_b1_7_21_r,temp_b1_7_21_i,temp_b1_7_22_r,temp_b1_7_22_i,temp_b1_8_21_r,temp_b1_8_21_i,temp_b1_8_22_r,temp_b1_8_22_i);
MULT MULT60 (clk,in_7_23_r,in_7_23_i,in_7_24_r,in_7_24_i,in_8_23_r,in_8_23_i,in_8_24_r,in_8_24_i,temp_m1_7_23_r,temp_m1_7_23_i,temp_m1_7_24_r,temp_m1_7_24_i,temp_m1_8_23_r,temp_m1_8_23_i,temp_m1_8_24_r,temp_m1_8_24_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly60 (clk,temp_m1_7_23_r,temp_m1_7_23_i,temp_m1_7_24_r,temp_m1_7_24_i,temp_m1_8_23_r,temp_m1_8_23_i,temp_m1_8_24_r,temp_m1_8_24_i,temp_b1_7_23_r,temp_b1_7_23_i,temp_b1_7_24_r,temp_b1_7_24_i,temp_b1_8_23_r,temp_b1_8_23_i,temp_b1_8_24_r,temp_b1_8_24_i);
MULT MULT61 (clk,in_7_25_r,in_7_25_i,in_7_26_r,in_7_26_i,in_8_25_r,in_8_25_i,in_8_26_r,in_8_26_i,temp_m1_7_25_r,temp_m1_7_25_i,temp_m1_7_26_r,temp_m1_7_26_i,temp_m1_8_25_r,temp_m1_8_25_i,temp_m1_8_26_r,temp_m1_8_26_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly61 (clk,temp_m1_7_25_r,temp_m1_7_25_i,temp_m1_7_26_r,temp_m1_7_26_i,temp_m1_8_25_r,temp_m1_8_25_i,temp_m1_8_26_r,temp_m1_8_26_i,temp_b1_7_25_r,temp_b1_7_25_i,temp_b1_7_26_r,temp_b1_7_26_i,temp_b1_8_25_r,temp_b1_8_25_i,temp_b1_8_26_r,temp_b1_8_26_i);
MULT MULT62 (clk,in_7_27_r,in_7_27_i,in_7_28_r,in_7_28_i,in_8_27_r,in_8_27_i,in_8_28_r,in_8_28_i,temp_m1_7_27_r,temp_m1_7_27_i,temp_m1_7_28_r,temp_m1_7_28_i,temp_m1_8_27_r,temp_m1_8_27_i,temp_m1_8_28_r,temp_m1_8_28_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly62 (clk,temp_m1_7_27_r,temp_m1_7_27_i,temp_m1_7_28_r,temp_m1_7_28_i,temp_m1_8_27_r,temp_m1_8_27_i,temp_m1_8_28_r,temp_m1_8_28_i,temp_b1_7_27_r,temp_b1_7_27_i,temp_b1_7_28_r,temp_b1_7_28_i,temp_b1_8_27_r,temp_b1_8_27_i,temp_b1_8_28_r,temp_b1_8_28_i);
MULT MULT63 (clk,in_7_29_r,in_7_29_i,in_7_30_r,in_7_30_i,in_8_29_r,in_8_29_i,in_8_30_r,in_8_30_i,temp_m1_7_29_r,temp_m1_7_29_i,temp_m1_7_30_r,temp_m1_7_30_i,temp_m1_8_29_r,temp_m1_8_29_i,temp_m1_8_30_r,temp_m1_8_30_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly63 (clk,temp_m1_7_29_r,temp_m1_7_29_i,temp_m1_7_30_r,temp_m1_7_30_i,temp_m1_8_29_r,temp_m1_8_29_i,temp_m1_8_30_r,temp_m1_8_30_i,temp_b1_7_29_r,temp_b1_7_29_i,temp_b1_7_30_r,temp_b1_7_30_i,temp_b1_8_29_r,temp_b1_8_29_i,temp_b1_8_30_r,temp_b1_8_30_i);
MULT MULT64 (clk,in_7_31_r,in_7_31_i,in_7_32_r,in_7_32_i,in_8_31_r,in_8_31_i,in_8_32_r,in_8_32_i,temp_m1_7_31_r,temp_m1_7_31_i,temp_m1_7_32_r,temp_m1_7_32_i,temp_m1_8_31_r,temp_m1_8_31_i,temp_m1_8_32_r,temp_m1_8_32_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly64 (clk,temp_m1_7_31_r,temp_m1_7_31_i,temp_m1_7_32_r,temp_m1_7_32_i,temp_m1_8_31_r,temp_m1_8_31_i,temp_m1_8_32_r,temp_m1_8_32_i,temp_b1_7_31_r,temp_b1_7_31_i,temp_b1_7_32_r,temp_b1_7_32_i,temp_b1_8_31_r,temp_b1_8_31_i,temp_b1_8_32_r,temp_b1_8_32_i);
MULT MULT65 (clk,in_9_1_r,in_9_1_i,in_9_2_r,in_9_2_i,in_10_1_r,in_10_1_i,in_10_2_r,in_10_2_i,temp_m1_9_1_r,temp_m1_9_1_i,temp_m1_9_2_r,temp_m1_9_2_i,temp_m1_10_1_r,temp_m1_10_1_i,temp_m1_10_2_r,temp_m1_10_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly65 (clk,temp_m1_9_1_r,temp_m1_9_1_i,temp_m1_9_2_r,temp_m1_9_2_i,temp_m1_10_1_r,temp_m1_10_1_i,temp_m1_10_2_r,temp_m1_10_2_i,temp_b1_9_1_r,temp_b1_9_1_i,temp_b1_9_2_r,temp_b1_9_2_i,temp_b1_10_1_r,temp_b1_10_1_i,temp_b1_10_2_r,temp_b1_10_2_i);
MULT MULT66 (clk,in_9_3_r,in_9_3_i,in_9_4_r,in_9_4_i,in_10_3_r,in_10_3_i,in_10_4_r,in_10_4_i,temp_m1_9_3_r,temp_m1_9_3_i,temp_m1_9_4_r,temp_m1_9_4_i,temp_m1_10_3_r,temp_m1_10_3_i,temp_m1_10_4_r,temp_m1_10_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly66 (clk,temp_m1_9_3_r,temp_m1_9_3_i,temp_m1_9_4_r,temp_m1_9_4_i,temp_m1_10_3_r,temp_m1_10_3_i,temp_m1_10_4_r,temp_m1_10_4_i,temp_b1_9_3_r,temp_b1_9_3_i,temp_b1_9_4_r,temp_b1_9_4_i,temp_b1_10_3_r,temp_b1_10_3_i,temp_b1_10_4_r,temp_b1_10_4_i);
MULT MULT67 (clk,in_9_5_r,in_9_5_i,in_9_6_r,in_9_6_i,in_10_5_r,in_10_5_i,in_10_6_r,in_10_6_i,temp_m1_9_5_r,temp_m1_9_5_i,temp_m1_9_6_r,temp_m1_9_6_i,temp_m1_10_5_r,temp_m1_10_5_i,temp_m1_10_6_r,temp_m1_10_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly67 (clk,temp_m1_9_5_r,temp_m1_9_5_i,temp_m1_9_6_r,temp_m1_9_6_i,temp_m1_10_5_r,temp_m1_10_5_i,temp_m1_10_6_r,temp_m1_10_6_i,temp_b1_9_5_r,temp_b1_9_5_i,temp_b1_9_6_r,temp_b1_9_6_i,temp_b1_10_5_r,temp_b1_10_5_i,temp_b1_10_6_r,temp_b1_10_6_i);
MULT MULT68 (clk,in_9_7_r,in_9_7_i,in_9_8_r,in_9_8_i,in_10_7_r,in_10_7_i,in_10_8_r,in_10_8_i,temp_m1_9_7_r,temp_m1_9_7_i,temp_m1_9_8_r,temp_m1_9_8_i,temp_m1_10_7_r,temp_m1_10_7_i,temp_m1_10_8_r,temp_m1_10_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly68 (clk,temp_m1_9_7_r,temp_m1_9_7_i,temp_m1_9_8_r,temp_m1_9_8_i,temp_m1_10_7_r,temp_m1_10_7_i,temp_m1_10_8_r,temp_m1_10_8_i,temp_b1_9_7_r,temp_b1_9_7_i,temp_b1_9_8_r,temp_b1_9_8_i,temp_b1_10_7_r,temp_b1_10_7_i,temp_b1_10_8_r,temp_b1_10_8_i);
MULT MULT69 (clk,in_9_9_r,in_9_9_i,in_9_10_r,in_9_10_i,in_10_9_r,in_10_9_i,in_10_10_r,in_10_10_i,temp_m1_9_9_r,temp_m1_9_9_i,temp_m1_9_10_r,temp_m1_9_10_i,temp_m1_10_9_r,temp_m1_10_9_i,temp_m1_10_10_r,temp_m1_10_10_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly69 (clk,temp_m1_9_9_r,temp_m1_9_9_i,temp_m1_9_10_r,temp_m1_9_10_i,temp_m1_10_9_r,temp_m1_10_9_i,temp_m1_10_10_r,temp_m1_10_10_i,temp_b1_9_9_r,temp_b1_9_9_i,temp_b1_9_10_r,temp_b1_9_10_i,temp_b1_10_9_r,temp_b1_10_9_i,temp_b1_10_10_r,temp_b1_10_10_i);
MULT MULT70 (clk,in_9_11_r,in_9_11_i,in_9_12_r,in_9_12_i,in_10_11_r,in_10_11_i,in_10_12_r,in_10_12_i,temp_m1_9_11_r,temp_m1_9_11_i,temp_m1_9_12_r,temp_m1_9_12_i,temp_m1_10_11_r,temp_m1_10_11_i,temp_m1_10_12_r,temp_m1_10_12_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly70 (clk,temp_m1_9_11_r,temp_m1_9_11_i,temp_m1_9_12_r,temp_m1_9_12_i,temp_m1_10_11_r,temp_m1_10_11_i,temp_m1_10_12_r,temp_m1_10_12_i,temp_b1_9_11_r,temp_b1_9_11_i,temp_b1_9_12_r,temp_b1_9_12_i,temp_b1_10_11_r,temp_b1_10_11_i,temp_b1_10_12_r,temp_b1_10_12_i);
MULT MULT71 (clk,in_9_13_r,in_9_13_i,in_9_14_r,in_9_14_i,in_10_13_r,in_10_13_i,in_10_14_r,in_10_14_i,temp_m1_9_13_r,temp_m1_9_13_i,temp_m1_9_14_r,temp_m1_9_14_i,temp_m1_10_13_r,temp_m1_10_13_i,temp_m1_10_14_r,temp_m1_10_14_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly71 (clk,temp_m1_9_13_r,temp_m1_9_13_i,temp_m1_9_14_r,temp_m1_9_14_i,temp_m1_10_13_r,temp_m1_10_13_i,temp_m1_10_14_r,temp_m1_10_14_i,temp_b1_9_13_r,temp_b1_9_13_i,temp_b1_9_14_r,temp_b1_9_14_i,temp_b1_10_13_r,temp_b1_10_13_i,temp_b1_10_14_r,temp_b1_10_14_i);
MULT MULT72 (clk,in_9_15_r,in_9_15_i,in_9_16_r,in_9_16_i,in_10_15_r,in_10_15_i,in_10_16_r,in_10_16_i,temp_m1_9_15_r,temp_m1_9_15_i,temp_m1_9_16_r,temp_m1_9_16_i,temp_m1_10_15_r,temp_m1_10_15_i,temp_m1_10_16_r,temp_m1_10_16_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly72 (clk,temp_m1_9_15_r,temp_m1_9_15_i,temp_m1_9_16_r,temp_m1_9_16_i,temp_m1_10_15_r,temp_m1_10_15_i,temp_m1_10_16_r,temp_m1_10_16_i,temp_b1_9_15_r,temp_b1_9_15_i,temp_b1_9_16_r,temp_b1_9_16_i,temp_b1_10_15_r,temp_b1_10_15_i,temp_b1_10_16_r,temp_b1_10_16_i);
MULT MULT73 (clk,in_9_17_r,in_9_17_i,in_9_18_r,in_9_18_i,in_10_17_r,in_10_17_i,in_10_18_r,in_10_18_i,temp_m1_9_17_r,temp_m1_9_17_i,temp_m1_9_18_r,temp_m1_9_18_i,temp_m1_10_17_r,temp_m1_10_17_i,temp_m1_10_18_r,temp_m1_10_18_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly73 (clk,temp_m1_9_17_r,temp_m1_9_17_i,temp_m1_9_18_r,temp_m1_9_18_i,temp_m1_10_17_r,temp_m1_10_17_i,temp_m1_10_18_r,temp_m1_10_18_i,temp_b1_9_17_r,temp_b1_9_17_i,temp_b1_9_18_r,temp_b1_9_18_i,temp_b1_10_17_r,temp_b1_10_17_i,temp_b1_10_18_r,temp_b1_10_18_i);
MULT MULT74 (clk,in_9_19_r,in_9_19_i,in_9_20_r,in_9_20_i,in_10_19_r,in_10_19_i,in_10_20_r,in_10_20_i,temp_m1_9_19_r,temp_m1_9_19_i,temp_m1_9_20_r,temp_m1_9_20_i,temp_m1_10_19_r,temp_m1_10_19_i,temp_m1_10_20_r,temp_m1_10_20_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly74 (clk,temp_m1_9_19_r,temp_m1_9_19_i,temp_m1_9_20_r,temp_m1_9_20_i,temp_m1_10_19_r,temp_m1_10_19_i,temp_m1_10_20_r,temp_m1_10_20_i,temp_b1_9_19_r,temp_b1_9_19_i,temp_b1_9_20_r,temp_b1_9_20_i,temp_b1_10_19_r,temp_b1_10_19_i,temp_b1_10_20_r,temp_b1_10_20_i);
MULT MULT75 (clk,in_9_21_r,in_9_21_i,in_9_22_r,in_9_22_i,in_10_21_r,in_10_21_i,in_10_22_r,in_10_22_i,temp_m1_9_21_r,temp_m1_9_21_i,temp_m1_9_22_r,temp_m1_9_22_i,temp_m1_10_21_r,temp_m1_10_21_i,temp_m1_10_22_r,temp_m1_10_22_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly75 (clk,temp_m1_9_21_r,temp_m1_9_21_i,temp_m1_9_22_r,temp_m1_9_22_i,temp_m1_10_21_r,temp_m1_10_21_i,temp_m1_10_22_r,temp_m1_10_22_i,temp_b1_9_21_r,temp_b1_9_21_i,temp_b1_9_22_r,temp_b1_9_22_i,temp_b1_10_21_r,temp_b1_10_21_i,temp_b1_10_22_r,temp_b1_10_22_i);
MULT MULT76 (clk,in_9_23_r,in_9_23_i,in_9_24_r,in_9_24_i,in_10_23_r,in_10_23_i,in_10_24_r,in_10_24_i,temp_m1_9_23_r,temp_m1_9_23_i,temp_m1_9_24_r,temp_m1_9_24_i,temp_m1_10_23_r,temp_m1_10_23_i,temp_m1_10_24_r,temp_m1_10_24_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly76 (clk,temp_m1_9_23_r,temp_m1_9_23_i,temp_m1_9_24_r,temp_m1_9_24_i,temp_m1_10_23_r,temp_m1_10_23_i,temp_m1_10_24_r,temp_m1_10_24_i,temp_b1_9_23_r,temp_b1_9_23_i,temp_b1_9_24_r,temp_b1_9_24_i,temp_b1_10_23_r,temp_b1_10_23_i,temp_b1_10_24_r,temp_b1_10_24_i);
MULT MULT77 (clk,in_9_25_r,in_9_25_i,in_9_26_r,in_9_26_i,in_10_25_r,in_10_25_i,in_10_26_r,in_10_26_i,temp_m1_9_25_r,temp_m1_9_25_i,temp_m1_9_26_r,temp_m1_9_26_i,temp_m1_10_25_r,temp_m1_10_25_i,temp_m1_10_26_r,temp_m1_10_26_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly77 (clk,temp_m1_9_25_r,temp_m1_9_25_i,temp_m1_9_26_r,temp_m1_9_26_i,temp_m1_10_25_r,temp_m1_10_25_i,temp_m1_10_26_r,temp_m1_10_26_i,temp_b1_9_25_r,temp_b1_9_25_i,temp_b1_9_26_r,temp_b1_9_26_i,temp_b1_10_25_r,temp_b1_10_25_i,temp_b1_10_26_r,temp_b1_10_26_i);
MULT MULT78 (clk,in_9_27_r,in_9_27_i,in_9_28_r,in_9_28_i,in_10_27_r,in_10_27_i,in_10_28_r,in_10_28_i,temp_m1_9_27_r,temp_m1_9_27_i,temp_m1_9_28_r,temp_m1_9_28_i,temp_m1_10_27_r,temp_m1_10_27_i,temp_m1_10_28_r,temp_m1_10_28_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly78 (clk,temp_m1_9_27_r,temp_m1_9_27_i,temp_m1_9_28_r,temp_m1_9_28_i,temp_m1_10_27_r,temp_m1_10_27_i,temp_m1_10_28_r,temp_m1_10_28_i,temp_b1_9_27_r,temp_b1_9_27_i,temp_b1_9_28_r,temp_b1_9_28_i,temp_b1_10_27_r,temp_b1_10_27_i,temp_b1_10_28_r,temp_b1_10_28_i);
MULT MULT79 (clk,in_9_29_r,in_9_29_i,in_9_30_r,in_9_30_i,in_10_29_r,in_10_29_i,in_10_30_r,in_10_30_i,temp_m1_9_29_r,temp_m1_9_29_i,temp_m1_9_30_r,temp_m1_9_30_i,temp_m1_10_29_r,temp_m1_10_29_i,temp_m1_10_30_r,temp_m1_10_30_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly79 (clk,temp_m1_9_29_r,temp_m1_9_29_i,temp_m1_9_30_r,temp_m1_9_30_i,temp_m1_10_29_r,temp_m1_10_29_i,temp_m1_10_30_r,temp_m1_10_30_i,temp_b1_9_29_r,temp_b1_9_29_i,temp_b1_9_30_r,temp_b1_9_30_i,temp_b1_10_29_r,temp_b1_10_29_i,temp_b1_10_30_r,temp_b1_10_30_i);
MULT MULT80 (clk,in_9_31_r,in_9_31_i,in_9_32_r,in_9_32_i,in_10_31_r,in_10_31_i,in_10_32_r,in_10_32_i,temp_m1_9_31_r,temp_m1_9_31_i,temp_m1_9_32_r,temp_m1_9_32_i,temp_m1_10_31_r,temp_m1_10_31_i,temp_m1_10_32_r,temp_m1_10_32_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly80 (clk,temp_m1_9_31_r,temp_m1_9_31_i,temp_m1_9_32_r,temp_m1_9_32_i,temp_m1_10_31_r,temp_m1_10_31_i,temp_m1_10_32_r,temp_m1_10_32_i,temp_b1_9_31_r,temp_b1_9_31_i,temp_b1_9_32_r,temp_b1_9_32_i,temp_b1_10_31_r,temp_b1_10_31_i,temp_b1_10_32_r,temp_b1_10_32_i);
MULT MULT81 (clk,in_11_1_r,in_11_1_i,in_11_2_r,in_11_2_i,in_12_1_r,in_12_1_i,in_12_2_r,in_12_2_i,temp_m1_11_1_r,temp_m1_11_1_i,temp_m1_11_2_r,temp_m1_11_2_i,temp_m1_12_1_r,temp_m1_12_1_i,temp_m1_12_2_r,temp_m1_12_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly81 (clk,temp_m1_11_1_r,temp_m1_11_1_i,temp_m1_11_2_r,temp_m1_11_2_i,temp_m1_12_1_r,temp_m1_12_1_i,temp_m1_12_2_r,temp_m1_12_2_i,temp_b1_11_1_r,temp_b1_11_1_i,temp_b1_11_2_r,temp_b1_11_2_i,temp_b1_12_1_r,temp_b1_12_1_i,temp_b1_12_2_r,temp_b1_12_2_i);
MULT MULT82 (clk,in_11_3_r,in_11_3_i,in_11_4_r,in_11_4_i,in_12_3_r,in_12_3_i,in_12_4_r,in_12_4_i,temp_m1_11_3_r,temp_m1_11_3_i,temp_m1_11_4_r,temp_m1_11_4_i,temp_m1_12_3_r,temp_m1_12_3_i,temp_m1_12_4_r,temp_m1_12_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly82 (clk,temp_m1_11_3_r,temp_m1_11_3_i,temp_m1_11_4_r,temp_m1_11_4_i,temp_m1_12_3_r,temp_m1_12_3_i,temp_m1_12_4_r,temp_m1_12_4_i,temp_b1_11_3_r,temp_b1_11_3_i,temp_b1_11_4_r,temp_b1_11_4_i,temp_b1_12_3_r,temp_b1_12_3_i,temp_b1_12_4_r,temp_b1_12_4_i);
MULT MULT83 (clk,in_11_5_r,in_11_5_i,in_11_6_r,in_11_6_i,in_12_5_r,in_12_5_i,in_12_6_r,in_12_6_i,temp_m1_11_5_r,temp_m1_11_5_i,temp_m1_11_6_r,temp_m1_11_6_i,temp_m1_12_5_r,temp_m1_12_5_i,temp_m1_12_6_r,temp_m1_12_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly83 (clk,temp_m1_11_5_r,temp_m1_11_5_i,temp_m1_11_6_r,temp_m1_11_6_i,temp_m1_12_5_r,temp_m1_12_5_i,temp_m1_12_6_r,temp_m1_12_6_i,temp_b1_11_5_r,temp_b1_11_5_i,temp_b1_11_6_r,temp_b1_11_6_i,temp_b1_12_5_r,temp_b1_12_5_i,temp_b1_12_6_r,temp_b1_12_6_i);
MULT MULT84 (clk,in_11_7_r,in_11_7_i,in_11_8_r,in_11_8_i,in_12_7_r,in_12_7_i,in_12_8_r,in_12_8_i,temp_m1_11_7_r,temp_m1_11_7_i,temp_m1_11_8_r,temp_m1_11_8_i,temp_m1_12_7_r,temp_m1_12_7_i,temp_m1_12_8_r,temp_m1_12_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly84 (clk,temp_m1_11_7_r,temp_m1_11_7_i,temp_m1_11_8_r,temp_m1_11_8_i,temp_m1_12_7_r,temp_m1_12_7_i,temp_m1_12_8_r,temp_m1_12_8_i,temp_b1_11_7_r,temp_b1_11_7_i,temp_b1_11_8_r,temp_b1_11_8_i,temp_b1_12_7_r,temp_b1_12_7_i,temp_b1_12_8_r,temp_b1_12_8_i);
MULT MULT85 (clk,in_11_9_r,in_11_9_i,in_11_10_r,in_11_10_i,in_12_9_r,in_12_9_i,in_12_10_r,in_12_10_i,temp_m1_11_9_r,temp_m1_11_9_i,temp_m1_11_10_r,temp_m1_11_10_i,temp_m1_12_9_r,temp_m1_12_9_i,temp_m1_12_10_r,temp_m1_12_10_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly85 (clk,temp_m1_11_9_r,temp_m1_11_9_i,temp_m1_11_10_r,temp_m1_11_10_i,temp_m1_12_9_r,temp_m1_12_9_i,temp_m1_12_10_r,temp_m1_12_10_i,temp_b1_11_9_r,temp_b1_11_9_i,temp_b1_11_10_r,temp_b1_11_10_i,temp_b1_12_9_r,temp_b1_12_9_i,temp_b1_12_10_r,temp_b1_12_10_i);
MULT MULT86 (clk,in_11_11_r,in_11_11_i,in_11_12_r,in_11_12_i,in_12_11_r,in_12_11_i,in_12_12_r,in_12_12_i,temp_m1_11_11_r,temp_m1_11_11_i,temp_m1_11_12_r,temp_m1_11_12_i,temp_m1_12_11_r,temp_m1_12_11_i,temp_m1_12_12_r,temp_m1_12_12_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly86 (clk,temp_m1_11_11_r,temp_m1_11_11_i,temp_m1_11_12_r,temp_m1_11_12_i,temp_m1_12_11_r,temp_m1_12_11_i,temp_m1_12_12_r,temp_m1_12_12_i,temp_b1_11_11_r,temp_b1_11_11_i,temp_b1_11_12_r,temp_b1_11_12_i,temp_b1_12_11_r,temp_b1_12_11_i,temp_b1_12_12_r,temp_b1_12_12_i);
MULT MULT87 (clk,in_11_13_r,in_11_13_i,in_11_14_r,in_11_14_i,in_12_13_r,in_12_13_i,in_12_14_r,in_12_14_i,temp_m1_11_13_r,temp_m1_11_13_i,temp_m1_11_14_r,temp_m1_11_14_i,temp_m1_12_13_r,temp_m1_12_13_i,temp_m1_12_14_r,temp_m1_12_14_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly87 (clk,temp_m1_11_13_r,temp_m1_11_13_i,temp_m1_11_14_r,temp_m1_11_14_i,temp_m1_12_13_r,temp_m1_12_13_i,temp_m1_12_14_r,temp_m1_12_14_i,temp_b1_11_13_r,temp_b1_11_13_i,temp_b1_11_14_r,temp_b1_11_14_i,temp_b1_12_13_r,temp_b1_12_13_i,temp_b1_12_14_r,temp_b1_12_14_i);
MULT MULT88 (clk,in_11_15_r,in_11_15_i,in_11_16_r,in_11_16_i,in_12_15_r,in_12_15_i,in_12_16_r,in_12_16_i,temp_m1_11_15_r,temp_m1_11_15_i,temp_m1_11_16_r,temp_m1_11_16_i,temp_m1_12_15_r,temp_m1_12_15_i,temp_m1_12_16_r,temp_m1_12_16_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly88 (clk,temp_m1_11_15_r,temp_m1_11_15_i,temp_m1_11_16_r,temp_m1_11_16_i,temp_m1_12_15_r,temp_m1_12_15_i,temp_m1_12_16_r,temp_m1_12_16_i,temp_b1_11_15_r,temp_b1_11_15_i,temp_b1_11_16_r,temp_b1_11_16_i,temp_b1_12_15_r,temp_b1_12_15_i,temp_b1_12_16_r,temp_b1_12_16_i);
MULT MULT89 (clk,in_11_17_r,in_11_17_i,in_11_18_r,in_11_18_i,in_12_17_r,in_12_17_i,in_12_18_r,in_12_18_i,temp_m1_11_17_r,temp_m1_11_17_i,temp_m1_11_18_r,temp_m1_11_18_i,temp_m1_12_17_r,temp_m1_12_17_i,temp_m1_12_18_r,temp_m1_12_18_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly89 (clk,temp_m1_11_17_r,temp_m1_11_17_i,temp_m1_11_18_r,temp_m1_11_18_i,temp_m1_12_17_r,temp_m1_12_17_i,temp_m1_12_18_r,temp_m1_12_18_i,temp_b1_11_17_r,temp_b1_11_17_i,temp_b1_11_18_r,temp_b1_11_18_i,temp_b1_12_17_r,temp_b1_12_17_i,temp_b1_12_18_r,temp_b1_12_18_i);
MULT MULT90 (clk,in_11_19_r,in_11_19_i,in_11_20_r,in_11_20_i,in_12_19_r,in_12_19_i,in_12_20_r,in_12_20_i,temp_m1_11_19_r,temp_m1_11_19_i,temp_m1_11_20_r,temp_m1_11_20_i,temp_m1_12_19_r,temp_m1_12_19_i,temp_m1_12_20_r,temp_m1_12_20_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly90 (clk,temp_m1_11_19_r,temp_m1_11_19_i,temp_m1_11_20_r,temp_m1_11_20_i,temp_m1_12_19_r,temp_m1_12_19_i,temp_m1_12_20_r,temp_m1_12_20_i,temp_b1_11_19_r,temp_b1_11_19_i,temp_b1_11_20_r,temp_b1_11_20_i,temp_b1_12_19_r,temp_b1_12_19_i,temp_b1_12_20_r,temp_b1_12_20_i);
MULT MULT91 (clk,in_11_21_r,in_11_21_i,in_11_22_r,in_11_22_i,in_12_21_r,in_12_21_i,in_12_22_r,in_12_22_i,temp_m1_11_21_r,temp_m1_11_21_i,temp_m1_11_22_r,temp_m1_11_22_i,temp_m1_12_21_r,temp_m1_12_21_i,temp_m1_12_22_r,temp_m1_12_22_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly91 (clk,temp_m1_11_21_r,temp_m1_11_21_i,temp_m1_11_22_r,temp_m1_11_22_i,temp_m1_12_21_r,temp_m1_12_21_i,temp_m1_12_22_r,temp_m1_12_22_i,temp_b1_11_21_r,temp_b1_11_21_i,temp_b1_11_22_r,temp_b1_11_22_i,temp_b1_12_21_r,temp_b1_12_21_i,temp_b1_12_22_r,temp_b1_12_22_i);
MULT MULT92 (clk,in_11_23_r,in_11_23_i,in_11_24_r,in_11_24_i,in_12_23_r,in_12_23_i,in_12_24_r,in_12_24_i,temp_m1_11_23_r,temp_m1_11_23_i,temp_m1_11_24_r,temp_m1_11_24_i,temp_m1_12_23_r,temp_m1_12_23_i,temp_m1_12_24_r,temp_m1_12_24_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly92 (clk,temp_m1_11_23_r,temp_m1_11_23_i,temp_m1_11_24_r,temp_m1_11_24_i,temp_m1_12_23_r,temp_m1_12_23_i,temp_m1_12_24_r,temp_m1_12_24_i,temp_b1_11_23_r,temp_b1_11_23_i,temp_b1_11_24_r,temp_b1_11_24_i,temp_b1_12_23_r,temp_b1_12_23_i,temp_b1_12_24_r,temp_b1_12_24_i);
MULT MULT93 (clk,in_11_25_r,in_11_25_i,in_11_26_r,in_11_26_i,in_12_25_r,in_12_25_i,in_12_26_r,in_12_26_i,temp_m1_11_25_r,temp_m1_11_25_i,temp_m1_11_26_r,temp_m1_11_26_i,temp_m1_12_25_r,temp_m1_12_25_i,temp_m1_12_26_r,temp_m1_12_26_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly93 (clk,temp_m1_11_25_r,temp_m1_11_25_i,temp_m1_11_26_r,temp_m1_11_26_i,temp_m1_12_25_r,temp_m1_12_25_i,temp_m1_12_26_r,temp_m1_12_26_i,temp_b1_11_25_r,temp_b1_11_25_i,temp_b1_11_26_r,temp_b1_11_26_i,temp_b1_12_25_r,temp_b1_12_25_i,temp_b1_12_26_r,temp_b1_12_26_i);
MULT MULT94 (clk,in_11_27_r,in_11_27_i,in_11_28_r,in_11_28_i,in_12_27_r,in_12_27_i,in_12_28_r,in_12_28_i,temp_m1_11_27_r,temp_m1_11_27_i,temp_m1_11_28_r,temp_m1_11_28_i,temp_m1_12_27_r,temp_m1_12_27_i,temp_m1_12_28_r,temp_m1_12_28_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly94 (clk,temp_m1_11_27_r,temp_m1_11_27_i,temp_m1_11_28_r,temp_m1_11_28_i,temp_m1_12_27_r,temp_m1_12_27_i,temp_m1_12_28_r,temp_m1_12_28_i,temp_b1_11_27_r,temp_b1_11_27_i,temp_b1_11_28_r,temp_b1_11_28_i,temp_b1_12_27_r,temp_b1_12_27_i,temp_b1_12_28_r,temp_b1_12_28_i);
MULT MULT95 (clk,in_11_29_r,in_11_29_i,in_11_30_r,in_11_30_i,in_12_29_r,in_12_29_i,in_12_30_r,in_12_30_i,temp_m1_11_29_r,temp_m1_11_29_i,temp_m1_11_30_r,temp_m1_11_30_i,temp_m1_12_29_r,temp_m1_12_29_i,temp_m1_12_30_r,temp_m1_12_30_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly95 (clk,temp_m1_11_29_r,temp_m1_11_29_i,temp_m1_11_30_r,temp_m1_11_30_i,temp_m1_12_29_r,temp_m1_12_29_i,temp_m1_12_30_r,temp_m1_12_30_i,temp_b1_11_29_r,temp_b1_11_29_i,temp_b1_11_30_r,temp_b1_11_30_i,temp_b1_12_29_r,temp_b1_12_29_i,temp_b1_12_30_r,temp_b1_12_30_i);
MULT MULT96 (clk,in_11_31_r,in_11_31_i,in_11_32_r,in_11_32_i,in_12_31_r,in_12_31_i,in_12_32_r,in_12_32_i,temp_m1_11_31_r,temp_m1_11_31_i,temp_m1_11_32_r,temp_m1_11_32_i,temp_m1_12_31_r,temp_m1_12_31_i,temp_m1_12_32_r,temp_m1_12_32_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly96 (clk,temp_m1_11_31_r,temp_m1_11_31_i,temp_m1_11_32_r,temp_m1_11_32_i,temp_m1_12_31_r,temp_m1_12_31_i,temp_m1_12_32_r,temp_m1_12_32_i,temp_b1_11_31_r,temp_b1_11_31_i,temp_b1_11_32_r,temp_b1_11_32_i,temp_b1_12_31_r,temp_b1_12_31_i,temp_b1_12_32_r,temp_b1_12_32_i);
MULT MULT97 (clk,in_13_1_r,in_13_1_i,in_13_2_r,in_13_2_i,in_14_1_r,in_14_1_i,in_14_2_r,in_14_2_i,temp_m1_13_1_r,temp_m1_13_1_i,temp_m1_13_2_r,temp_m1_13_2_i,temp_m1_14_1_r,temp_m1_14_1_i,temp_m1_14_2_r,temp_m1_14_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly97 (clk,temp_m1_13_1_r,temp_m1_13_1_i,temp_m1_13_2_r,temp_m1_13_2_i,temp_m1_14_1_r,temp_m1_14_1_i,temp_m1_14_2_r,temp_m1_14_2_i,temp_b1_13_1_r,temp_b1_13_1_i,temp_b1_13_2_r,temp_b1_13_2_i,temp_b1_14_1_r,temp_b1_14_1_i,temp_b1_14_2_r,temp_b1_14_2_i);
MULT MULT98 (clk,in_13_3_r,in_13_3_i,in_13_4_r,in_13_4_i,in_14_3_r,in_14_3_i,in_14_4_r,in_14_4_i,temp_m1_13_3_r,temp_m1_13_3_i,temp_m1_13_4_r,temp_m1_13_4_i,temp_m1_14_3_r,temp_m1_14_3_i,temp_m1_14_4_r,temp_m1_14_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly98 (clk,temp_m1_13_3_r,temp_m1_13_3_i,temp_m1_13_4_r,temp_m1_13_4_i,temp_m1_14_3_r,temp_m1_14_3_i,temp_m1_14_4_r,temp_m1_14_4_i,temp_b1_13_3_r,temp_b1_13_3_i,temp_b1_13_4_r,temp_b1_13_4_i,temp_b1_14_3_r,temp_b1_14_3_i,temp_b1_14_4_r,temp_b1_14_4_i);
MULT MULT99 (clk,in_13_5_r,in_13_5_i,in_13_6_r,in_13_6_i,in_14_5_r,in_14_5_i,in_14_6_r,in_14_6_i,temp_m1_13_5_r,temp_m1_13_5_i,temp_m1_13_6_r,temp_m1_13_6_i,temp_m1_14_5_r,temp_m1_14_5_i,temp_m1_14_6_r,temp_m1_14_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly99 (clk,temp_m1_13_5_r,temp_m1_13_5_i,temp_m1_13_6_r,temp_m1_13_6_i,temp_m1_14_5_r,temp_m1_14_5_i,temp_m1_14_6_r,temp_m1_14_6_i,temp_b1_13_5_r,temp_b1_13_5_i,temp_b1_13_6_r,temp_b1_13_6_i,temp_b1_14_5_r,temp_b1_14_5_i,temp_b1_14_6_r,temp_b1_14_6_i);
MULT MULT100 (clk,in_13_7_r,in_13_7_i,in_13_8_r,in_13_8_i,in_14_7_r,in_14_7_i,in_14_8_r,in_14_8_i,temp_m1_13_7_r,temp_m1_13_7_i,temp_m1_13_8_r,temp_m1_13_8_i,temp_m1_14_7_r,temp_m1_14_7_i,temp_m1_14_8_r,temp_m1_14_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly100 (clk,temp_m1_13_7_r,temp_m1_13_7_i,temp_m1_13_8_r,temp_m1_13_8_i,temp_m1_14_7_r,temp_m1_14_7_i,temp_m1_14_8_r,temp_m1_14_8_i,temp_b1_13_7_r,temp_b1_13_7_i,temp_b1_13_8_r,temp_b1_13_8_i,temp_b1_14_7_r,temp_b1_14_7_i,temp_b1_14_8_r,temp_b1_14_8_i);
MULT MULT101 (clk,in_13_9_r,in_13_9_i,in_13_10_r,in_13_10_i,in_14_9_r,in_14_9_i,in_14_10_r,in_14_10_i,temp_m1_13_9_r,temp_m1_13_9_i,temp_m1_13_10_r,temp_m1_13_10_i,temp_m1_14_9_r,temp_m1_14_9_i,temp_m1_14_10_r,temp_m1_14_10_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly101 (clk,temp_m1_13_9_r,temp_m1_13_9_i,temp_m1_13_10_r,temp_m1_13_10_i,temp_m1_14_9_r,temp_m1_14_9_i,temp_m1_14_10_r,temp_m1_14_10_i,temp_b1_13_9_r,temp_b1_13_9_i,temp_b1_13_10_r,temp_b1_13_10_i,temp_b1_14_9_r,temp_b1_14_9_i,temp_b1_14_10_r,temp_b1_14_10_i);
MULT MULT102 (clk,in_13_11_r,in_13_11_i,in_13_12_r,in_13_12_i,in_14_11_r,in_14_11_i,in_14_12_r,in_14_12_i,temp_m1_13_11_r,temp_m1_13_11_i,temp_m1_13_12_r,temp_m1_13_12_i,temp_m1_14_11_r,temp_m1_14_11_i,temp_m1_14_12_r,temp_m1_14_12_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly102 (clk,temp_m1_13_11_r,temp_m1_13_11_i,temp_m1_13_12_r,temp_m1_13_12_i,temp_m1_14_11_r,temp_m1_14_11_i,temp_m1_14_12_r,temp_m1_14_12_i,temp_b1_13_11_r,temp_b1_13_11_i,temp_b1_13_12_r,temp_b1_13_12_i,temp_b1_14_11_r,temp_b1_14_11_i,temp_b1_14_12_r,temp_b1_14_12_i);
MULT MULT103 (clk,in_13_13_r,in_13_13_i,in_13_14_r,in_13_14_i,in_14_13_r,in_14_13_i,in_14_14_r,in_14_14_i,temp_m1_13_13_r,temp_m1_13_13_i,temp_m1_13_14_r,temp_m1_13_14_i,temp_m1_14_13_r,temp_m1_14_13_i,temp_m1_14_14_r,temp_m1_14_14_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly103 (clk,temp_m1_13_13_r,temp_m1_13_13_i,temp_m1_13_14_r,temp_m1_13_14_i,temp_m1_14_13_r,temp_m1_14_13_i,temp_m1_14_14_r,temp_m1_14_14_i,temp_b1_13_13_r,temp_b1_13_13_i,temp_b1_13_14_r,temp_b1_13_14_i,temp_b1_14_13_r,temp_b1_14_13_i,temp_b1_14_14_r,temp_b1_14_14_i);
MULT MULT104 (clk,in_13_15_r,in_13_15_i,in_13_16_r,in_13_16_i,in_14_15_r,in_14_15_i,in_14_16_r,in_14_16_i,temp_m1_13_15_r,temp_m1_13_15_i,temp_m1_13_16_r,temp_m1_13_16_i,temp_m1_14_15_r,temp_m1_14_15_i,temp_m1_14_16_r,temp_m1_14_16_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly104 (clk,temp_m1_13_15_r,temp_m1_13_15_i,temp_m1_13_16_r,temp_m1_13_16_i,temp_m1_14_15_r,temp_m1_14_15_i,temp_m1_14_16_r,temp_m1_14_16_i,temp_b1_13_15_r,temp_b1_13_15_i,temp_b1_13_16_r,temp_b1_13_16_i,temp_b1_14_15_r,temp_b1_14_15_i,temp_b1_14_16_r,temp_b1_14_16_i);
MULT MULT105 (clk,in_13_17_r,in_13_17_i,in_13_18_r,in_13_18_i,in_14_17_r,in_14_17_i,in_14_18_r,in_14_18_i,temp_m1_13_17_r,temp_m1_13_17_i,temp_m1_13_18_r,temp_m1_13_18_i,temp_m1_14_17_r,temp_m1_14_17_i,temp_m1_14_18_r,temp_m1_14_18_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly105 (clk,temp_m1_13_17_r,temp_m1_13_17_i,temp_m1_13_18_r,temp_m1_13_18_i,temp_m1_14_17_r,temp_m1_14_17_i,temp_m1_14_18_r,temp_m1_14_18_i,temp_b1_13_17_r,temp_b1_13_17_i,temp_b1_13_18_r,temp_b1_13_18_i,temp_b1_14_17_r,temp_b1_14_17_i,temp_b1_14_18_r,temp_b1_14_18_i);
MULT MULT106 (clk,in_13_19_r,in_13_19_i,in_13_20_r,in_13_20_i,in_14_19_r,in_14_19_i,in_14_20_r,in_14_20_i,temp_m1_13_19_r,temp_m1_13_19_i,temp_m1_13_20_r,temp_m1_13_20_i,temp_m1_14_19_r,temp_m1_14_19_i,temp_m1_14_20_r,temp_m1_14_20_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly106 (clk,temp_m1_13_19_r,temp_m1_13_19_i,temp_m1_13_20_r,temp_m1_13_20_i,temp_m1_14_19_r,temp_m1_14_19_i,temp_m1_14_20_r,temp_m1_14_20_i,temp_b1_13_19_r,temp_b1_13_19_i,temp_b1_13_20_r,temp_b1_13_20_i,temp_b1_14_19_r,temp_b1_14_19_i,temp_b1_14_20_r,temp_b1_14_20_i);
MULT MULT107 (clk,in_13_21_r,in_13_21_i,in_13_22_r,in_13_22_i,in_14_21_r,in_14_21_i,in_14_22_r,in_14_22_i,temp_m1_13_21_r,temp_m1_13_21_i,temp_m1_13_22_r,temp_m1_13_22_i,temp_m1_14_21_r,temp_m1_14_21_i,temp_m1_14_22_r,temp_m1_14_22_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly107 (clk,temp_m1_13_21_r,temp_m1_13_21_i,temp_m1_13_22_r,temp_m1_13_22_i,temp_m1_14_21_r,temp_m1_14_21_i,temp_m1_14_22_r,temp_m1_14_22_i,temp_b1_13_21_r,temp_b1_13_21_i,temp_b1_13_22_r,temp_b1_13_22_i,temp_b1_14_21_r,temp_b1_14_21_i,temp_b1_14_22_r,temp_b1_14_22_i);
MULT MULT108 (clk,in_13_23_r,in_13_23_i,in_13_24_r,in_13_24_i,in_14_23_r,in_14_23_i,in_14_24_r,in_14_24_i,temp_m1_13_23_r,temp_m1_13_23_i,temp_m1_13_24_r,temp_m1_13_24_i,temp_m1_14_23_r,temp_m1_14_23_i,temp_m1_14_24_r,temp_m1_14_24_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly108 (clk,temp_m1_13_23_r,temp_m1_13_23_i,temp_m1_13_24_r,temp_m1_13_24_i,temp_m1_14_23_r,temp_m1_14_23_i,temp_m1_14_24_r,temp_m1_14_24_i,temp_b1_13_23_r,temp_b1_13_23_i,temp_b1_13_24_r,temp_b1_13_24_i,temp_b1_14_23_r,temp_b1_14_23_i,temp_b1_14_24_r,temp_b1_14_24_i);
MULT MULT109 (clk,in_13_25_r,in_13_25_i,in_13_26_r,in_13_26_i,in_14_25_r,in_14_25_i,in_14_26_r,in_14_26_i,temp_m1_13_25_r,temp_m1_13_25_i,temp_m1_13_26_r,temp_m1_13_26_i,temp_m1_14_25_r,temp_m1_14_25_i,temp_m1_14_26_r,temp_m1_14_26_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly109 (clk,temp_m1_13_25_r,temp_m1_13_25_i,temp_m1_13_26_r,temp_m1_13_26_i,temp_m1_14_25_r,temp_m1_14_25_i,temp_m1_14_26_r,temp_m1_14_26_i,temp_b1_13_25_r,temp_b1_13_25_i,temp_b1_13_26_r,temp_b1_13_26_i,temp_b1_14_25_r,temp_b1_14_25_i,temp_b1_14_26_r,temp_b1_14_26_i);
MULT MULT110 (clk,in_13_27_r,in_13_27_i,in_13_28_r,in_13_28_i,in_14_27_r,in_14_27_i,in_14_28_r,in_14_28_i,temp_m1_13_27_r,temp_m1_13_27_i,temp_m1_13_28_r,temp_m1_13_28_i,temp_m1_14_27_r,temp_m1_14_27_i,temp_m1_14_28_r,temp_m1_14_28_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly110 (clk,temp_m1_13_27_r,temp_m1_13_27_i,temp_m1_13_28_r,temp_m1_13_28_i,temp_m1_14_27_r,temp_m1_14_27_i,temp_m1_14_28_r,temp_m1_14_28_i,temp_b1_13_27_r,temp_b1_13_27_i,temp_b1_13_28_r,temp_b1_13_28_i,temp_b1_14_27_r,temp_b1_14_27_i,temp_b1_14_28_r,temp_b1_14_28_i);
MULT MULT111 (clk,in_13_29_r,in_13_29_i,in_13_30_r,in_13_30_i,in_14_29_r,in_14_29_i,in_14_30_r,in_14_30_i,temp_m1_13_29_r,temp_m1_13_29_i,temp_m1_13_30_r,temp_m1_13_30_i,temp_m1_14_29_r,temp_m1_14_29_i,temp_m1_14_30_r,temp_m1_14_30_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly111 (clk,temp_m1_13_29_r,temp_m1_13_29_i,temp_m1_13_30_r,temp_m1_13_30_i,temp_m1_14_29_r,temp_m1_14_29_i,temp_m1_14_30_r,temp_m1_14_30_i,temp_b1_13_29_r,temp_b1_13_29_i,temp_b1_13_30_r,temp_b1_13_30_i,temp_b1_14_29_r,temp_b1_14_29_i,temp_b1_14_30_r,temp_b1_14_30_i);
MULT MULT112 (clk,in_13_31_r,in_13_31_i,in_13_32_r,in_13_32_i,in_14_31_r,in_14_31_i,in_14_32_r,in_14_32_i,temp_m1_13_31_r,temp_m1_13_31_i,temp_m1_13_32_r,temp_m1_13_32_i,temp_m1_14_31_r,temp_m1_14_31_i,temp_m1_14_32_r,temp_m1_14_32_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly112 (clk,temp_m1_13_31_r,temp_m1_13_31_i,temp_m1_13_32_r,temp_m1_13_32_i,temp_m1_14_31_r,temp_m1_14_31_i,temp_m1_14_32_r,temp_m1_14_32_i,temp_b1_13_31_r,temp_b1_13_31_i,temp_b1_13_32_r,temp_b1_13_32_i,temp_b1_14_31_r,temp_b1_14_31_i,temp_b1_14_32_r,temp_b1_14_32_i);
MULT MULT113 (clk,in_15_1_r,in_15_1_i,in_15_2_r,in_15_2_i,in_16_1_r,in_16_1_i,in_16_2_r,in_16_2_i,temp_m1_15_1_r,temp_m1_15_1_i,temp_m1_15_2_r,temp_m1_15_2_i,temp_m1_16_1_r,temp_m1_16_1_i,temp_m1_16_2_r,temp_m1_16_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly113 (clk,temp_m1_15_1_r,temp_m1_15_1_i,temp_m1_15_2_r,temp_m1_15_2_i,temp_m1_16_1_r,temp_m1_16_1_i,temp_m1_16_2_r,temp_m1_16_2_i,temp_b1_15_1_r,temp_b1_15_1_i,temp_b1_15_2_r,temp_b1_15_2_i,temp_b1_16_1_r,temp_b1_16_1_i,temp_b1_16_2_r,temp_b1_16_2_i);
MULT MULT114 (clk,in_15_3_r,in_15_3_i,in_15_4_r,in_15_4_i,in_16_3_r,in_16_3_i,in_16_4_r,in_16_4_i,temp_m1_15_3_r,temp_m1_15_3_i,temp_m1_15_4_r,temp_m1_15_4_i,temp_m1_16_3_r,temp_m1_16_3_i,temp_m1_16_4_r,temp_m1_16_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly114 (clk,temp_m1_15_3_r,temp_m1_15_3_i,temp_m1_15_4_r,temp_m1_15_4_i,temp_m1_16_3_r,temp_m1_16_3_i,temp_m1_16_4_r,temp_m1_16_4_i,temp_b1_15_3_r,temp_b1_15_3_i,temp_b1_15_4_r,temp_b1_15_4_i,temp_b1_16_3_r,temp_b1_16_3_i,temp_b1_16_4_r,temp_b1_16_4_i);
MULT MULT115 (clk,in_15_5_r,in_15_5_i,in_15_6_r,in_15_6_i,in_16_5_r,in_16_5_i,in_16_6_r,in_16_6_i,temp_m1_15_5_r,temp_m1_15_5_i,temp_m1_15_6_r,temp_m1_15_6_i,temp_m1_16_5_r,temp_m1_16_5_i,temp_m1_16_6_r,temp_m1_16_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly115 (clk,temp_m1_15_5_r,temp_m1_15_5_i,temp_m1_15_6_r,temp_m1_15_6_i,temp_m1_16_5_r,temp_m1_16_5_i,temp_m1_16_6_r,temp_m1_16_6_i,temp_b1_15_5_r,temp_b1_15_5_i,temp_b1_15_6_r,temp_b1_15_6_i,temp_b1_16_5_r,temp_b1_16_5_i,temp_b1_16_6_r,temp_b1_16_6_i);
MULT MULT116 (clk,in_15_7_r,in_15_7_i,in_15_8_r,in_15_8_i,in_16_7_r,in_16_7_i,in_16_8_r,in_16_8_i,temp_m1_15_7_r,temp_m1_15_7_i,temp_m1_15_8_r,temp_m1_15_8_i,temp_m1_16_7_r,temp_m1_16_7_i,temp_m1_16_8_r,temp_m1_16_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly116 (clk,temp_m1_15_7_r,temp_m1_15_7_i,temp_m1_15_8_r,temp_m1_15_8_i,temp_m1_16_7_r,temp_m1_16_7_i,temp_m1_16_8_r,temp_m1_16_8_i,temp_b1_15_7_r,temp_b1_15_7_i,temp_b1_15_8_r,temp_b1_15_8_i,temp_b1_16_7_r,temp_b1_16_7_i,temp_b1_16_8_r,temp_b1_16_8_i);
MULT MULT117 (clk,in_15_9_r,in_15_9_i,in_15_10_r,in_15_10_i,in_16_9_r,in_16_9_i,in_16_10_r,in_16_10_i,temp_m1_15_9_r,temp_m1_15_9_i,temp_m1_15_10_r,temp_m1_15_10_i,temp_m1_16_9_r,temp_m1_16_9_i,temp_m1_16_10_r,temp_m1_16_10_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly117 (clk,temp_m1_15_9_r,temp_m1_15_9_i,temp_m1_15_10_r,temp_m1_15_10_i,temp_m1_16_9_r,temp_m1_16_9_i,temp_m1_16_10_r,temp_m1_16_10_i,temp_b1_15_9_r,temp_b1_15_9_i,temp_b1_15_10_r,temp_b1_15_10_i,temp_b1_16_9_r,temp_b1_16_9_i,temp_b1_16_10_r,temp_b1_16_10_i);
MULT MULT118 (clk,in_15_11_r,in_15_11_i,in_15_12_r,in_15_12_i,in_16_11_r,in_16_11_i,in_16_12_r,in_16_12_i,temp_m1_15_11_r,temp_m1_15_11_i,temp_m1_15_12_r,temp_m1_15_12_i,temp_m1_16_11_r,temp_m1_16_11_i,temp_m1_16_12_r,temp_m1_16_12_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly118 (clk,temp_m1_15_11_r,temp_m1_15_11_i,temp_m1_15_12_r,temp_m1_15_12_i,temp_m1_16_11_r,temp_m1_16_11_i,temp_m1_16_12_r,temp_m1_16_12_i,temp_b1_15_11_r,temp_b1_15_11_i,temp_b1_15_12_r,temp_b1_15_12_i,temp_b1_16_11_r,temp_b1_16_11_i,temp_b1_16_12_r,temp_b1_16_12_i);
MULT MULT119 (clk,in_15_13_r,in_15_13_i,in_15_14_r,in_15_14_i,in_16_13_r,in_16_13_i,in_16_14_r,in_16_14_i,temp_m1_15_13_r,temp_m1_15_13_i,temp_m1_15_14_r,temp_m1_15_14_i,temp_m1_16_13_r,temp_m1_16_13_i,temp_m1_16_14_r,temp_m1_16_14_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly119 (clk,temp_m1_15_13_r,temp_m1_15_13_i,temp_m1_15_14_r,temp_m1_15_14_i,temp_m1_16_13_r,temp_m1_16_13_i,temp_m1_16_14_r,temp_m1_16_14_i,temp_b1_15_13_r,temp_b1_15_13_i,temp_b1_15_14_r,temp_b1_15_14_i,temp_b1_16_13_r,temp_b1_16_13_i,temp_b1_16_14_r,temp_b1_16_14_i);
MULT MULT120 (clk,in_15_15_r,in_15_15_i,in_15_16_r,in_15_16_i,in_16_15_r,in_16_15_i,in_16_16_r,in_16_16_i,temp_m1_15_15_r,temp_m1_15_15_i,temp_m1_15_16_r,temp_m1_15_16_i,temp_m1_16_15_r,temp_m1_16_15_i,temp_m1_16_16_r,temp_m1_16_16_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly120 (clk,temp_m1_15_15_r,temp_m1_15_15_i,temp_m1_15_16_r,temp_m1_15_16_i,temp_m1_16_15_r,temp_m1_16_15_i,temp_m1_16_16_r,temp_m1_16_16_i,temp_b1_15_15_r,temp_b1_15_15_i,temp_b1_15_16_r,temp_b1_15_16_i,temp_b1_16_15_r,temp_b1_16_15_i,temp_b1_16_16_r,temp_b1_16_16_i);
MULT MULT121 (clk,in_15_17_r,in_15_17_i,in_15_18_r,in_15_18_i,in_16_17_r,in_16_17_i,in_16_18_r,in_16_18_i,temp_m1_15_17_r,temp_m1_15_17_i,temp_m1_15_18_r,temp_m1_15_18_i,temp_m1_16_17_r,temp_m1_16_17_i,temp_m1_16_18_r,temp_m1_16_18_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly121 (clk,temp_m1_15_17_r,temp_m1_15_17_i,temp_m1_15_18_r,temp_m1_15_18_i,temp_m1_16_17_r,temp_m1_16_17_i,temp_m1_16_18_r,temp_m1_16_18_i,temp_b1_15_17_r,temp_b1_15_17_i,temp_b1_15_18_r,temp_b1_15_18_i,temp_b1_16_17_r,temp_b1_16_17_i,temp_b1_16_18_r,temp_b1_16_18_i);
MULT MULT122 (clk,in_15_19_r,in_15_19_i,in_15_20_r,in_15_20_i,in_16_19_r,in_16_19_i,in_16_20_r,in_16_20_i,temp_m1_15_19_r,temp_m1_15_19_i,temp_m1_15_20_r,temp_m1_15_20_i,temp_m1_16_19_r,temp_m1_16_19_i,temp_m1_16_20_r,temp_m1_16_20_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly122 (clk,temp_m1_15_19_r,temp_m1_15_19_i,temp_m1_15_20_r,temp_m1_15_20_i,temp_m1_16_19_r,temp_m1_16_19_i,temp_m1_16_20_r,temp_m1_16_20_i,temp_b1_15_19_r,temp_b1_15_19_i,temp_b1_15_20_r,temp_b1_15_20_i,temp_b1_16_19_r,temp_b1_16_19_i,temp_b1_16_20_r,temp_b1_16_20_i);
MULT MULT123 (clk,in_15_21_r,in_15_21_i,in_15_22_r,in_15_22_i,in_16_21_r,in_16_21_i,in_16_22_r,in_16_22_i,temp_m1_15_21_r,temp_m1_15_21_i,temp_m1_15_22_r,temp_m1_15_22_i,temp_m1_16_21_r,temp_m1_16_21_i,temp_m1_16_22_r,temp_m1_16_22_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly123 (clk,temp_m1_15_21_r,temp_m1_15_21_i,temp_m1_15_22_r,temp_m1_15_22_i,temp_m1_16_21_r,temp_m1_16_21_i,temp_m1_16_22_r,temp_m1_16_22_i,temp_b1_15_21_r,temp_b1_15_21_i,temp_b1_15_22_r,temp_b1_15_22_i,temp_b1_16_21_r,temp_b1_16_21_i,temp_b1_16_22_r,temp_b1_16_22_i);
MULT MULT124 (clk,in_15_23_r,in_15_23_i,in_15_24_r,in_15_24_i,in_16_23_r,in_16_23_i,in_16_24_r,in_16_24_i,temp_m1_15_23_r,temp_m1_15_23_i,temp_m1_15_24_r,temp_m1_15_24_i,temp_m1_16_23_r,temp_m1_16_23_i,temp_m1_16_24_r,temp_m1_16_24_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly124 (clk,temp_m1_15_23_r,temp_m1_15_23_i,temp_m1_15_24_r,temp_m1_15_24_i,temp_m1_16_23_r,temp_m1_16_23_i,temp_m1_16_24_r,temp_m1_16_24_i,temp_b1_15_23_r,temp_b1_15_23_i,temp_b1_15_24_r,temp_b1_15_24_i,temp_b1_16_23_r,temp_b1_16_23_i,temp_b1_16_24_r,temp_b1_16_24_i);
MULT MULT125 (clk,in_15_25_r,in_15_25_i,in_15_26_r,in_15_26_i,in_16_25_r,in_16_25_i,in_16_26_r,in_16_26_i,temp_m1_15_25_r,temp_m1_15_25_i,temp_m1_15_26_r,temp_m1_15_26_i,temp_m1_16_25_r,temp_m1_16_25_i,temp_m1_16_26_r,temp_m1_16_26_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly125 (clk,temp_m1_15_25_r,temp_m1_15_25_i,temp_m1_15_26_r,temp_m1_15_26_i,temp_m1_16_25_r,temp_m1_16_25_i,temp_m1_16_26_r,temp_m1_16_26_i,temp_b1_15_25_r,temp_b1_15_25_i,temp_b1_15_26_r,temp_b1_15_26_i,temp_b1_16_25_r,temp_b1_16_25_i,temp_b1_16_26_r,temp_b1_16_26_i);
MULT MULT126 (clk,in_15_27_r,in_15_27_i,in_15_28_r,in_15_28_i,in_16_27_r,in_16_27_i,in_16_28_r,in_16_28_i,temp_m1_15_27_r,temp_m1_15_27_i,temp_m1_15_28_r,temp_m1_15_28_i,temp_m1_16_27_r,temp_m1_16_27_i,temp_m1_16_28_r,temp_m1_16_28_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly126 (clk,temp_m1_15_27_r,temp_m1_15_27_i,temp_m1_15_28_r,temp_m1_15_28_i,temp_m1_16_27_r,temp_m1_16_27_i,temp_m1_16_28_r,temp_m1_16_28_i,temp_b1_15_27_r,temp_b1_15_27_i,temp_b1_15_28_r,temp_b1_15_28_i,temp_b1_16_27_r,temp_b1_16_27_i,temp_b1_16_28_r,temp_b1_16_28_i);
MULT MULT127 (clk,in_15_29_r,in_15_29_i,in_15_30_r,in_15_30_i,in_16_29_r,in_16_29_i,in_16_30_r,in_16_30_i,temp_m1_15_29_r,temp_m1_15_29_i,temp_m1_15_30_r,temp_m1_15_30_i,temp_m1_16_29_r,temp_m1_16_29_i,temp_m1_16_30_r,temp_m1_16_30_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly127 (clk,temp_m1_15_29_r,temp_m1_15_29_i,temp_m1_15_30_r,temp_m1_15_30_i,temp_m1_16_29_r,temp_m1_16_29_i,temp_m1_16_30_r,temp_m1_16_30_i,temp_b1_15_29_r,temp_b1_15_29_i,temp_b1_15_30_r,temp_b1_15_30_i,temp_b1_16_29_r,temp_b1_16_29_i,temp_b1_16_30_r,temp_b1_16_30_i);
MULT MULT128 (clk,in_15_31_r,in_15_31_i,in_15_32_r,in_15_32_i,in_16_31_r,in_16_31_i,in_16_32_r,in_16_32_i,temp_m1_15_31_r,temp_m1_15_31_i,temp_m1_15_32_r,temp_m1_15_32_i,temp_m1_16_31_r,temp_m1_16_31_i,temp_m1_16_32_r,temp_m1_16_32_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly128 (clk,temp_m1_15_31_r,temp_m1_15_31_i,temp_m1_15_32_r,temp_m1_15_32_i,temp_m1_16_31_r,temp_m1_16_31_i,temp_m1_16_32_r,temp_m1_16_32_i,temp_b1_15_31_r,temp_b1_15_31_i,temp_b1_15_32_r,temp_b1_15_32_i,temp_b1_16_31_r,temp_b1_16_31_i,temp_b1_16_32_r,temp_b1_16_32_i);
MULT MULT129 (clk,in_17_1_r,in_17_1_i,in_17_2_r,in_17_2_i,in_18_1_r,in_18_1_i,in_18_2_r,in_18_2_i,temp_m1_17_1_r,temp_m1_17_1_i,temp_m1_17_2_r,temp_m1_17_2_i,temp_m1_18_1_r,temp_m1_18_1_i,temp_m1_18_2_r,temp_m1_18_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly129 (clk,temp_m1_17_1_r,temp_m1_17_1_i,temp_m1_17_2_r,temp_m1_17_2_i,temp_m1_18_1_r,temp_m1_18_1_i,temp_m1_18_2_r,temp_m1_18_2_i,temp_b1_17_1_r,temp_b1_17_1_i,temp_b1_17_2_r,temp_b1_17_2_i,temp_b1_18_1_r,temp_b1_18_1_i,temp_b1_18_2_r,temp_b1_18_2_i);
MULT MULT130 (clk,in_17_3_r,in_17_3_i,in_17_4_r,in_17_4_i,in_18_3_r,in_18_3_i,in_18_4_r,in_18_4_i,temp_m1_17_3_r,temp_m1_17_3_i,temp_m1_17_4_r,temp_m1_17_4_i,temp_m1_18_3_r,temp_m1_18_3_i,temp_m1_18_4_r,temp_m1_18_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly130 (clk,temp_m1_17_3_r,temp_m1_17_3_i,temp_m1_17_4_r,temp_m1_17_4_i,temp_m1_18_3_r,temp_m1_18_3_i,temp_m1_18_4_r,temp_m1_18_4_i,temp_b1_17_3_r,temp_b1_17_3_i,temp_b1_17_4_r,temp_b1_17_4_i,temp_b1_18_3_r,temp_b1_18_3_i,temp_b1_18_4_r,temp_b1_18_4_i);
MULT MULT131 (clk,in_17_5_r,in_17_5_i,in_17_6_r,in_17_6_i,in_18_5_r,in_18_5_i,in_18_6_r,in_18_6_i,temp_m1_17_5_r,temp_m1_17_5_i,temp_m1_17_6_r,temp_m1_17_6_i,temp_m1_18_5_r,temp_m1_18_5_i,temp_m1_18_6_r,temp_m1_18_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly131 (clk,temp_m1_17_5_r,temp_m1_17_5_i,temp_m1_17_6_r,temp_m1_17_6_i,temp_m1_18_5_r,temp_m1_18_5_i,temp_m1_18_6_r,temp_m1_18_6_i,temp_b1_17_5_r,temp_b1_17_5_i,temp_b1_17_6_r,temp_b1_17_6_i,temp_b1_18_5_r,temp_b1_18_5_i,temp_b1_18_6_r,temp_b1_18_6_i);
MULT MULT132 (clk,in_17_7_r,in_17_7_i,in_17_8_r,in_17_8_i,in_18_7_r,in_18_7_i,in_18_8_r,in_18_8_i,temp_m1_17_7_r,temp_m1_17_7_i,temp_m1_17_8_r,temp_m1_17_8_i,temp_m1_18_7_r,temp_m1_18_7_i,temp_m1_18_8_r,temp_m1_18_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly132 (clk,temp_m1_17_7_r,temp_m1_17_7_i,temp_m1_17_8_r,temp_m1_17_8_i,temp_m1_18_7_r,temp_m1_18_7_i,temp_m1_18_8_r,temp_m1_18_8_i,temp_b1_17_7_r,temp_b1_17_7_i,temp_b1_17_8_r,temp_b1_17_8_i,temp_b1_18_7_r,temp_b1_18_7_i,temp_b1_18_8_r,temp_b1_18_8_i);
MULT MULT133 (clk,in_17_9_r,in_17_9_i,in_17_10_r,in_17_10_i,in_18_9_r,in_18_9_i,in_18_10_r,in_18_10_i,temp_m1_17_9_r,temp_m1_17_9_i,temp_m1_17_10_r,temp_m1_17_10_i,temp_m1_18_9_r,temp_m1_18_9_i,temp_m1_18_10_r,temp_m1_18_10_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly133 (clk,temp_m1_17_9_r,temp_m1_17_9_i,temp_m1_17_10_r,temp_m1_17_10_i,temp_m1_18_9_r,temp_m1_18_9_i,temp_m1_18_10_r,temp_m1_18_10_i,temp_b1_17_9_r,temp_b1_17_9_i,temp_b1_17_10_r,temp_b1_17_10_i,temp_b1_18_9_r,temp_b1_18_9_i,temp_b1_18_10_r,temp_b1_18_10_i);
MULT MULT134 (clk,in_17_11_r,in_17_11_i,in_17_12_r,in_17_12_i,in_18_11_r,in_18_11_i,in_18_12_r,in_18_12_i,temp_m1_17_11_r,temp_m1_17_11_i,temp_m1_17_12_r,temp_m1_17_12_i,temp_m1_18_11_r,temp_m1_18_11_i,temp_m1_18_12_r,temp_m1_18_12_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly134 (clk,temp_m1_17_11_r,temp_m1_17_11_i,temp_m1_17_12_r,temp_m1_17_12_i,temp_m1_18_11_r,temp_m1_18_11_i,temp_m1_18_12_r,temp_m1_18_12_i,temp_b1_17_11_r,temp_b1_17_11_i,temp_b1_17_12_r,temp_b1_17_12_i,temp_b1_18_11_r,temp_b1_18_11_i,temp_b1_18_12_r,temp_b1_18_12_i);
MULT MULT135 (clk,in_17_13_r,in_17_13_i,in_17_14_r,in_17_14_i,in_18_13_r,in_18_13_i,in_18_14_r,in_18_14_i,temp_m1_17_13_r,temp_m1_17_13_i,temp_m1_17_14_r,temp_m1_17_14_i,temp_m1_18_13_r,temp_m1_18_13_i,temp_m1_18_14_r,temp_m1_18_14_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly135 (clk,temp_m1_17_13_r,temp_m1_17_13_i,temp_m1_17_14_r,temp_m1_17_14_i,temp_m1_18_13_r,temp_m1_18_13_i,temp_m1_18_14_r,temp_m1_18_14_i,temp_b1_17_13_r,temp_b1_17_13_i,temp_b1_17_14_r,temp_b1_17_14_i,temp_b1_18_13_r,temp_b1_18_13_i,temp_b1_18_14_r,temp_b1_18_14_i);
MULT MULT136 (clk,in_17_15_r,in_17_15_i,in_17_16_r,in_17_16_i,in_18_15_r,in_18_15_i,in_18_16_r,in_18_16_i,temp_m1_17_15_r,temp_m1_17_15_i,temp_m1_17_16_r,temp_m1_17_16_i,temp_m1_18_15_r,temp_m1_18_15_i,temp_m1_18_16_r,temp_m1_18_16_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly136 (clk,temp_m1_17_15_r,temp_m1_17_15_i,temp_m1_17_16_r,temp_m1_17_16_i,temp_m1_18_15_r,temp_m1_18_15_i,temp_m1_18_16_r,temp_m1_18_16_i,temp_b1_17_15_r,temp_b1_17_15_i,temp_b1_17_16_r,temp_b1_17_16_i,temp_b1_18_15_r,temp_b1_18_15_i,temp_b1_18_16_r,temp_b1_18_16_i);
MULT MULT137 (clk,in_17_17_r,in_17_17_i,in_17_18_r,in_17_18_i,in_18_17_r,in_18_17_i,in_18_18_r,in_18_18_i,temp_m1_17_17_r,temp_m1_17_17_i,temp_m1_17_18_r,temp_m1_17_18_i,temp_m1_18_17_r,temp_m1_18_17_i,temp_m1_18_18_r,temp_m1_18_18_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly137 (clk,temp_m1_17_17_r,temp_m1_17_17_i,temp_m1_17_18_r,temp_m1_17_18_i,temp_m1_18_17_r,temp_m1_18_17_i,temp_m1_18_18_r,temp_m1_18_18_i,temp_b1_17_17_r,temp_b1_17_17_i,temp_b1_17_18_r,temp_b1_17_18_i,temp_b1_18_17_r,temp_b1_18_17_i,temp_b1_18_18_r,temp_b1_18_18_i);
MULT MULT138 (clk,in_17_19_r,in_17_19_i,in_17_20_r,in_17_20_i,in_18_19_r,in_18_19_i,in_18_20_r,in_18_20_i,temp_m1_17_19_r,temp_m1_17_19_i,temp_m1_17_20_r,temp_m1_17_20_i,temp_m1_18_19_r,temp_m1_18_19_i,temp_m1_18_20_r,temp_m1_18_20_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly138 (clk,temp_m1_17_19_r,temp_m1_17_19_i,temp_m1_17_20_r,temp_m1_17_20_i,temp_m1_18_19_r,temp_m1_18_19_i,temp_m1_18_20_r,temp_m1_18_20_i,temp_b1_17_19_r,temp_b1_17_19_i,temp_b1_17_20_r,temp_b1_17_20_i,temp_b1_18_19_r,temp_b1_18_19_i,temp_b1_18_20_r,temp_b1_18_20_i);
MULT MULT139 (clk,in_17_21_r,in_17_21_i,in_17_22_r,in_17_22_i,in_18_21_r,in_18_21_i,in_18_22_r,in_18_22_i,temp_m1_17_21_r,temp_m1_17_21_i,temp_m1_17_22_r,temp_m1_17_22_i,temp_m1_18_21_r,temp_m1_18_21_i,temp_m1_18_22_r,temp_m1_18_22_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly139 (clk,temp_m1_17_21_r,temp_m1_17_21_i,temp_m1_17_22_r,temp_m1_17_22_i,temp_m1_18_21_r,temp_m1_18_21_i,temp_m1_18_22_r,temp_m1_18_22_i,temp_b1_17_21_r,temp_b1_17_21_i,temp_b1_17_22_r,temp_b1_17_22_i,temp_b1_18_21_r,temp_b1_18_21_i,temp_b1_18_22_r,temp_b1_18_22_i);
MULT MULT140 (clk,in_17_23_r,in_17_23_i,in_17_24_r,in_17_24_i,in_18_23_r,in_18_23_i,in_18_24_r,in_18_24_i,temp_m1_17_23_r,temp_m1_17_23_i,temp_m1_17_24_r,temp_m1_17_24_i,temp_m1_18_23_r,temp_m1_18_23_i,temp_m1_18_24_r,temp_m1_18_24_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly140 (clk,temp_m1_17_23_r,temp_m1_17_23_i,temp_m1_17_24_r,temp_m1_17_24_i,temp_m1_18_23_r,temp_m1_18_23_i,temp_m1_18_24_r,temp_m1_18_24_i,temp_b1_17_23_r,temp_b1_17_23_i,temp_b1_17_24_r,temp_b1_17_24_i,temp_b1_18_23_r,temp_b1_18_23_i,temp_b1_18_24_r,temp_b1_18_24_i);
MULT MULT141 (clk,in_17_25_r,in_17_25_i,in_17_26_r,in_17_26_i,in_18_25_r,in_18_25_i,in_18_26_r,in_18_26_i,temp_m1_17_25_r,temp_m1_17_25_i,temp_m1_17_26_r,temp_m1_17_26_i,temp_m1_18_25_r,temp_m1_18_25_i,temp_m1_18_26_r,temp_m1_18_26_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly141 (clk,temp_m1_17_25_r,temp_m1_17_25_i,temp_m1_17_26_r,temp_m1_17_26_i,temp_m1_18_25_r,temp_m1_18_25_i,temp_m1_18_26_r,temp_m1_18_26_i,temp_b1_17_25_r,temp_b1_17_25_i,temp_b1_17_26_r,temp_b1_17_26_i,temp_b1_18_25_r,temp_b1_18_25_i,temp_b1_18_26_r,temp_b1_18_26_i);
MULT MULT142 (clk,in_17_27_r,in_17_27_i,in_17_28_r,in_17_28_i,in_18_27_r,in_18_27_i,in_18_28_r,in_18_28_i,temp_m1_17_27_r,temp_m1_17_27_i,temp_m1_17_28_r,temp_m1_17_28_i,temp_m1_18_27_r,temp_m1_18_27_i,temp_m1_18_28_r,temp_m1_18_28_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly142 (clk,temp_m1_17_27_r,temp_m1_17_27_i,temp_m1_17_28_r,temp_m1_17_28_i,temp_m1_18_27_r,temp_m1_18_27_i,temp_m1_18_28_r,temp_m1_18_28_i,temp_b1_17_27_r,temp_b1_17_27_i,temp_b1_17_28_r,temp_b1_17_28_i,temp_b1_18_27_r,temp_b1_18_27_i,temp_b1_18_28_r,temp_b1_18_28_i);
MULT MULT143 (clk,in_17_29_r,in_17_29_i,in_17_30_r,in_17_30_i,in_18_29_r,in_18_29_i,in_18_30_r,in_18_30_i,temp_m1_17_29_r,temp_m1_17_29_i,temp_m1_17_30_r,temp_m1_17_30_i,temp_m1_18_29_r,temp_m1_18_29_i,temp_m1_18_30_r,temp_m1_18_30_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly143 (clk,temp_m1_17_29_r,temp_m1_17_29_i,temp_m1_17_30_r,temp_m1_17_30_i,temp_m1_18_29_r,temp_m1_18_29_i,temp_m1_18_30_r,temp_m1_18_30_i,temp_b1_17_29_r,temp_b1_17_29_i,temp_b1_17_30_r,temp_b1_17_30_i,temp_b1_18_29_r,temp_b1_18_29_i,temp_b1_18_30_r,temp_b1_18_30_i);
MULT MULT144 (clk,in_17_31_r,in_17_31_i,in_17_32_r,in_17_32_i,in_18_31_r,in_18_31_i,in_18_32_r,in_18_32_i,temp_m1_17_31_r,temp_m1_17_31_i,temp_m1_17_32_r,temp_m1_17_32_i,temp_m1_18_31_r,temp_m1_18_31_i,temp_m1_18_32_r,temp_m1_18_32_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly144 (clk,temp_m1_17_31_r,temp_m1_17_31_i,temp_m1_17_32_r,temp_m1_17_32_i,temp_m1_18_31_r,temp_m1_18_31_i,temp_m1_18_32_r,temp_m1_18_32_i,temp_b1_17_31_r,temp_b1_17_31_i,temp_b1_17_32_r,temp_b1_17_32_i,temp_b1_18_31_r,temp_b1_18_31_i,temp_b1_18_32_r,temp_b1_18_32_i);
MULT MULT145 (clk,in_19_1_r,in_19_1_i,in_19_2_r,in_19_2_i,in_20_1_r,in_20_1_i,in_20_2_r,in_20_2_i,temp_m1_19_1_r,temp_m1_19_1_i,temp_m1_19_2_r,temp_m1_19_2_i,temp_m1_20_1_r,temp_m1_20_1_i,temp_m1_20_2_r,temp_m1_20_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly145 (clk,temp_m1_19_1_r,temp_m1_19_1_i,temp_m1_19_2_r,temp_m1_19_2_i,temp_m1_20_1_r,temp_m1_20_1_i,temp_m1_20_2_r,temp_m1_20_2_i,temp_b1_19_1_r,temp_b1_19_1_i,temp_b1_19_2_r,temp_b1_19_2_i,temp_b1_20_1_r,temp_b1_20_1_i,temp_b1_20_2_r,temp_b1_20_2_i);
MULT MULT146 (clk,in_19_3_r,in_19_3_i,in_19_4_r,in_19_4_i,in_20_3_r,in_20_3_i,in_20_4_r,in_20_4_i,temp_m1_19_3_r,temp_m1_19_3_i,temp_m1_19_4_r,temp_m1_19_4_i,temp_m1_20_3_r,temp_m1_20_3_i,temp_m1_20_4_r,temp_m1_20_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly146 (clk,temp_m1_19_3_r,temp_m1_19_3_i,temp_m1_19_4_r,temp_m1_19_4_i,temp_m1_20_3_r,temp_m1_20_3_i,temp_m1_20_4_r,temp_m1_20_4_i,temp_b1_19_3_r,temp_b1_19_3_i,temp_b1_19_4_r,temp_b1_19_4_i,temp_b1_20_3_r,temp_b1_20_3_i,temp_b1_20_4_r,temp_b1_20_4_i);
MULT MULT147 (clk,in_19_5_r,in_19_5_i,in_19_6_r,in_19_6_i,in_20_5_r,in_20_5_i,in_20_6_r,in_20_6_i,temp_m1_19_5_r,temp_m1_19_5_i,temp_m1_19_6_r,temp_m1_19_6_i,temp_m1_20_5_r,temp_m1_20_5_i,temp_m1_20_6_r,temp_m1_20_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly147 (clk,temp_m1_19_5_r,temp_m1_19_5_i,temp_m1_19_6_r,temp_m1_19_6_i,temp_m1_20_5_r,temp_m1_20_5_i,temp_m1_20_6_r,temp_m1_20_6_i,temp_b1_19_5_r,temp_b1_19_5_i,temp_b1_19_6_r,temp_b1_19_6_i,temp_b1_20_5_r,temp_b1_20_5_i,temp_b1_20_6_r,temp_b1_20_6_i);
MULT MULT148 (clk,in_19_7_r,in_19_7_i,in_19_8_r,in_19_8_i,in_20_7_r,in_20_7_i,in_20_8_r,in_20_8_i,temp_m1_19_7_r,temp_m1_19_7_i,temp_m1_19_8_r,temp_m1_19_8_i,temp_m1_20_7_r,temp_m1_20_7_i,temp_m1_20_8_r,temp_m1_20_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly148 (clk,temp_m1_19_7_r,temp_m1_19_7_i,temp_m1_19_8_r,temp_m1_19_8_i,temp_m1_20_7_r,temp_m1_20_7_i,temp_m1_20_8_r,temp_m1_20_8_i,temp_b1_19_7_r,temp_b1_19_7_i,temp_b1_19_8_r,temp_b1_19_8_i,temp_b1_20_7_r,temp_b1_20_7_i,temp_b1_20_8_r,temp_b1_20_8_i);
MULT MULT149 (clk,in_19_9_r,in_19_9_i,in_19_10_r,in_19_10_i,in_20_9_r,in_20_9_i,in_20_10_r,in_20_10_i,temp_m1_19_9_r,temp_m1_19_9_i,temp_m1_19_10_r,temp_m1_19_10_i,temp_m1_20_9_r,temp_m1_20_9_i,temp_m1_20_10_r,temp_m1_20_10_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly149 (clk,temp_m1_19_9_r,temp_m1_19_9_i,temp_m1_19_10_r,temp_m1_19_10_i,temp_m1_20_9_r,temp_m1_20_9_i,temp_m1_20_10_r,temp_m1_20_10_i,temp_b1_19_9_r,temp_b1_19_9_i,temp_b1_19_10_r,temp_b1_19_10_i,temp_b1_20_9_r,temp_b1_20_9_i,temp_b1_20_10_r,temp_b1_20_10_i);
MULT MULT150 (clk,in_19_11_r,in_19_11_i,in_19_12_r,in_19_12_i,in_20_11_r,in_20_11_i,in_20_12_r,in_20_12_i,temp_m1_19_11_r,temp_m1_19_11_i,temp_m1_19_12_r,temp_m1_19_12_i,temp_m1_20_11_r,temp_m1_20_11_i,temp_m1_20_12_r,temp_m1_20_12_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly150 (clk,temp_m1_19_11_r,temp_m1_19_11_i,temp_m1_19_12_r,temp_m1_19_12_i,temp_m1_20_11_r,temp_m1_20_11_i,temp_m1_20_12_r,temp_m1_20_12_i,temp_b1_19_11_r,temp_b1_19_11_i,temp_b1_19_12_r,temp_b1_19_12_i,temp_b1_20_11_r,temp_b1_20_11_i,temp_b1_20_12_r,temp_b1_20_12_i);
MULT MULT151 (clk,in_19_13_r,in_19_13_i,in_19_14_r,in_19_14_i,in_20_13_r,in_20_13_i,in_20_14_r,in_20_14_i,temp_m1_19_13_r,temp_m1_19_13_i,temp_m1_19_14_r,temp_m1_19_14_i,temp_m1_20_13_r,temp_m1_20_13_i,temp_m1_20_14_r,temp_m1_20_14_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly151 (clk,temp_m1_19_13_r,temp_m1_19_13_i,temp_m1_19_14_r,temp_m1_19_14_i,temp_m1_20_13_r,temp_m1_20_13_i,temp_m1_20_14_r,temp_m1_20_14_i,temp_b1_19_13_r,temp_b1_19_13_i,temp_b1_19_14_r,temp_b1_19_14_i,temp_b1_20_13_r,temp_b1_20_13_i,temp_b1_20_14_r,temp_b1_20_14_i);
MULT MULT152 (clk,in_19_15_r,in_19_15_i,in_19_16_r,in_19_16_i,in_20_15_r,in_20_15_i,in_20_16_r,in_20_16_i,temp_m1_19_15_r,temp_m1_19_15_i,temp_m1_19_16_r,temp_m1_19_16_i,temp_m1_20_15_r,temp_m1_20_15_i,temp_m1_20_16_r,temp_m1_20_16_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly152 (clk,temp_m1_19_15_r,temp_m1_19_15_i,temp_m1_19_16_r,temp_m1_19_16_i,temp_m1_20_15_r,temp_m1_20_15_i,temp_m1_20_16_r,temp_m1_20_16_i,temp_b1_19_15_r,temp_b1_19_15_i,temp_b1_19_16_r,temp_b1_19_16_i,temp_b1_20_15_r,temp_b1_20_15_i,temp_b1_20_16_r,temp_b1_20_16_i);
MULT MULT153 (clk,in_19_17_r,in_19_17_i,in_19_18_r,in_19_18_i,in_20_17_r,in_20_17_i,in_20_18_r,in_20_18_i,temp_m1_19_17_r,temp_m1_19_17_i,temp_m1_19_18_r,temp_m1_19_18_i,temp_m1_20_17_r,temp_m1_20_17_i,temp_m1_20_18_r,temp_m1_20_18_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly153 (clk,temp_m1_19_17_r,temp_m1_19_17_i,temp_m1_19_18_r,temp_m1_19_18_i,temp_m1_20_17_r,temp_m1_20_17_i,temp_m1_20_18_r,temp_m1_20_18_i,temp_b1_19_17_r,temp_b1_19_17_i,temp_b1_19_18_r,temp_b1_19_18_i,temp_b1_20_17_r,temp_b1_20_17_i,temp_b1_20_18_r,temp_b1_20_18_i);
MULT MULT154 (clk,in_19_19_r,in_19_19_i,in_19_20_r,in_19_20_i,in_20_19_r,in_20_19_i,in_20_20_r,in_20_20_i,temp_m1_19_19_r,temp_m1_19_19_i,temp_m1_19_20_r,temp_m1_19_20_i,temp_m1_20_19_r,temp_m1_20_19_i,temp_m1_20_20_r,temp_m1_20_20_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly154 (clk,temp_m1_19_19_r,temp_m1_19_19_i,temp_m1_19_20_r,temp_m1_19_20_i,temp_m1_20_19_r,temp_m1_20_19_i,temp_m1_20_20_r,temp_m1_20_20_i,temp_b1_19_19_r,temp_b1_19_19_i,temp_b1_19_20_r,temp_b1_19_20_i,temp_b1_20_19_r,temp_b1_20_19_i,temp_b1_20_20_r,temp_b1_20_20_i);
MULT MULT155 (clk,in_19_21_r,in_19_21_i,in_19_22_r,in_19_22_i,in_20_21_r,in_20_21_i,in_20_22_r,in_20_22_i,temp_m1_19_21_r,temp_m1_19_21_i,temp_m1_19_22_r,temp_m1_19_22_i,temp_m1_20_21_r,temp_m1_20_21_i,temp_m1_20_22_r,temp_m1_20_22_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly155 (clk,temp_m1_19_21_r,temp_m1_19_21_i,temp_m1_19_22_r,temp_m1_19_22_i,temp_m1_20_21_r,temp_m1_20_21_i,temp_m1_20_22_r,temp_m1_20_22_i,temp_b1_19_21_r,temp_b1_19_21_i,temp_b1_19_22_r,temp_b1_19_22_i,temp_b1_20_21_r,temp_b1_20_21_i,temp_b1_20_22_r,temp_b1_20_22_i);
MULT MULT156 (clk,in_19_23_r,in_19_23_i,in_19_24_r,in_19_24_i,in_20_23_r,in_20_23_i,in_20_24_r,in_20_24_i,temp_m1_19_23_r,temp_m1_19_23_i,temp_m1_19_24_r,temp_m1_19_24_i,temp_m1_20_23_r,temp_m1_20_23_i,temp_m1_20_24_r,temp_m1_20_24_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly156 (clk,temp_m1_19_23_r,temp_m1_19_23_i,temp_m1_19_24_r,temp_m1_19_24_i,temp_m1_20_23_r,temp_m1_20_23_i,temp_m1_20_24_r,temp_m1_20_24_i,temp_b1_19_23_r,temp_b1_19_23_i,temp_b1_19_24_r,temp_b1_19_24_i,temp_b1_20_23_r,temp_b1_20_23_i,temp_b1_20_24_r,temp_b1_20_24_i);
MULT MULT157 (clk,in_19_25_r,in_19_25_i,in_19_26_r,in_19_26_i,in_20_25_r,in_20_25_i,in_20_26_r,in_20_26_i,temp_m1_19_25_r,temp_m1_19_25_i,temp_m1_19_26_r,temp_m1_19_26_i,temp_m1_20_25_r,temp_m1_20_25_i,temp_m1_20_26_r,temp_m1_20_26_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly157 (clk,temp_m1_19_25_r,temp_m1_19_25_i,temp_m1_19_26_r,temp_m1_19_26_i,temp_m1_20_25_r,temp_m1_20_25_i,temp_m1_20_26_r,temp_m1_20_26_i,temp_b1_19_25_r,temp_b1_19_25_i,temp_b1_19_26_r,temp_b1_19_26_i,temp_b1_20_25_r,temp_b1_20_25_i,temp_b1_20_26_r,temp_b1_20_26_i);
MULT MULT158 (clk,in_19_27_r,in_19_27_i,in_19_28_r,in_19_28_i,in_20_27_r,in_20_27_i,in_20_28_r,in_20_28_i,temp_m1_19_27_r,temp_m1_19_27_i,temp_m1_19_28_r,temp_m1_19_28_i,temp_m1_20_27_r,temp_m1_20_27_i,temp_m1_20_28_r,temp_m1_20_28_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly158 (clk,temp_m1_19_27_r,temp_m1_19_27_i,temp_m1_19_28_r,temp_m1_19_28_i,temp_m1_20_27_r,temp_m1_20_27_i,temp_m1_20_28_r,temp_m1_20_28_i,temp_b1_19_27_r,temp_b1_19_27_i,temp_b1_19_28_r,temp_b1_19_28_i,temp_b1_20_27_r,temp_b1_20_27_i,temp_b1_20_28_r,temp_b1_20_28_i);
MULT MULT159 (clk,in_19_29_r,in_19_29_i,in_19_30_r,in_19_30_i,in_20_29_r,in_20_29_i,in_20_30_r,in_20_30_i,temp_m1_19_29_r,temp_m1_19_29_i,temp_m1_19_30_r,temp_m1_19_30_i,temp_m1_20_29_r,temp_m1_20_29_i,temp_m1_20_30_r,temp_m1_20_30_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly159 (clk,temp_m1_19_29_r,temp_m1_19_29_i,temp_m1_19_30_r,temp_m1_19_30_i,temp_m1_20_29_r,temp_m1_20_29_i,temp_m1_20_30_r,temp_m1_20_30_i,temp_b1_19_29_r,temp_b1_19_29_i,temp_b1_19_30_r,temp_b1_19_30_i,temp_b1_20_29_r,temp_b1_20_29_i,temp_b1_20_30_r,temp_b1_20_30_i);
MULT MULT160 (clk,in_19_31_r,in_19_31_i,in_19_32_r,in_19_32_i,in_20_31_r,in_20_31_i,in_20_32_r,in_20_32_i,temp_m1_19_31_r,temp_m1_19_31_i,temp_m1_19_32_r,temp_m1_19_32_i,temp_m1_20_31_r,temp_m1_20_31_i,temp_m1_20_32_r,temp_m1_20_32_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly160 (clk,temp_m1_19_31_r,temp_m1_19_31_i,temp_m1_19_32_r,temp_m1_19_32_i,temp_m1_20_31_r,temp_m1_20_31_i,temp_m1_20_32_r,temp_m1_20_32_i,temp_b1_19_31_r,temp_b1_19_31_i,temp_b1_19_32_r,temp_b1_19_32_i,temp_b1_20_31_r,temp_b1_20_31_i,temp_b1_20_32_r,temp_b1_20_32_i);
MULT MULT161 (clk,in_21_1_r,in_21_1_i,in_21_2_r,in_21_2_i,in_22_1_r,in_22_1_i,in_22_2_r,in_22_2_i,temp_m1_21_1_r,temp_m1_21_1_i,temp_m1_21_2_r,temp_m1_21_2_i,temp_m1_22_1_r,temp_m1_22_1_i,temp_m1_22_2_r,temp_m1_22_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly161 (clk,temp_m1_21_1_r,temp_m1_21_1_i,temp_m1_21_2_r,temp_m1_21_2_i,temp_m1_22_1_r,temp_m1_22_1_i,temp_m1_22_2_r,temp_m1_22_2_i,temp_b1_21_1_r,temp_b1_21_1_i,temp_b1_21_2_r,temp_b1_21_2_i,temp_b1_22_1_r,temp_b1_22_1_i,temp_b1_22_2_r,temp_b1_22_2_i);
MULT MULT162 (clk,in_21_3_r,in_21_3_i,in_21_4_r,in_21_4_i,in_22_3_r,in_22_3_i,in_22_4_r,in_22_4_i,temp_m1_21_3_r,temp_m1_21_3_i,temp_m1_21_4_r,temp_m1_21_4_i,temp_m1_22_3_r,temp_m1_22_3_i,temp_m1_22_4_r,temp_m1_22_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly162 (clk,temp_m1_21_3_r,temp_m1_21_3_i,temp_m1_21_4_r,temp_m1_21_4_i,temp_m1_22_3_r,temp_m1_22_3_i,temp_m1_22_4_r,temp_m1_22_4_i,temp_b1_21_3_r,temp_b1_21_3_i,temp_b1_21_4_r,temp_b1_21_4_i,temp_b1_22_3_r,temp_b1_22_3_i,temp_b1_22_4_r,temp_b1_22_4_i);
MULT MULT163 (clk,in_21_5_r,in_21_5_i,in_21_6_r,in_21_6_i,in_22_5_r,in_22_5_i,in_22_6_r,in_22_6_i,temp_m1_21_5_r,temp_m1_21_5_i,temp_m1_21_6_r,temp_m1_21_6_i,temp_m1_22_5_r,temp_m1_22_5_i,temp_m1_22_6_r,temp_m1_22_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly163 (clk,temp_m1_21_5_r,temp_m1_21_5_i,temp_m1_21_6_r,temp_m1_21_6_i,temp_m1_22_5_r,temp_m1_22_5_i,temp_m1_22_6_r,temp_m1_22_6_i,temp_b1_21_5_r,temp_b1_21_5_i,temp_b1_21_6_r,temp_b1_21_6_i,temp_b1_22_5_r,temp_b1_22_5_i,temp_b1_22_6_r,temp_b1_22_6_i);
MULT MULT164 (clk,in_21_7_r,in_21_7_i,in_21_8_r,in_21_8_i,in_22_7_r,in_22_7_i,in_22_8_r,in_22_8_i,temp_m1_21_7_r,temp_m1_21_7_i,temp_m1_21_8_r,temp_m1_21_8_i,temp_m1_22_7_r,temp_m1_22_7_i,temp_m1_22_8_r,temp_m1_22_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly164 (clk,temp_m1_21_7_r,temp_m1_21_7_i,temp_m1_21_8_r,temp_m1_21_8_i,temp_m1_22_7_r,temp_m1_22_7_i,temp_m1_22_8_r,temp_m1_22_8_i,temp_b1_21_7_r,temp_b1_21_7_i,temp_b1_21_8_r,temp_b1_21_8_i,temp_b1_22_7_r,temp_b1_22_7_i,temp_b1_22_8_r,temp_b1_22_8_i);
MULT MULT165 (clk,in_21_9_r,in_21_9_i,in_21_10_r,in_21_10_i,in_22_9_r,in_22_9_i,in_22_10_r,in_22_10_i,temp_m1_21_9_r,temp_m1_21_9_i,temp_m1_21_10_r,temp_m1_21_10_i,temp_m1_22_9_r,temp_m1_22_9_i,temp_m1_22_10_r,temp_m1_22_10_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly165 (clk,temp_m1_21_9_r,temp_m1_21_9_i,temp_m1_21_10_r,temp_m1_21_10_i,temp_m1_22_9_r,temp_m1_22_9_i,temp_m1_22_10_r,temp_m1_22_10_i,temp_b1_21_9_r,temp_b1_21_9_i,temp_b1_21_10_r,temp_b1_21_10_i,temp_b1_22_9_r,temp_b1_22_9_i,temp_b1_22_10_r,temp_b1_22_10_i);
MULT MULT166 (clk,in_21_11_r,in_21_11_i,in_21_12_r,in_21_12_i,in_22_11_r,in_22_11_i,in_22_12_r,in_22_12_i,temp_m1_21_11_r,temp_m1_21_11_i,temp_m1_21_12_r,temp_m1_21_12_i,temp_m1_22_11_r,temp_m1_22_11_i,temp_m1_22_12_r,temp_m1_22_12_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly166 (clk,temp_m1_21_11_r,temp_m1_21_11_i,temp_m1_21_12_r,temp_m1_21_12_i,temp_m1_22_11_r,temp_m1_22_11_i,temp_m1_22_12_r,temp_m1_22_12_i,temp_b1_21_11_r,temp_b1_21_11_i,temp_b1_21_12_r,temp_b1_21_12_i,temp_b1_22_11_r,temp_b1_22_11_i,temp_b1_22_12_r,temp_b1_22_12_i);
MULT MULT167 (clk,in_21_13_r,in_21_13_i,in_21_14_r,in_21_14_i,in_22_13_r,in_22_13_i,in_22_14_r,in_22_14_i,temp_m1_21_13_r,temp_m1_21_13_i,temp_m1_21_14_r,temp_m1_21_14_i,temp_m1_22_13_r,temp_m1_22_13_i,temp_m1_22_14_r,temp_m1_22_14_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly167 (clk,temp_m1_21_13_r,temp_m1_21_13_i,temp_m1_21_14_r,temp_m1_21_14_i,temp_m1_22_13_r,temp_m1_22_13_i,temp_m1_22_14_r,temp_m1_22_14_i,temp_b1_21_13_r,temp_b1_21_13_i,temp_b1_21_14_r,temp_b1_21_14_i,temp_b1_22_13_r,temp_b1_22_13_i,temp_b1_22_14_r,temp_b1_22_14_i);
MULT MULT168 (clk,in_21_15_r,in_21_15_i,in_21_16_r,in_21_16_i,in_22_15_r,in_22_15_i,in_22_16_r,in_22_16_i,temp_m1_21_15_r,temp_m1_21_15_i,temp_m1_21_16_r,temp_m1_21_16_i,temp_m1_22_15_r,temp_m1_22_15_i,temp_m1_22_16_r,temp_m1_22_16_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly168 (clk,temp_m1_21_15_r,temp_m1_21_15_i,temp_m1_21_16_r,temp_m1_21_16_i,temp_m1_22_15_r,temp_m1_22_15_i,temp_m1_22_16_r,temp_m1_22_16_i,temp_b1_21_15_r,temp_b1_21_15_i,temp_b1_21_16_r,temp_b1_21_16_i,temp_b1_22_15_r,temp_b1_22_15_i,temp_b1_22_16_r,temp_b1_22_16_i);
MULT MULT169 (clk,in_21_17_r,in_21_17_i,in_21_18_r,in_21_18_i,in_22_17_r,in_22_17_i,in_22_18_r,in_22_18_i,temp_m1_21_17_r,temp_m1_21_17_i,temp_m1_21_18_r,temp_m1_21_18_i,temp_m1_22_17_r,temp_m1_22_17_i,temp_m1_22_18_r,temp_m1_22_18_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly169 (clk,temp_m1_21_17_r,temp_m1_21_17_i,temp_m1_21_18_r,temp_m1_21_18_i,temp_m1_22_17_r,temp_m1_22_17_i,temp_m1_22_18_r,temp_m1_22_18_i,temp_b1_21_17_r,temp_b1_21_17_i,temp_b1_21_18_r,temp_b1_21_18_i,temp_b1_22_17_r,temp_b1_22_17_i,temp_b1_22_18_r,temp_b1_22_18_i);
MULT MULT170 (clk,in_21_19_r,in_21_19_i,in_21_20_r,in_21_20_i,in_22_19_r,in_22_19_i,in_22_20_r,in_22_20_i,temp_m1_21_19_r,temp_m1_21_19_i,temp_m1_21_20_r,temp_m1_21_20_i,temp_m1_22_19_r,temp_m1_22_19_i,temp_m1_22_20_r,temp_m1_22_20_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly170 (clk,temp_m1_21_19_r,temp_m1_21_19_i,temp_m1_21_20_r,temp_m1_21_20_i,temp_m1_22_19_r,temp_m1_22_19_i,temp_m1_22_20_r,temp_m1_22_20_i,temp_b1_21_19_r,temp_b1_21_19_i,temp_b1_21_20_r,temp_b1_21_20_i,temp_b1_22_19_r,temp_b1_22_19_i,temp_b1_22_20_r,temp_b1_22_20_i);
MULT MULT171 (clk,in_21_21_r,in_21_21_i,in_21_22_r,in_21_22_i,in_22_21_r,in_22_21_i,in_22_22_r,in_22_22_i,temp_m1_21_21_r,temp_m1_21_21_i,temp_m1_21_22_r,temp_m1_21_22_i,temp_m1_22_21_r,temp_m1_22_21_i,temp_m1_22_22_r,temp_m1_22_22_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly171 (clk,temp_m1_21_21_r,temp_m1_21_21_i,temp_m1_21_22_r,temp_m1_21_22_i,temp_m1_22_21_r,temp_m1_22_21_i,temp_m1_22_22_r,temp_m1_22_22_i,temp_b1_21_21_r,temp_b1_21_21_i,temp_b1_21_22_r,temp_b1_21_22_i,temp_b1_22_21_r,temp_b1_22_21_i,temp_b1_22_22_r,temp_b1_22_22_i);
MULT MULT172 (clk,in_21_23_r,in_21_23_i,in_21_24_r,in_21_24_i,in_22_23_r,in_22_23_i,in_22_24_r,in_22_24_i,temp_m1_21_23_r,temp_m1_21_23_i,temp_m1_21_24_r,temp_m1_21_24_i,temp_m1_22_23_r,temp_m1_22_23_i,temp_m1_22_24_r,temp_m1_22_24_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly172 (clk,temp_m1_21_23_r,temp_m1_21_23_i,temp_m1_21_24_r,temp_m1_21_24_i,temp_m1_22_23_r,temp_m1_22_23_i,temp_m1_22_24_r,temp_m1_22_24_i,temp_b1_21_23_r,temp_b1_21_23_i,temp_b1_21_24_r,temp_b1_21_24_i,temp_b1_22_23_r,temp_b1_22_23_i,temp_b1_22_24_r,temp_b1_22_24_i);
MULT MULT173 (clk,in_21_25_r,in_21_25_i,in_21_26_r,in_21_26_i,in_22_25_r,in_22_25_i,in_22_26_r,in_22_26_i,temp_m1_21_25_r,temp_m1_21_25_i,temp_m1_21_26_r,temp_m1_21_26_i,temp_m1_22_25_r,temp_m1_22_25_i,temp_m1_22_26_r,temp_m1_22_26_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly173 (clk,temp_m1_21_25_r,temp_m1_21_25_i,temp_m1_21_26_r,temp_m1_21_26_i,temp_m1_22_25_r,temp_m1_22_25_i,temp_m1_22_26_r,temp_m1_22_26_i,temp_b1_21_25_r,temp_b1_21_25_i,temp_b1_21_26_r,temp_b1_21_26_i,temp_b1_22_25_r,temp_b1_22_25_i,temp_b1_22_26_r,temp_b1_22_26_i);
MULT MULT174 (clk,in_21_27_r,in_21_27_i,in_21_28_r,in_21_28_i,in_22_27_r,in_22_27_i,in_22_28_r,in_22_28_i,temp_m1_21_27_r,temp_m1_21_27_i,temp_m1_21_28_r,temp_m1_21_28_i,temp_m1_22_27_r,temp_m1_22_27_i,temp_m1_22_28_r,temp_m1_22_28_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly174 (clk,temp_m1_21_27_r,temp_m1_21_27_i,temp_m1_21_28_r,temp_m1_21_28_i,temp_m1_22_27_r,temp_m1_22_27_i,temp_m1_22_28_r,temp_m1_22_28_i,temp_b1_21_27_r,temp_b1_21_27_i,temp_b1_21_28_r,temp_b1_21_28_i,temp_b1_22_27_r,temp_b1_22_27_i,temp_b1_22_28_r,temp_b1_22_28_i);
MULT MULT175 (clk,in_21_29_r,in_21_29_i,in_21_30_r,in_21_30_i,in_22_29_r,in_22_29_i,in_22_30_r,in_22_30_i,temp_m1_21_29_r,temp_m1_21_29_i,temp_m1_21_30_r,temp_m1_21_30_i,temp_m1_22_29_r,temp_m1_22_29_i,temp_m1_22_30_r,temp_m1_22_30_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly175 (clk,temp_m1_21_29_r,temp_m1_21_29_i,temp_m1_21_30_r,temp_m1_21_30_i,temp_m1_22_29_r,temp_m1_22_29_i,temp_m1_22_30_r,temp_m1_22_30_i,temp_b1_21_29_r,temp_b1_21_29_i,temp_b1_21_30_r,temp_b1_21_30_i,temp_b1_22_29_r,temp_b1_22_29_i,temp_b1_22_30_r,temp_b1_22_30_i);
MULT MULT176 (clk,in_21_31_r,in_21_31_i,in_21_32_r,in_21_32_i,in_22_31_r,in_22_31_i,in_22_32_r,in_22_32_i,temp_m1_21_31_r,temp_m1_21_31_i,temp_m1_21_32_r,temp_m1_21_32_i,temp_m1_22_31_r,temp_m1_22_31_i,temp_m1_22_32_r,temp_m1_22_32_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly176 (clk,temp_m1_21_31_r,temp_m1_21_31_i,temp_m1_21_32_r,temp_m1_21_32_i,temp_m1_22_31_r,temp_m1_22_31_i,temp_m1_22_32_r,temp_m1_22_32_i,temp_b1_21_31_r,temp_b1_21_31_i,temp_b1_21_32_r,temp_b1_21_32_i,temp_b1_22_31_r,temp_b1_22_31_i,temp_b1_22_32_r,temp_b1_22_32_i);
MULT MULT177 (clk,in_23_1_r,in_23_1_i,in_23_2_r,in_23_2_i,in_24_1_r,in_24_1_i,in_24_2_r,in_24_2_i,temp_m1_23_1_r,temp_m1_23_1_i,temp_m1_23_2_r,temp_m1_23_2_i,temp_m1_24_1_r,temp_m1_24_1_i,temp_m1_24_2_r,temp_m1_24_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly177 (clk,temp_m1_23_1_r,temp_m1_23_1_i,temp_m1_23_2_r,temp_m1_23_2_i,temp_m1_24_1_r,temp_m1_24_1_i,temp_m1_24_2_r,temp_m1_24_2_i,temp_b1_23_1_r,temp_b1_23_1_i,temp_b1_23_2_r,temp_b1_23_2_i,temp_b1_24_1_r,temp_b1_24_1_i,temp_b1_24_2_r,temp_b1_24_2_i);
MULT MULT178 (clk,in_23_3_r,in_23_3_i,in_23_4_r,in_23_4_i,in_24_3_r,in_24_3_i,in_24_4_r,in_24_4_i,temp_m1_23_3_r,temp_m1_23_3_i,temp_m1_23_4_r,temp_m1_23_4_i,temp_m1_24_3_r,temp_m1_24_3_i,temp_m1_24_4_r,temp_m1_24_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly178 (clk,temp_m1_23_3_r,temp_m1_23_3_i,temp_m1_23_4_r,temp_m1_23_4_i,temp_m1_24_3_r,temp_m1_24_3_i,temp_m1_24_4_r,temp_m1_24_4_i,temp_b1_23_3_r,temp_b1_23_3_i,temp_b1_23_4_r,temp_b1_23_4_i,temp_b1_24_3_r,temp_b1_24_3_i,temp_b1_24_4_r,temp_b1_24_4_i);
MULT MULT179 (clk,in_23_5_r,in_23_5_i,in_23_6_r,in_23_6_i,in_24_5_r,in_24_5_i,in_24_6_r,in_24_6_i,temp_m1_23_5_r,temp_m1_23_5_i,temp_m1_23_6_r,temp_m1_23_6_i,temp_m1_24_5_r,temp_m1_24_5_i,temp_m1_24_6_r,temp_m1_24_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly179 (clk,temp_m1_23_5_r,temp_m1_23_5_i,temp_m1_23_6_r,temp_m1_23_6_i,temp_m1_24_5_r,temp_m1_24_5_i,temp_m1_24_6_r,temp_m1_24_6_i,temp_b1_23_5_r,temp_b1_23_5_i,temp_b1_23_6_r,temp_b1_23_6_i,temp_b1_24_5_r,temp_b1_24_5_i,temp_b1_24_6_r,temp_b1_24_6_i);
MULT MULT180 (clk,in_23_7_r,in_23_7_i,in_23_8_r,in_23_8_i,in_24_7_r,in_24_7_i,in_24_8_r,in_24_8_i,temp_m1_23_7_r,temp_m1_23_7_i,temp_m1_23_8_r,temp_m1_23_8_i,temp_m1_24_7_r,temp_m1_24_7_i,temp_m1_24_8_r,temp_m1_24_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly180 (clk,temp_m1_23_7_r,temp_m1_23_7_i,temp_m1_23_8_r,temp_m1_23_8_i,temp_m1_24_7_r,temp_m1_24_7_i,temp_m1_24_8_r,temp_m1_24_8_i,temp_b1_23_7_r,temp_b1_23_7_i,temp_b1_23_8_r,temp_b1_23_8_i,temp_b1_24_7_r,temp_b1_24_7_i,temp_b1_24_8_r,temp_b1_24_8_i);
MULT MULT181 (clk,in_23_9_r,in_23_9_i,in_23_10_r,in_23_10_i,in_24_9_r,in_24_9_i,in_24_10_r,in_24_10_i,temp_m1_23_9_r,temp_m1_23_9_i,temp_m1_23_10_r,temp_m1_23_10_i,temp_m1_24_9_r,temp_m1_24_9_i,temp_m1_24_10_r,temp_m1_24_10_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly181 (clk,temp_m1_23_9_r,temp_m1_23_9_i,temp_m1_23_10_r,temp_m1_23_10_i,temp_m1_24_9_r,temp_m1_24_9_i,temp_m1_24_10_r,temp_m1_24_10_i,temp_b1_23_9_r,temp_b1_23_9_i,temp_b1_23_10_r,temp_b1_23_10_i,temp_b1_24_9_r,temp_b1_24_9_i,temp_b1_24_10_r,temp_b1_24_10_i);
MULT MULT182 (clk,in_23_11_r,in_23_11_i,in_23_12_r,in_23_12_i,in_24_11_r,in_24_11_i,in_24_12_r,in_24_12_i,temp_m1_23_11_r,temp_m1_23_11_i,temp_m1_23_12_r,temp_m1_23_12_i,temp_m1_24_11_r,temp_m1_24_11_i,temp_m1_24_12_r,temp_m1_24_12_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly182 (clk,temp_m1_23_11_r,temp_m1_23_11_i,temp_m1_23_12_r,temp_m1_23_12_i,temp_m1_24_11_r,temp_m1_24_11_i,temp_m1_24_12_r,temp_m1_24_12_i,temp_b1_23_11_r,temp_b1_23_11_i,temp_b1_23_12_r,temp_b1_23_12_i,temp_b1_24_11_r,temp_b1_24_11_i,temp_b1_24_12_r,temp_b1_24_12_i);
MULT MULT183 (clk,in_23_13_r,in_23_13_i,in_23_14_r,in_23_14_i,in_24_13_r,in_24_13_i,in_24_14_r,in_24_14_i,temp_m1_23_13_r,temp_m1_23_13_i,temp_m1_23_14_r,temp_m1_23_14_i,temp_m1_24_13_r,temp_m1_24_13_i,temp_m1_24_14_r,temp_m1_24_14_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly183 (clk,temp_m1_23_13_r,temp_m1_23_13_i,temp_m1_23_14_r,temp_m1_23_14_i,temp_m1_24_13_r,temp_m1_24_13_i,temp_m1_24_14_r,temp_m1_24_14_i,temp_b1_23_13_r,temp_b1_23_13_i,temp_b1_23_14_r,temp_b1_23_14_i,temp_b1_24_13_r,temp_b1_24_13_i,temp_b1_24_14_r,temp_b1_24_14_i);
MULT MULT184 (clk,in_23_15_r,in_23_15_i,in_23_16_r,in_23_16_i,in_24_15_r,in_24_15_i,in_24_16_r,in_24_16_i,temp_m1_23_15_r,temp_m1_23_15_i,temp_m1_23_16_r,temp_m1_23_16_i,temp_m1_24_15_r,temp_m1_24_15_i,temp_m1_24_16_r,temp_m1_24_16_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly184 (clk,temp_m1_23_15_r,temp_m1_23_15_i,temp_m1_23_16_r,temp_m1_23_16_i,temp_m1_24_15_r,temp_m1_24_15_i,temp_m1_24_16_r,temp_m1_24_16_i,temp_b1_23_15_r,temp_b1_23_15_i,temp_b1_23_16_r,temp_b1_23_16_i,temp_b1_24_15_r,temp_b1_24_15_i,temp_b1_24_16_r,temp_b1_24_16_i);
MULT MULT185 (clk,in_23_17_r,in_23_17_i,in_23_18_r,in_23_18_i,in_24_17_r,in_24_17_i,in_24_18_r,in_24_18_i,temp_m1_23_17_r,temp_m1_23_17_i,temp_m1_23_18_r,temp_m1_23_18_i,temp_m1_24_17_r,temp_m1_24_17_i,temp_m1_24_18_r,temp_m1_24_18_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly185 (clk,temp_m1_23_17_r,temp_m1_23_17_i,temp_m1_23_18_r,temp_m1_23_18_i,temp_m1_24_17_r,temp_m1_24_17_i,temp_m1_24_18_r,temp_m1_24_18_i,temp_b1_23_17_r,temp_b1_23_17_i,temp_b1_23_18_r,temp_b1_23_18_i,temp_b1_24_17_r,temp_b1_24_17_i,temp_b1_24_18_r,temp_b1_24_18_i);
MULT MULT186 (clk,in_23_19_r,in_23_19_i,in_23_20_r,in_23_20_i,in_24_19_r,in_24_19_i,in_24_20_r,in_24_20_i,temp_m1_23_19_r,temp_m1_23_19_i,temp_m1_23_20_r,temp_m1_23_20_i,temp_m1_24_19_r,temp_m1_24_19_i,temp_m1_24_20_r,temp_m1_24_20_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly186 (clk,temp_m1_23_19_r,temp_m1_23_19_i,temp_m1_23_20_r,temp_m1_23_20_i,temp_m1_24_19_r,temp_m1_24_19_i,temp_m1_24_20_r,temp_m1_24_20_i,temp_b1_23_19_r,temp_b1_23_19_i,temp_b1_23_20_r,temp_b1_23_20_i,temp_b1_24_19_r,temp_b1_24_19_i,temp_b1_24_20_r,temp_b1_24_20_i);
MULT MULT187 (clk,in_23_21_r,in_23_21_i,in_23_22_r,in_23_22_i,in_24_21_r,in_24_21_i,in_24_22_r,in_24_22_i,temp_m1_23_21_r,temp_m1_23_21_i,temp_m1_23_22_r,temp_m1_23_22_i,temp_m1_24_21_r,temp_m1_24_21_i,temp_m1_24_22_r,temp_m1_24_22_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly187 (clk,temp_m1_23_21_r,temp_m1_23_21_i,temp_m1_23_22_r,temp_m1_23_22_i,temp_m1_24_21_r,temp_m1_24_21_i,temp_m1_24_22_r,temp_m1_24_22_i,temp_b1_23_21_r,temp_b1_23_21_i,temp_b1_23_22_r,temp_b1_23_22_i,temp_b1_24_21_r,temp_b1_24_21_i,temp_b1_24_22_r,temp_b1_24_22_i);
MULT MULT188 (clk,in_23_23_r,in_23_23_i,in_23_24_r,in_23_24_i,in_24_23_r,in_24_23_i,in_24_24_r,in_24_24_i,temp_m1_23_23_r,temp_m1_23_23_i,temp_m1_23_24_r,temp_m1_23_24_i,temp_m1_24_23_r,temp_m1_24_23_i,temp_m1_24_24_r,temp_m1_24_24_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly188 (clk,temp_m1_23_23_r,temp_m1_23_23_i,temp_m1_23_24_r,temp_m1_23_24_i,temp_m1_24_23_r,temp_m1_24_23_i,temp_m1_24_24_r,temp_m1_24_24_i,temp_b1_23_23_r,temp_b1_23_23_i,temp_b1_23_24_r,temp_b1_23_24_i,temp_b1_24_23_r,temp_b1_24_23_i,temp_b1_24_24_r,temp_b1_24_24_i);
MULT MULT189 (clk,in_23_25_r,in_23_25_i,in_23_26_r,in_23_26_i,in_24_25_r,in_24_25_i,in_24_26_r,in_24_26_i,temp_m1_23_25_r,temp_m1_23_25_i,temp_m1_23_26_r,temp_m1_23_26_i,temp_m1_24_25_r,temp_m1_24_25_i,temp_m1_24_26_r,temp_m1_24_26_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly189 (clk,temp_m1_23_25_r,temp_m1_23_25_i,temp_m1_23_26_r,temp_m1_23_26_i,temp_m1_24_25_r,temp_m1_24_25_i,temp_m1_24_26_r,temp_m1_24_26_i,temp_b1_23_25_r,temp_b1_23_25_i,temp_b1_23_26_r,temp_b1_23_26_i,temp_b1_24_25_r,temp_b1_24_25_i,temp_b1_24_26_r,temp_b1_24_26_i);
MULT MULT190 (clk,in_23_27_r,in_23_27_i,in_23_28_r,in_23_28_i,in_24_27_r,in_24_27_i,in_24_28_r,in_24_28_i,temp_m1_23_27_r,temp_m1_23_27_i,temp_m1_23_28_r,temp_m1_23_28_i,temp_m1_24_27_r,temp_m1_24_27_i,temp_m1_24_28_r,temp_m1_24_28_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly190 (clk,temp_m1_23_27_r,temp_m1_23_27_i,temp_m1_23_28_r,temp_m1_23_28_i,temp_m1_24_27_r,temp_m1_24_27_i,temp_m1_24_28_r,temp_m1_24_28_i,temp_b1_23_27_r,temp_b1_23_27_i,temp_b1_23_28_r,temp_b1_23_28_i,temp_b1_24_27_r,temp_b1_24_27_i,temp_b1_24_28_r,temp_b1_24_28_i);
MULT MULT191 (clk,in_23_29_r,in_23_29_i,in_23_30_r,in_23_30_i,in_24_29_r,in_24_29_i,in_24_30_r,in_24_30_i,temp_m1_23_29_r,temp_m1_23_29_i,temp_m1_23_30_r,temp_m1_23_30_i,temp_m1_24_29_r,temp_m1_24_29_i,temp_m1_24_30_r,temp_m1_24_30_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly191 (clk,temp_m1_23_29_r,temp_m1_23_29_i,temp_m1_23_30_r,temp_m1_23_30_i,temp_m1_24_29_r,temp_m1_24_29_i,temp_m1_24_30_r,temp_m1_24_30_i,temp_b1_23_29_r,temp_b1_23_29_i,temp_b1_23_30_r,temp_b1_23_30_i,temp_b1_24_29_r,temp_b1_24_29_i,temp_b1_24_30_r,temp_b1_24_30_i);
MULT MULT192 (clk,in_23_31_r,in_23_31_i,in_23_32_r,in_23_32_i,in_24_31_r,in_24_31_i,in_24_32_r,in_24_32_i,temp_m1_23_31_r,temp_m1_23_31_i,temp_m1_23_32_r,temp_m1_23_32_i,temp_m1_24_31_r,temp_m1_24_31_i,temp_m1_24_32_r,temp_m1_24_32_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly192 (clk,temp_m1_23_31_r,temp_m1_23_31_i,temp_m1_23_32_r,temp_m1_23_32_i,temp_m1_24_31_r,temp_m1_24_31_i,temp_m1_24_32_r,temp_m1_24_32_i,temp_b1_23_31_r,temp_b1_23_31_i,temp_b1_23_32_r,temp_b1_23_32_i,temp_b1_24_31_r,temp_b1_24_31_i,temp_b1_24_32_r,temp_b1_24_32_i);
MULT MULT193 (clk,in_25_1_r,in_25_1_i,in_25_2_r,in_25_2_i,in_26_1_r,in_26_1_i,in_26_2_r,in_26_2_i,temp_m1_25_1_r,temp_m1_25_1_i,temp_m1_25_2_r,temp_m1_25_2_i,temp_m1_26_1_r,temp_m1_26_1_i,temp_m1_26_2_r,temp_m1_26_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly193 (clk,temp_m1_25_1_r,temp_m1_25_1_i,temp_m1_25_2_r,temp_m1_25_2_i,temp_m1_26_1_r,temp_m1_26_1_i,temp_m1_26_2_r,temp_m1_26_2_i,temp_b1_25_1_r,temp_b1_25_1_i,temp_b1_25_2_r,temp_b1_25_2_i,temp_b1_26_1_r,temp_b1_26_1_i,temp_b1_26_2_r,temp_b1_26_2_i);
MULT MULT194 (clk,in_25_3_r,in_25_3_i,in_25_4_r,in_25_4_i,in_26_3_r,in_26_3_i,in_26_4_r,in_26_4_i,temp_m1_25_3_r,temp_m1_25_3_i,temp_m1_25_4_r,temp_m1_25_4_i,temp_m1_26_3_r,temp_m1_26_3_i,temp_m1_26_4_r,temp_m1_26_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly194 (clk,temp_m1_25_3_r,temp_m1_25_3_i,temp_m1_25_4_r,temp_m1_25_4_i,temp_m1_26_3_r,temp_m1_26_3_i,temp_m1_26_4_r,temp_m1_26_4_i,temp_b1_25_3_r,temp_b1_25_3_i,temp_b1_25_4_r,temp_b1_25_4_i,temp_b1_26_3_r,temp_b1_26_3_i,temp_b1_26_4_r,temp_b1_26_4_i);
MULT MULT195 (clk,in_25_5_r,in_25_5_i,in_25_6_r,in_25_6_i,in_26_5_r,in_26_5_i,in_26_6_r,in_26_6_i,temp_m1_25_5_r,temp_m1_25_5_i,temp_m1_25_6_r,temp_m1_25_6_i,temp_m1_26_5_r,temp_m1_26_5_i,temp_m1_26_6_r,temp_m1_26_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly195 (clk,temp_m1_25_5_r,temp_m1_25_5_i,temp_m1_25_6_r,temp_m1_25_6_i,temp_m1_26_5_r,temp_m1_26_5_i,temp_m1_26_6_r,temp_m1_26_6_i,temp_b1_25_5_r,temp_b1_25_5_i,temp_b1_25_6_r,temp_b1_25_6_i,temp_b1_26_5_r,temp_b1_26_5_i,temp_b1_26_6_r,temp_b1_26_6_i);
MULT MULT196 (clk,in_25_7_r,in_25_7_i,in_25_8_r,in_25_8_i,in_26_7_r,in_26_7_i,in_26_8_r,in_26_8_i,temp_m1_25_7_r,temp_m1_25_7_i,temp_m1_25_8_r,temp_m1_25_8_i,temp_m1_26_7_r,temp_m1_26_7_i,temp_m1_26_8_r,temp_m1_26_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly196 (clk,temp_m1_25_7_r,temp_m1_25_7_i,temp_m1_25_8_r,temp_m1_25_8_i,temp_m1_26_7_r,temp_m1_26_7_i,temp_m1_26_8_r,temp_m1_26_8_i,temp_b1_25_7_r,temp_b1_25_7_i,temp_b1_25_8_r,temp_b1_25_8_i,temp_b1_26_7_r,temp_b1_26_7_i,temp_b1_26_8_r,temp_b1_26_8_i);
MULT MULT197 (clk,in_25_9_r,in_25_9_i,in_25_10_r,in_25_10_i,in_26_9_r,in_26_9_i,in_26_10_r,in_26_10_i,temp_m1_25_9_r,temp_m1_25_9_i,temp_m1_25_10_r,temp_m1_25_10_i,temp_m1_26_9_r,temp_m1_26_9_i,temp_m1_26_10_r,temp_m1_26_10_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly197 (clk,temp_m1_25_9_r,temp_m1_25_9_i,temp_m1_25_10_r,temp_m1_25_10_i,temp_m1_26_9_r,temp_m1_26_9_i,temp_m1_26_10_r,temp_m1_26_10_i,temp_b1_25_9_r,temp_b1_25_9_i,temp_b1_25_10_r,temp_b1_25_10_i,temp_b1_26_9_r,temp_b1_26_9_i,temp_b1_26_10_r,temp_b1_26_10_i);
MULT MULT198 (clk,in_25_11_r,in_25_11_i,in_25_12_r,in_25_12_i,in_26_11_r,in_26_11_i,in_26_12_r,in_26_12_i,temp_m1_25_11_r,temp_m1_25_11_i,temp_m1_25_12_r,temp_m1_25_12_i,temp_m1_26_11_r,temp_m1_26_11_i,temp_m1_26_12_r,temp_m1_26_12_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly198 (clk,temp_m1_25_11_r,temp_m1_25_11_i,temp_m1_25_12_r,temp_m1_25_12_i,temp_m1_26_11_r,temp_m1_26_11_i,temp_m1_26_12_r,temp_m1_26_12_i,temp_b1_25_11_r,temp_b1_25_11_i,temp_b1_25_12_r,temp_b1_25_12_i,temp_b1_26_11_r,temp_b1_26_11_i,temp_b1_26_12_r,temp_b1_26_12_i);
MULT MULT199 (clk,in_25_13_r,in_25_13_i,in_25_14_r,in_25_14_i,in_26_13_r,in_26_13_i,in_26_14_r,in_26_14_i,temp_m1_25_13_r,temp_m1_25_13_i,temp_m1_25_14_r,temp_m1_25_14_i,temp_m1_26_13_r,temp_m1_26_13_i,temp_m1_26_14_r,temp_m1_26_14_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly199 (clk,temp_m1_25_13_r,temp_m1_25_13_i,temp_m1_25_14_r,temp_m1_25_14_i,temp_m1_26_13_r,temp_m1_26_13_i,temp_m1_26_14_r,temp_m1_26_14_i,temp_b1_25_13_r,temp_b1_25_13_i,temp_b1_25_14_r,temp_b1_25_14_i,temp_b1_26_13_r,temp_b1_26_13_i,temp_b1_26_14_r,temp_b1_26_14_i);
MULT MULT200 (clk,in_25_15_r,in_25_15_i,in_25_16_r,in_25_16_i,in_26_15_r,in_26_15_i,in_26_16_r,in_26_16_i,temp_m1_25_15_r,temp_m1_25_15_i,temp_m1_25_16_r,temp_m1_25_16_i,temp_m1_26_15_r,temp_m1_26_15_i,temp_m1_26_16_r,temp_m1_26_16_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly200 (clk,temp_m1_25_15_r,temp_m1_25_15_i,temp_m1_25_16_r,temp_m1_25_16_i,temp_m1_26_15_r,temp_m1_26_15_i,temp_m1_26_16_r,temp_m1_26_16_i,temp_b1_25_15_r,temp_b1_25_15_i,temp_b1_25_16_r,temp_b1_25_16_i,temp_b1_26_15_r,temp_b1_26_15_i,temp_b1_26_16_r,temp_b1_26_16_i);
MULT MULT201 (clk,in_25_17_r,in_25_17_i,in_25_18_r,in_25_18_i,in_26_17_r,in_26_17_i,in_26_18_r,in_26_18_i,temp_m1_25_17_r,temp_m1_25_17_i,temp_m1_25_18_r,temp_m1_25_18_i,temp_m1_26_17_r,temp_m1_26_17_i,temp_m1_26_18_r,temp_m1_26_18_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly201 (clk,temp_m1_25_17_r,temp_m1_25_17_i,temp_m1_25_18_r,temp_m1_25_18_i,temp_m1_26_17_r,temp_m1_26_17_i,temp_m1_26_18_r,temp_m1_26_18_i,temp_b1_25_17_r,temp_b1_25_17_i,temp_b1_25_18_r,temp_b1_25_18_i,temp_b1_26_17_r,temp_b1_26_17_i,temp_b1_26_18_r,temp_b1_26_18_i);
MULT MULT202 (clk,in_25_19_r,in_25_19_i,in_25_20_r,in_25_20_i,in_26_19_r,in_26_19_i,in_26_20_r,in_26_20_i,temp_m1_25_19_r,temp_m1_25_19_i,temp_m1_25_20_r,temp_m1_25_20_i,temp_m1_26_19_r,temp_m1_26_19_i,temp_m1_26_20_r,temp_m1_26_20_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly202 (clk,temp_m1_25_19_r,temp_m1_25_19_i,temp_m1_25_20_r,temp_m1_25_20_i,temp_m1_26_19_r,temp_m1_26_19_i,temp_m1_26_20_r,temp_m1_26_20_i,temp_b1_25_19_r,temp_b1_25_19_i,temp_b1_25_20_r,temp_b1_25_20_i,temp_b1_26_19_r,temp_b1_26_19_i,temp_b1_26_20_r,temp_b1_26_20_i);
MULT MULT203 (clk,in_25_21_r,in_25_21_i,in_25_22_r,in_25_22_i,in_26_21_r,in_26_21_i,in_26_22_r,in_26_22_i,temp_m1_25_21_r,temp_m1_25_21_i,temp_m1_25_22_r,temp_m1_25_22_i,temp_m1_26_21_r,temp_m1_26_21_i,temp_m1_26_22_r,temp_m1_26_22_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly203 (clk,temp_m1_25_21_r,temp_m1_25_21_i,temp_m1_25_22_r,temp_m1_25_22_i,temp_m1_26_21_r,temp_m1_26_21_i,temp_m1_26_22_r,temp_m1_26_22_i,temp_b1_25_21_r,temp_b1_25_21_i,temp_b1_25_22_r,temp_b1_25_22_i,temp_b1_26_21_r,temp_b1_26_21_i,temp_b1_26_22_r,temp_b1_26_22_i);
MULT MULT204 (clk,in_25_23_r,in_25_23_i,in_25_24_r,in_25_24_i,in_26_23_r,in_26_23_i,in_26_24_r,in_26_24_i,temp_m1_25_23_r,temp_m1_25_23_i,temp_m1_25_24_r,temp_m1_25_24_i,temp_m1_26_23_r,temp_m1_26_23_i,temp_m1_26_24_r,temp_m1_26_24_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly204 (clk,temp_m1_25_23_r,temp_m1_25_23_i,temp_m1_25_24_r,temp_m1_25_24_i,temp_m1_26_23_r,temp_m1_26_23_i,temp_m1_26_24_r,temp_m1_26_24_i,temp_b1_25_23_r,temp_b1_25_23_i,temp_b1_25_24_r,temp_b1_25_24_i,temp_b1_26_23_r,temp_b1_26_23_i,temp_b1_26_24_r,temp_b1_26_24_i);
MULT MULT205 (clk,in_25_25_r,in_25_25_i,in_25_26_r,in_25_26_i,in_26_25_r,in_26_25_i,in_26_26_r,in_26_26_i,temp_m1_25_25_r,temp_m1_25_25_i,temp_m1_25_26_r,temp_m1_25_26_i,temp_m1_26_25_r,temp_m1_26_25_i,temp_m1_26_26_r,temp_m1_26_26_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly205 (clk,temp_m1_25_25_r,temp_m1_25_25_i,temp_m1_25_26_r,temp_m1_25_26_i,temp_m1_26_25_r,temp_m1_26_25_i,temp_m1_26_26_r,temp_m1_26_26_i,temp_b1_25_25_r,temp_b1_25_25_i,temp_b1_25_26_r,temp_b1_25_26_i,temp_b1_26_25_r,temp_b1_26_25_i,temp_b1_26_26_r,temp_b1_26_26_i);
MULT MULT206 (clk,in_25_27_r,in_25_27_i,in_25_28_r,in_25_28_i,in_26_27_r,in_26_27_i,in_26_28_r,in_26_28_i,temp_m1_25_27_r,temp_m1_25_27_i,temp_m1_25_28_r,temp_m1_25_28_i,temp_m1_26_27_r,temp_m1_26_27_i,temp_m1_26_28_r,temp_m1_26_28_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly206 (clk,temp_m1_25_27_r,temp_m1_25_27_i,temp_m1_25_28_r,temp_m1_25_28_i,temp_m1_26_27_r,temp_m1_26_27_i,temp_m1_26_28_r,temp_m1_26_28_i,temp_b1_25_27_r,temp_b1_25_27_i,temp_b1_25_28_r,temp_b1_25_28_i,temp_b1_26_27_r,temp_b1_26_27_i,temp_b1_26_28_r,temp_b1_26_28_i);
MULT MULT207 (clk,in_25_29_r,in_25_29_i,in_25_30_r,in_25_30_i,in_26_29_r,in_26_29_i,in_26_30_r,in_26_30_i,temp_m1_25_29_r,temp_m1_25_29_i,temp_m1_25_30_r,temp_m1_25_30_i,temp_m1_26_29_r,temp_m1_26_29_i,temp_m1_26_30_r,temp_m1_26_30_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly207 (clk,temp_m1_25_29_r,temp_m1_25_29_i,temp_m1_25_30_r,temp_m1_25_30_i,temp_m1_26_29_r,temp_m1_26_29_i,temp_m1_26_30_r,temp_m1_26_30_i,temp_b1_25_29_r,temp_b1_25_29_i,temp_b1_25_30_r,temp_b1_25_30_i,temp_b1_26_29_r,temp_b1_26_29_i,temp_b1_26_30_r,temp_b1_26_30_i);
MULT MULT208 (clk,in_25_31_r,in_25_31_i,in_25_32_r,in_25_32_i,in_26_31_r,in_26_31_i,in_26_32_r,in_26_32_i,temp_m1_25_31_r,temp_m1_25_31_i,temp_m1_25_32_r,temp_m1_25_32_i,temp_m1_26_31_r,temp_m1_26_31_i,temp_m1_26_32_r,temp_m1_26_32_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly208 (clk,temp_m1_25_31_r,temp_m1_25_31_i,temp_m1_25_32_r,temp_m1_25_32_i,temp_m1_26_31_r,temp_m1_26_31_i,temp_m1_26_32_r,temp_m1_26_32_i,temp_b1_25_31_r,temp_b1_25_31_i,temp_b1_25_32_r,temp_b1_25_32_i,temp_b1_26_31_r,temp_b1_26_31_i,temp_b1_26_32_r,temp_b1_26_32_i);
MULT MULT209 (clk,in_27_1_r,in_27_1_i,in_27_2_r,in_27_2_i,in_28_1_r,in_28_1_i,in_28_2_r,in_28_2_i,temp_m1_27_1_r,temp_m1_27_1_i,temp_m1_27_2_r,temp_m1_27_2_i,temp_m1_28_1_r,temp_m1_28_1_i,temp_m1_28_2_r,temp_m1_28_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly209 (clk,temp_m1_27_1_r,temp_m1_27_1_i,temp_m1_27_2_r,temp_m1_27_2_i,temp_m1_28_1_r,temp_m1_28_1_i,temp_m1_28_2_r,temp_m1_28_2_i,temp_b1_27_1_r,temp_b1_27_1_i,temp_b1_27_2_r,temp_b1_27_2_i,temp_b1_28_1_r,temp_b1_28_1_i,temp_b1_28_2_r,temp_b1_28_2_i);
MULT MULT210 (clk,in_27_3_r,in_27_3_i,in_27_4_r,in_27_4_i,in_28_3_r,in_28_3_i,in_28_4_r,in_28_4_i,temp_m1_27_3_r,temp_m1_27_3_i,temp_m1_27_4_r,temp_m1_27_4_i,temp_m1_28_3_r,temp_m1_28_3_i,temp_m1_28_4_r,temp_m1_28_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly210 (clk,temp_m1_27_3_r,temp_m1_27_3_i,temp_m1_27_4_r,temp_m1_27_4_i,temp_m1_28_3_r,temp_m1_28_3_i,temp_m1_28_4_r,temp_m1_28_4_i,temp_b1_27_3_r,temp_b1_27_3_i,temp_b1_27_4_r,temp_b1_27_4_i,temp_b1_28_3_r,temp_b1_28_3_i,temp_b1_28_4_r,temp_b1_28_4_i);
MULT MULT211 (clk,in_27_5_r,in_27_5_i,in_27_6_r,in_27_6_i,in_28_5_r,in_28_5_i,in_28_6_r,in_28_6_i,temp_m1_27_5_r,temp_m1_27_5_i,temp_m1_27_6_r,temp_m1_27_6_i,temp_m1_28_5_r,temp_m1_28_5_i,temp_m1_28_6_r,temp_m1_28_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly211 (clk,temp_m1_27_5_r,temp_m1_27_5_i,temp_m1_27_6_r,temp_m1_27_6_i,temp_m1_28_5_r,temp_m1_28_5_i,temp_m1_28_6_r,temp_m1_28_6_i,temp_b1_27_5_r,temp_b1_27_5_i,temp_b1_27_6_r,temp_b1_27_6_i,temp_b1_28_5_r,temp_b1_28_5_i,temp_b1_28_6_r,temp_b1_28_6_i);
MULT MULT212 (clk,in_27_7_r,in_27_7_i,in_27_8_r,in_27_8_i,in_28_7_r,in_28_7_i,in_28_8_r,in_28_8_i,temp_m1_27_7_r,temp_m1_27_7_i,temp_m1_27_8_r,temp_m1_27_8_i,temp_m1_28_7_r,temp_m1_28_7_i,temp_m1_28_8_r,temp_m1_28_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly212 (clk,temp_m1_27_7_r,temp_m1_27_7_i,temp_m1_27_8_r,temp_m1_27_8_i,temp_m1_28_7_r,temp_m1_28_7_i,temp_m1_28_8_r,temp_m1_28_8_i,temp_b1_27_7_r,temp_b1_27_7_i,temp_b1_27_8_r,temp_b1_27_8_i,temp_b1_28_7_r,temp_b1_28_7_i,temp_b1_28_8_r,temp_b1_28_8_i);
MULT MULT213 (clk,in_27_9_r,in_27_9_i,in_27_10_r,in_27_10_i,in_28_9_r,in_28_9_i,in_28_10_r,in_28_10_i,temp_m1_27_9_r,temp_m1_27_9_i,temp_m1_27_10_r,temp_m1_27_10_i,temp_m1_28_9_r,temp_m1_28_9_i,temp_m1_28_10_r,temp_m1_28_10_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly213 (clk,temp_m1_27_9_r,temp_m1_27_9_i,temp_m1_27_10_r,temp_m1_27_10_i,temp_m1_28_9_r,temp_m1_28_9_i,temp_m1_28_10_r,temp_m1_28_10_i,temp_b1_27_9_r,temp_b1_27_9_i,temp_b1_27_10_r,temp_b1_27_10_i,temp_b1_28_9_r,temp_b1_28_9_i,temp_b1_28_10_r,temp_b1_28_10_i);
MULT MULT214 (clk,in_27_11_r,in_27_11_i,in_27_12_r,in_27_12_i,in_28_11_r,in_28_11_i,in_28_12_r,in_28_12_i,temp_m1_27_11_r,temp_m1_27_11_i,temp_m1_27_12_r,temp_m1_27_12_i,temp_m1_28_11_r,temp_m1_28_11_i,temp_m1_28_12_r,temp_m1_28_12_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly214 (clk,temp_m1_27_11_r,temp_m1_27_11_i,temp_m1_27_12_r,temp_m1_27_12_i,temp_m1_28_11_r,temp_m1_28_11_i,temp_m1_28_12_r,temp_m1_28_12_i,temp_b1_27_11_r,temp_b1_27_11_i,temp_b1_27_12_r,temp_b1_27_12_i,temp_b1_28_11_r,temp_b1_28_11_i,temp_b1_28_12_r,temp_b1_28_12_i);
MULT MULT215 (clk,in_27_13_r,in_27_13_i,in_27_14_r,in_27_14_i,in_28_13_r,in_28_13_i,in_28_14_r,in_28_14_i,temp_m1_27_13_r,temp_m1_27_13_i,temp_m1_27_14_r,temp_m1_27_14_i,temp_m1_28_13_r,temp_m1_28_13_i,temp_m1_28_14_r,temp_m1_28_14_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly215 (clk,temp_m1_27_13_r,temp_m1_27_13_i,temp_m1_27_14_r,temp_m1_27_14_i,temp_m1_28_13_r,temp_m1_28_13_i,temp_m1_28_14_r,temp_m1_28_14_i,temp_b1_27_13_r,temp_b1_27_13_i,temp_b1_27_14_r,temp_b1_27_14_i,temp_b1_28_13_r,temp_b1_28_13_i,temp_b1_28_14_r,temp_b1_28_14_i);
MULT MULT216 (clk,in_27_15_r,in_27_15_i,in_27_16_r,in_27_16_i,in_28_15_r,in_28_15_i,in_28_16_r,in_28_16_i,temp_m1_27_15_r,temp_m1_27_15_i,temp_m1_27_16_r,temp_m1_27_16_i,temp_m1_28_15_r,temp_m1_28_15_i,temp_m1_28_16_r,temp_m1_28_16_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly216 (clk,temp_m1_27_15_r,temp_m1_27_15_i,temp_m1_27_16_r,temp_m1_27_16_i,temp_m1_28_15_r,temp_m1_28_15_i,temp_m1_28_16_r,temp_m1_28_16_i,temp_b1_27_15_r,temp_b1_27_15_i,temp_b1_27_16_r,temp_b1_27_16_i,temp_b1_28_15_r,temp_b1_28_15_i,temp_b1_28_16_r,temp_b1_28_16_i);
MULT MULT217 (clk,in_27_17_r,in_27_17_i,in_27_18_r,in_27_18_i,in_28_17_r,in_28_17_i,in_28_18_r,in_28_18_i,temp_m1_27_17_r,temp_m1_27_17_i,temp_m1_27_18_r,temp_m1_27_18_i,temp_m1_28_17_r,temp_m1_28_17_i,temp_m1_28_18_r,temp_m1_28_18_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly217 (clk,temp_m1_27_17_r,temp_m1_27_17_i,temp_m1_27_18_r,temp_m1_27_18_i,temp_m1_28_17_r,temp_m1_28_17_i,temp_m1_28_18_r,temp_m1_28_18_i,temp_b1_27_17_r,temp_b1_27_17_i,temp_b1_27_18_r,temp_b1_27_18_i,temp_b1_28_17_r,temp_b1_28_17_i,temp_b1_28_18_r,temp_b1_28_18_i);
MULT MULT218 (clk,in_27_19_r,in_27_19_i,in_27_20_r,in_27_20_i,in_28_19_r,in_28_19_i,in_28_20_r,in_28_20_i,temp_m1_27_19_r,temp_m1_27_19_i,temp_m1_27_20_r,temp_m1_27_20_i,temp_m1_28_19_r,temp_m1_28_19_i,temp_m1_28_20_r,temp_m1_28_20_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly218 (clk,temp_m1_27_19_r,temp_m1_27_19_i,temp_m1_27_20_r,temp_m1_27_20_i,temp_m1_28_19_r,temp_m1_28_19_i,temp_m1_28_20_r,temp_m1_28_20_i,temp_b1_27_19_r,temp_b1_27_19_i,temp_b1_27_20_r,temp_b1_27_20_i,temp_b1_28_19_r,temp_b1_28_19_i,temp_b1_28_20_r,temp_b1_28_20_i);
MULT MULT219 (clk,in_27_21_r,in_27_21_i,in_27_22_r,in_27_22_i,in_28_21_r,in_28_21_i,in_28_22_r,in_28_22_i,temp_m1_27_21_r,temp_m1_27_21_i,temp_m1_27_22_r,temp_m1_27_22_i,temp_m1_28_21_r,temp_m1_28_21_i,temp_m1_28_22_r,temp_m1_28_22_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly219 (clk,temp_m1_27_21_r,temp_m1_27_21_i,temp_m1_27_22_r,temp_m1_27_22_i,temp_m1_28_21_r,temp_m1_28_21_i,temp_m1_28_22_r,temp_m1_28_22_i,temp_b1_27_21_r,temp_b1_27_21_i,temp_b1_27_22_r,temp_b1_27_22_i,temp_b1_28_21_r,temp_b1_28_21_i,temp_b1_28_22_r,temp_b1_28_22_i);
MULT MULT220 (clk,in_27_23_r,in_27_23_i,in_27_24_r,in_27_24_i,in_28_23_r,in_28_23_i,in_28_24_r,in_28_24_i,temp_m1_27_23_r,temp_m1_27_23_i,temp_m1_27_24_r,temp_m1_27_24_i,temp_m1_28_23_r,temp_m1_28_23_i,temp_m1_28_24_r,temp_m1_28_24_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly220 (clk,temp_m1_27_23_r,temp_m1_27_23_i,temp_m1_27_24_r,temp_m1_27_24_i,temp_m1_28_23_r,temp_m1_28_23_i,temp_m1_28_24_r,temp_m1_28_24_i,temp_b1_27_23_r,temp_b1_27_23_i,temp_b1_27_24_r,temp_b1_27_24_i,temp_b1_28_23_r,temp_b1_28_23_i,temp_b1_28_24_r,temp_b1_28_24_i);
MULT MULT221 (clk,in_27_25_r,in_27_25_i,in_27_26_r,in_27_26_i,in_28_25_r,in_28_25_i,in_28_26_r,in_28_26_i,temp_m1_27_25_r,temp_m1_27_25_i,temp_m1_27_26_r,temp_m1_27_26_i,temp_m1_28_25_r,temp_m1_28_25_i,temp_m1_28_26_r,temp_m1_28_26_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly221 (clk,temp_m1_27_25_r,temp_m1_27_25_i,temp_m1_27_26_r,temp_m1_27_26_i,temp_m1_28_25_r,temp_m1_28_25_i,temp_m1_28_26_r,temp_m1_28_26_i,temp_b1_27_25_r,temp_b1_27_25_i,temp_b1_27_26_r,temp_b1_27_26_i,temp_b1_28_25_r,temp_b1_28_25_i,temp_b1_28_26_r,temp_b1_28_26_i);
MULT MULT222 (clk,in_27_27_r,in_27_27_i,in_27_28_r,in_27_28_i,in_28_27_r,in_28_27_i,in_28_28_r,in_28_28_i,temp_m1_27_27_r,temp_m1_27_27_i,temp_m1_27_28_r,temp_m1_27_28_i,temp_m1_28_27_r,temp_m1_28_27_i,temp_m1_28_28_r,temp_m1_28_28_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly222 (clk,temp_m1_27_27_r,temp_m1_27_27_i,temp_m1_27_28_r,temp_m1_27_28_i,temp_m1_28_27_r,temp_m1_28_27_i,temp_m1_28_28_r,temp_m1_28_28_i,temp_b1_27_27_r,temp_b1_27_27_i,temp_b1_27_28_r,temp_b1_27_28_i,temp_b1_28_27_r,temp_b1_28_27_i,temp_b1_28_28_r,temp_b1_28_28_i);
MULT MULT223 (clk,in_27_29_r,in_27_29_i,in_27_30_r,in_27_30_i,in_28_29_r,in_28_29_i,in_28_30_r,in_28_30_i,temp_m1_27_29_r,temp_m1_27_29_i,temp_m1_27_30_r,temp_m1_27_30_i,temp_m1_28_29_r,temp_m1_28_29_i,temp_m1_28_30_r,temp_m1_28_30_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly223 (clk,temp_m1_27_29_r,temp_m1_27_29_i,temp_m1_27_30_r,temp_m1_27_30_i,temp_m1_28_29_r,temp_m1_28_29_i,temp_m1_28_30_r,temp_m1_28_30_i,temp_b1_27_29_r,temp_b1_27_29_i,temp_b1_27_30_r,temp_b1_27_30_i,temp_b1_28_29_r,temp_b1_28_29_i,temp_b1_28_30_r,temp_b1_28_30_i);
MULT MULT224 (clk,in_27_31_r,in_27_31_i,in_27_32_r,in_27_32_i,in_28_31_r,in_28_31_i,in_28_32_r,in_28_32_i,temp_m1_27_31_r,temp_m1_27_31_i,temp_m1_27_32_r,temp_m1_27_32_i,temp_m1_28_31_r,temp_m1_28_31_i,temp_m1_28_32_r,temp_m1_28_32_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly224 (clk,temp_m1_27_31_r,temp_m1_27_31_i,temp_m1_27_32_r,temp_m1_27_32_i,temp_m1_28_31_r,temp_m1_28_31_i,temp_m1_28_32_r,temp_m1_28_32_i,temp_b1_27_31_r,temp_b1_27_31_i,temp_b1_27_32_r,temp_b1_27_32_i,temp_b1_28_31_r,temp_b1_28_31_i,temp_b1_28_32_r,temp_b1_28_32_i);
MULT MULT225 (clk,in_29_1_r,in_29_1_i,in_29_2_r,in_29_2_i,in_30_1_r,in_30_1_i,in_30_2_r,in_30_2_i,temp_m1_29_1_r,temp_m1_29_1_i,temp_m1_29_2_r,temp_m1_29_2_i,temp_m1_30_1_r,temp_m1_30_1_i,temp_m1_30_2_r,temp_m1_30_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly225 (clk,temp_m1_29_1_r,temp_m1_29_1_i,temp_m1_29_2_r,temp_m1_29_2_i,temp_m1_30_1_r,temp_m1_30_1_i,temp_m1_30_2_r,temp_m1_30_2_i,temp_b1_29_1_r,temp_b1_29_1_i,temp_b1_29_2_r,temp_b1_29_2_i,temp_b1_30_1_r,temp_b1_30_1_i,temp_b1_30_2_r,temp_b1_30_2_i);
MULT MULT226 (clk,in_29_3_r,in_29_3_i,in_29_4_r,in_29_4_i,in_30_3_r,in_30_3_i,in_30_4_r,in_30_4_i,temp_m1_29_3_r,temp_m1_29_3_i,temp_m1_29_4_r,temp_m1_29_4_i,temp_m1_30_3_r,temp_m1_30_3_i,temp_m1_30_4_r,temp_m1_30_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly226 (clk,temp_m1_29_3_r,temp_m1_29_3_i,temp_m1_29_4_r,temp_m1_29_4_i,temp_m1_30_3_r,temp_m1_30_3_i,temp_m1_30_4_r,temp_m1_30_4_i,temp_b1_29_3_r,temp_b1_29_3_i,temp_b1_29_4_r,temp_b1_29_4_i,temp_b1_30_3_r,temp_b1_30_3_i,temp_b1_30_4_r,temp_b1_30_4_i);
MULT MULT227 (clk,in_29_5_r,in_29_5_i,in_29_6_r,in_29_6_i,in_30_5_r,in_30_5_i,in_30_6_r,in_30_6_i,temp_m1_29_5_r,temp_m1_29_5_i,temp_m1_29_6_r,temp_m1_29_6_i,temp_m1_30_5_r,temp_m1_30_5_i,temp_m1_30_6_r,temp_m1_30_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly227 (clk,temp_m1_29_5_r,temp_m1_29_5_i,temp_m1_29_6_r,temp_m1_29_6_i,temp_m1_30_5_r,temp_m1_30_5_i,temp_m1_30_6_r,temp_m1_30_6_i,temp_b1_29_5_r,temp_b1_29_5_i,temp_b1_29_6_r,temp_b1_29_6_i,temp_b1_30_5_r,temp_b1_30_5_i,temp_b1_30_6_r,temp_b1_30_6_i);
MULT MULT228 (clk,in_29_7_r,in_29_7_i,in_29_8_r,in_29_8_i,in_30_7_r,in_30_7_i,in_30_8_r,in_30_8_i,temp_m1_29_7_r,temp_m1_29_7_i,temp_m1_29_8_r,temp_m1_29_8_i,temp_m1_30_7_r,temp_m1_30_7_i,temp_m1_30_8_r,temp_m1_30_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly228 (clk,temp_m1_29_7_r,temp_m1_29_7_i,temp_m1_29_8_r,temp_m1_29_8_i,temp_m1_30_7_r,temp_m1_30_7_i,temp_m1_30_8_r,temp_m1_30_8_i,temp_b1_29_7_r,temp_b1_29_7_i,temp_b1_29_8_r,temp_b1_29_8_i,temp_b1_30_7_r,temp_b1_30_7_i,temp_b1_30_8_r,temp_b1_30_8_i);
MULT MULT229 (clk,in_29_9_r,in_29_9_i,in_29_10_r,in_29_10_i,in_30_9_r,in_30_9_i,in_30_10_r,in_30_10_i,temp_m1_29_9_r,temp_m1_29_9_i,temp_m1_29_10_r,temp_m1_29_10_i,temp_m1_30_9_r,temp_m1_30_9_i,temp_m1_30_10_r,temp_m1_30_10_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly229 (clk,temp_m1_29_9_r,temp_m1_29_9_i,temp_m1_29_10_r,temp_m1_29_10_i,temp_m1_30_9_r,temp_m1_30_9_i,temp_m1_30_10_r,temp_m1_30_10_i,temp_b1_29_9_r,temp_b1_29_9_i,temp_b1_29_10_r,temp_b1_29_10_i,temp_b1_30_9_r,temp_b1_30_9_i,temp_b1_30_10_r,temp_b1_30_10_i);
MULT MULT230 (clk,in_29_11_r,in_29_11_i,in_29_12_r,in_29_12_i,in_30_11_r,in_30_11_i,in_30_12_r,in_30_12_i,temp_m1_29_11_r,temp_m1_29_11_i,temp_m1_29_12_r,temp_m1_29_12_i,temp_m1_30_11_r,temp_m1_30_11_i,temp_m1_30_12_r,temp_m1_30_12_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly230 (clk,temp_m1_29_11_r,temp_m1_29_11_i,temp_m1_29_12_r,temp_m1_29_12_i,temp_m1_30_11_r,temp_m1_30_11_i,temp_m1_30_12_r,temp_m1_30_12_i,temp_b1_29_11_r,temp_b1_29_11_i,temp_b1_29_12_r,temp_b1_29_12_i,temp_b1_30_11_r,temp_b1_30_11_i,temp_b1_30_12_r,temp_b1_30_12_i);
MULT MULT231 (clk,in_29_13_r,in_29_13_i,in_29_14_r,in_29_14_i,in_30_13_r,in_30_13_i,in_30_14_r,in_30_14_i,temp_m1_29_13_r,temp_m1_29_13_i,temp_m1_29_14_r,temp_m1_29_14_i,temp_m1_30_13_r,temp_m1_30_13_i,temp_m1_30_14_r,temp_m1_30_14_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly231 (clk,temp_m1_29_13_r,temp_m1_29_13_i,temp_m1_29_14_r,temp_m1_29_14_i,temp_m1_30_13_r,temp_m1_30_13_i,temp_m1_30_14_r,temp_m1_30_14_i,temp_b1_29_13_r,temp_b1_29_13_i,temp_b1_29_14_r,temp_b1_29_14_i,temp_b1_30_13_r,temp_b1_30_13_i,temp_b1_30_14_r,temp_b1_30_14_i);
MULT MULT232 (clk,in_29_15_r,in_29_15_i,in_29_16_r,in_29_16_i,in_30_15_r,in_30_15_i,in_30_16_r,in_30_16_i,temp_m1_29_15_r,temp_m1_29_15_i,temp_m1_29_16_r,temp_m1_29_16_i,temp_m1_30_15_r,temp_m1_30_15_i,temp_m1_30_16_r,temp_m1_30_16_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly232 (clk,temp_m1_29_15_r,temp_m1_29_15_i,temp_m1_29_16_r,temp_m1_29_16_i,temp_m1_30_15_r,temp_m1_30_15_i,temp_m1_30_16_r,temp_m1_30_16_i,temp_b1_29_15_r,temp_b1_29_15_i,temp_b1_29_16_r,temp_b1_29_16_i,temp_b1_30_15_r,temp_b1_30_15_i,temp_b1_30_16_r,temp_b1_30_16_i);
MULT MULT233 (clk,in_29_17_r,in_29_17_i,in_29_18_r,in_29_18_i,in_30_17_r,in_30_17_i,in_30_18_r,in_30_18_i,temp_m1_29_17_r,temp_m1_29_17_i,temp_m1_29_18_r,temp_m1_29_18_i,temp_m1_30_17_r,temp_m1_30_17_i,temp_m1_30_18_r,temp_m1_30_18_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly233 (clk,temp_m1_29_17_r,temp_m1_29_17_i,temp_m1_29_18_r,temp_m1_29_18_i,temp_m1_30_17_r,temp_m1_30_17_i,temp_m1_30_18_r,temp_m1_30_18_i,temp_b1_29_17_r,temp_b1_29_17_i,temp_b1_29_18_r,temp_b1_29_18_i,temp_b1_30_17_r,temp_b1_30_17_i,temp_b1_30_18_r,temp_b1_30_18_i);
MULT MULT234 (clk,in_29_19_r,in_29_19_i,in_29_20_r,in_29_20_i,in_30_19_r,in_30_19_i,in_30_20_r,in_30_20_i,temp_m1_29_19_r,temp_m1_29_19_i,temp_m1_29_20_r,temp_m1_29_20_i,temp_m1_30_19_r,temp_m1_30_19_i,temp_m1_30_20_r,temp_m1_30_20_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly234 (clk,temp_m1_29_19_r,temp_m1_29_19_i,temp_m1_29_20_r,temp_m1_29_20_i,temp_m1_30_19_r,temp_m1_30_19_i,temp_m1_30_20_r,temp_m1_30_20_i,temp_b1_29_19_r,temp_b1_29_19_i,temp_b1_29_20_r,temp_b1_29_20_i,temp_b1_30_19_r,temp_b1_30_19_i,temp_b1_30_20_r,temp_b1_30_20_i);
MULT MULT235 (clk,in_29_21_r,in_29_21_i,in_29_22_r,in_29_22_i,in_30_21_r,in_30_21_i,in_30_22_r,in_30_22_i,temp_m1_29_21_r,temp_m1_29_21_i,temp_m1_29_22_r,temp_m1_29_22_i,temp_m1_30_21_r,temp_m1_30_21_i,temp_m1_30_22_r,temp_m1_30_22_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly235 (clk,temp_m1_29_21_r,temp_m1_29_21_i,temp_m1_29_22_r,temp_m1_29_22_i,temp_m1_30_21_r,temp_m1_30_21_i,temp_m1_30_22_r,temp_m1_30_22_i,temp_b1_29_21_r,temp_b1_29_21_i,temp_b1_29_22_r,temp_b1_29_22_i,temp_b1_30_21_r,temp_b1_30_21_i,temp_b1_30_22_r,temp_b1_30_22_i);
MULT MULT236 (clk,in_29_23_r,in_29_23_i,in_29_24_r,in_29_24_i,in_30_23_r,in_30_23_i,in_30_24_r,in_30_24_i,temp_m1_29_23_r,temp_m1_29_23_i,temp_m1_29_24_r,temp_m1_29_24_i,temp_m1_30_23_r,temp_m1_30_23_i,temp_m1_30_24_r,temp_m1_30_24_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly236 (clk,temp_m1_29_23_r,temp_m1_29_23_i,temp_m1_29_24_r,temp_m1_29_24_i,temp_m1_30_23_r,temp_m1_30_23_i,temp_m1_30_24_r,temp_m1_30_24_i,temp_b1_29_23_r,temp_b1_29_23_i,temp_b1_29_24_r,temp_b1_29_24_i,temp_b1_30_23_r,temp_b1_30_23_i,temp_b1_30_24_r,temp_b1_30_24_i);
MULT MULT237 (clk,in_29_25_r,in_29_25_i,in_29_26_r,in_29_26_i,in_30_25_r,in_30_25_i,in_30_26_r,in_30_26_i,temp_m1_29_25_r,temp_m1_29_25_i,temp_m1_29_26_r,temp_m1_29_26_i,temp_m1_30_25_r,temp_m1_30_25_i,temp_m1_30_26_r,temp_m1_30_26_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly237 (clk,temp_m1_29_25_r,temp_m1_29_25_i,temp_m1_29_26_r,temp_m1_29_26_i,temp_m1_30_25_r,temp_m1_30_25_i,temp_m1_30_26_r,temp_m1_30_26_i,temp_b1_29_25_r,temp_b1_29_25_i,temp_b1_29_26_r,temp_b1_29_26_i,temp_b1_30_25_r,temp_b1_30_25_i,temp_b1_30_26_r,temp_b1_30_26_i);
MULT MULT238 (clk,in_29_27_r,in_29_27_i,in_29_28_r,in_29_28_i,in_30_27_r,in_30_27_i,in_30_28_r,in_30_28_i,temp_m1_29_27_r,temp_m1_29_27_i,temp_m1_29_28_r,temp_m1_29_28_i,temp_m1_30_27_r,temp_m1_30_27_i,temp_m1_30_28_r,temp_m1_30_28_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly238 (clk,temp_m1_29_27_r,temp_m1_29_27_i,temp_m1_29_28_r,temp_m1_29_28_i,temp_m1_30_27_r,temp_m1_30_27_i,temp_m1_30_28_r,temp_m1_30_28_i,temp_b1_29_27_r,temp_b1_29_27_i,temp_b1_29_28_r,temp_b1_29_28_i,temp_b1_30_27_r,temp_b1_30_27_i,temp_b1_30_28_r,temp_b1_30_28_i);
MULT MULT239 (clk,in_29_29_r,in_29_29_i,in_29_30_r,in_29_30_i,in_30_29_r,in_30_29_i,in_30_30_r,in_30_30_i,temp_m1_29_29_r,temp_m1_29_29_i,temp_m1_29_30_r,temp_m1_29_30_i,temp_m1_30_29_r,temp_m1_30_29_i,temp_m1_30_30_r,temp_m1_30_30_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly239 (clk,temp_m1_29_29_r,temp_m1_29_29_i,temp_m1_29_30_r,temp_m1_29_30_i,temp_m1_30_29_r,temp_m1_30_29_i,temp_m1_30_30_r,temp_m1_30_30_i,temp_b1_29_29_r,temp_b1_29_29_i,temp_b1_29_30_r,temp_b1_29_30_i,temp_b1_30_29_r,temp_b1_30_29_i,temp_b1_30_30_r,temp_b1_30_30_i);
MULT MULT240 (clk,in_29_31_r,in_29_31_i,in_29_32_r,in_29_32_i,in_30_31_r,in_30_31_i,in_30_32_r,in_30_32_i,temp_m1_29_31_r,temp_m1_29_31_i,temp_m1_29_32_r,temp_m1_29_32_i,temp_m1_30_31_r,temp_m1_30_31_i,temp_m1_30_32_r,temp_m1_30_32_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly240 (clk,temp_m1_29_31_r,temp_m1_29_31_i,temp_m1_29_32_r,temp_m1_29_32_i,temp_m1_30_31_r,temp_m1_30_31_i,temp_m1_30_32_r,temp_m1_30_32_i,temp_b1_29_31_r,temp_b1_29_31_i,temp_b1_29_32_r,temp_b1_29_32_i,temp_b1_30_31_r,temp_b1_30_31_i,temp_b1_30_32_r,temp_b1_30_32_i);
MULT MULT241 (clk,in_31_1_r,in_31_1_i,in_31_2_r,in_31_2_i,in_32_1_r,in_32_1_i,in_32_2_r,in_32_2_i,temp_m1_31_1_r,temp_m1_31_1_i,temp_m1_31_2_r,temp_m1_31_2_i,temp_m1_32_1_r,temp_m1_32_1_i,temp_m1_32_2_r,temp_m1_32_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly241 (clk,temp_m1_31_1_r,temp_m1_31_1_i,temp_m1_31_2_r,temp_m1_31_2_i,temp_m1_32_1_r,temp_m1_32_1_i,temp_m1_32_2_r,temp_m1_32_2_i,temp_b1_31_1_r,temp_b1_31_1_i,temp_b1_31_2_r,temp_b1_31_2_i,temp_b1_32_1_r,temp_b1_32_1_i,temp_b1_32_2_r,temp_b1_32_2_i);
MULT MULT242 (clk,in_31_3_r,in_31_3_i,in_31_4_r,in_31_4_i,in_32_3_r,in_32_3_i,in_32_4_r,in_32_4_i,temp_m1_31_3_r,temp_m1_31_3_i,temp_m1_31_4_r,temp_m1_31_4_i,temp_m1_32_3_r,temp_m1_32_3_i,temp_m1_32_4_r,temp_m1_32_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly242 (clk,temp_m1_31_3_r,temp_m1_31_3_i,temp_m1_31_4_r,temp_m1_31_4_i,temp_m1_32_3_r,temp_m1_32_3_i,temp_m1_32_4_r,temp_m1_32_4_i,temp_b1_31_3_r,temp_b1_31_3_i,temp_b1_31_4_r,temp_b1_31_4_i,temp_b1_32_3_r,temp_b1_32_3_i,temp_b1_32_4_r,temp_b1_32_4_i);
MULT MULT243 (clk,in_31_5_r,in_31_5_i,in_31_6_r,in_31_6_i,in_32_5_r,in_32_5_i,in_32_6_r,in_32_6_i,temp_m1_31_5_r,temp_m1_31_5_i,temp_m1_31_6_r,temp_m1_31_6_i,temp_m1_32_5_r,temp_m1_32_5_i,temp_m1_32_6_r,temp_m1_32_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly243 (clk,temp_m1_31_5_r,temp_m1_31_5_i,temp_m1_31_6_r,temp_m1_31_6_i,temp_m1_32_5_r,temp_m1_32_5_i,temp_m1_32_6_r,temp_m1_32_6_i,temp_b1_31_5_r,temp_b1_31_5_i,temp_b1_31_6_r,temp_b1_31_6_i,temp_b1_32_5_r,temp_b1_32_5_i,temp_b1_32_6_r,temp_b1_32_6_i);
MULT MULT244 (clk,in_31_7_r,in_31_7_i,in_31_8_r,in_31_8_i,in_32_7_r,in_32_7_i,in_32_8_r,in_32_8_i,temp_m1_31_7_r,temp_m1_31_7_i,temp_m1_31_8_r,temp_m1_31_8_i,temp_m1_32_7_r,temp_m1_32_7_i,temp_m1_32_8_r,temp_m1_32_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly244 (clk,temp_m1_31_7_r,temp_m1_31_7_i,temp_m1_31_8_r,temp_m1_31_8_i,temp_m1_32_7_r,temp_m1_32_7_i,temp_m1_32_8_r,temp_m1_32_8_i,temp_b1_31_7_r,temp_b1_31_7_i,temp_b1_31_8_r,temp_b1_31_8_i,temp_b1_32_7_r,temp_b1_32_7_i,temp_b1_32_8_r,temp_b1_32_8_i);
MULT MULT245 (clk,in_31_9_r,in_31_9_i,in_31_10_r,in_31_10_i,in_32_9_r,in_32_9_i,in_32_10_r,in_32_10_i,temp_m1_31_9_r,temp_m1_31_9_i,temp_m1_31_10_r,temp_m1_31_10_i,temp_m1_32_9_r,temp_m1_32_9_i,temp_m1_32_10_r,temp_m1_32_10_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly245 (clk,temp_m1_31_9_r,temp_m1_31_9_i,temp_m1_31_10_r,temp_m1_31_10_i,temp_m1_32_9_r,temp_m1_32_9_i,temp_m1_32_10_r,temp_m1_32_10_i,temp_b1_31_9_r,temp_b1_31_9_i,temp_b1_31_10_r,temp_b1_31_10_i,temp_b1_32_9_r,temp_b1_32_9_i,temp_b1_32_10_r,temp_b1_32_10_i);
MULT MULT246 (clk,in_31_11_r,in_31_11_i,in_31_12_r,in_31_12_i,in_32_11_r,in_32_11_i,in_32_12_r,in_32_12_i,temp_m1_31_11_r,temp_m1_31_11_i,temp_m1_31_12_r,temp_m1_31_12_i,temp_m1_32_11_r,temp_m1_32_11_i,temp_m1_32_12_r,temp_m1_32_12_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly246 (clk,temp_m1_31_11_r,temp_m1_31_11_i,temp_m1_31_12_r,temp_m1_31_12_i,temp_m1_32_11_r,temp_m1_32_11_i,temp_m1_32_12_r,temp_m1_32_12_i,temp_b1_31_11_r,temp_b1_31_11_i,temp_b1_31_12_r,temp_b1_31_12_i,temp_b1_32_11_r,temp_b1_32_11_i,temp_b1_32_12_r,temp_b1_32_12_i);
MULT MULT247 (clk,in_31_13_r,in_31_13_i,in_31_14_r,in_31_14_i,in_32_13_r,in_32_13_i,in_32_14_r,in_32_14_i,temp_m1_31_13_r,temp_m1_31_13_i,temp_m1_31_14_r,temp_m1_31_14_i,temp_m1_32_13_r,temp_m1_32_13_i,temp_m1_32_14_r,temp_m1_32_14_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly247 (clk,temp_m1_31_13_r,temp_m1_31_13_i,temp_m1_31_14_r,temp_m1_31_14_i,temp_m1_32_13_r,temp_m1_32_13_i,temp_m1_32_14_r,temp_m1_32_14_i,temp_b1_31_13_r,temp_b1_31_13_i,temp_b1_31_14_r,temp_b1_31_14_i,temp_b1_32_13_r,temp_b1_32_13_i,temp_b1_32_14_r,temp_b1_32_14_i);
MULT MULT248 (clk,in_31_15_r,in_31_15_i,in_31_16_r,in_31_16_i,in_32_15_r,in_32_15_i,in_32_16_r,in_32_16_i,temp_m1_31_15_r,temp_m1_31_15_i,temp_m1_31_16_r,temp_m1_31_16_i,temp_m1_32_15_r,temp_m1_32_15_i,temp_m1_32_16_r,temp_m1_32_16_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly248 (clk,temp_m1_31_15_r,temp_m1_31_15_i,temp_m1_31_16_r,temp_m1_31_16_i,temp_m1_32_15_r,temp_m1_32_15_i,temp_m1_32_16_r,temp_m1_32_16_i,temp_b1_31_15_r,temp_b1_31_15_i,temp_b1_31_16_r,temp_b1_31_16_i,temp_b1_32_15_r,temp_b1_32_15_i,temp_b1_32_16_r,temp_b1_32_16_i);
MULT MULT249 (clk,in_31_17_r,in_31_17_i,in_31_18_r,in_31_18_i,in_32_17_r,in_32_17_i,in_32_18_r,in_32_18_i,temp_m1_31_17_r,temp_m1_31_17_i,temp_m1_31_18_r,temp_m1_31_18_i,temp_m1_32_17_r,temp_m1_32_17_i,temp_m1_32_18_r,temp_m1_32_18_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly249 (clk,temp_m1_31_17_r,temp_m1_31_17_i,temp_m1_31_18_r,temp_m1_31_18_i,temp_m1_32_17_r,temp_m1_32_17_i,temp_m1_32_18_r,temp_m1_32_18_i,temp_b1_31_17_r,temp_b1_31_17_i,temp_b1_31_18_r,temp_b1_31_18_i,temp_b1_32_17_r,temp_b1_32_17_i,temp_b1_32_18_r,temp_b1_32_18_i);
MULT MULT250 (clk,in_31_19_r,in_31_19_i,in_31_20_r,in_31_20_i,in_32_19_r,in_32_19_i,in_32_20_r,in_32_20_i,temp_m1_31_19_r,temp_m1_31_19_i,temp_m1_31_20_r,temp_m1_31_20_i,temp_m1_32_19_r,temp_m1_32_19_i,temp_m1_32_20_r,temp_m1_32_20_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly250 (clk,temp_m1_31_19_r,temp_m1_31_19_i,temp_m1_31_20_r,temp_m1_31_20_i,temp_m1_32_19_r,temp_m1_32_19_i,temp_m1_32_20_r,temp_m1_32_20_i,temp_b1_31_19_r,temp_b1_31_19_i,temp_b1_31_20_r,temp_b1_31_20_i,temp_b1_32_19_r,temp_b1_32_19_i,temp_b1_32_20_r,temp_b1_32_20_i);
MULT MULT251 (clk,in_31_21_r,in_31_21_i,in_31_22_r,in_31_22_i,in_32_21_r,in_32_21_i,in_32_22_r,in_32_22_i,temp_m1_31_21_r,temp_m1_31_21_i,temp_m1_31_22_r,temp_m1_31_22_i,temp_m1_32_21_r,temp_m1_32_21_i,temp_m1_32_22_r,temp_m1_32_22_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly251 (clk,temp_m1_31_21_r,temp_m1_31_21_i,temp_m1_31_22_r,temp_m1_31_22_i,temp_m1_32_21_r,temp_m1_32_21_i,temp_m1_32_22_r,temp_m1_32_22_i,temp_b1_31_21_r,temp_b1_31_21_i,temp_b1_31_22_r,temp_b1_31_22_i,temp_b1_32_21_r,temp_b1_32_21_i,temp_b1_32_22_r,temp_b1_32_22_i);
MULT MULT252 (clk,in_31_23_r,in_31_23_i,in_31_24_r,in_31_24_i,in_32_23_r,in_32_23_i,in_32_24_r,in_32_24_i,temp_m1_31_23_r,temp_m1_31_23_i,temp_m1_31_24_r,temp_m1_31_24_i,temp_m1_32_23_r,temp_m1_32_23_i,temp_m1_32_24_r,temp_m1_32_24_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly252 (clk,temp_m1_31_23_r,temp_m1_31_23_i,temp_m1_31_24_r,temp_m1_31_24_i,temp_m1_32_23_r,temp_m1_32_23_i,temp_m1_32_24_r,temp_m1_32_24_i,temp_b1_31_23_r,temp_b1_31_23_i,temp_b1_31_24_r,temp_b1_31_24_i,temp_b1_32_23_r,temp_b1_32_23_i,temp_b1_32_24_r,temp_b1_32_24_i);
MULT MULT253 (clk,in_31_25_r,in_31_25_i,in_31_26_r,in_31_26_i,in_32_25_r,in_32_25_i,in_32_26_r,in_32_26_i,temp_m1_31_25_r,temp_m1_31_25_i,temp_m1_31_26_r,temp_m1_31_26_i,temp_m1_32_25_r,temp_m1_32_25_i,temp_m1_32_26_r,temp_m1_32_26_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly253 (clk,temp_m1_31_25_r,temp_m1_31_25_i,temp_m1_31_26_r,temp_m1_31_26_i,temp_m1_32_25_r,temp_m1_32_25_i,temp_m1_32_26_r,temp_m1_32_26_i,temp_b1_31_25_r,temp_b1_31_25_i,temp_b1_31_26_r,temp_b1_31_26_i,temp_b1_32_25_r,temp_b1_32_25_i,temp_b1_32_26_r,temp_b1_32_26_i);
MULT MULT254 (clk,in_31_27_r,in_31_27_i,in_31_28_r,in_31_28_i,in_32_27_r,in_32_27_i,in_32_28_r,in_32_28_i,temp_m1_31_27_r,temp_m1_31_27_i,temp_m1_31_28_r,temp_m1_31_28_i,temp_m1_32_27_r,temp_m1_32_27_i,temp_m1_32_28_r,temp_m1_32_28_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly254 (clk,temp_m1_31_27_r,temp_m1_31_27_i,temp_m1_31_28_r,temp_m1_31_28_i,temp_m1_32_27_r,temp_m1_32_27_i,temp_m1_32_28_r,temp_m1_32_28_i,temp_b1_31_27_r,temp_b1_31_27_i,temp_b1_31_28_r,temp_b1_31_28_i,temp_b1_32_27_r,temp_b1_32_27_i,temp_b1_32_28_r,temp_b1_32_28_i);
MULT MULT255 (clk,in_31_29_r,in_31_29_i,in_31_30_r,in_31_30_i,in_32_29_r,in_32_29_i,in_32_30_r,in_32_30_i,temp_m1_31_29_r,temp_m1_31_29_i,temp_m1_31_30_r,temp_m1_31_30_i,temp_m1_32_29_r,temp_m1_32_29_i,temp_m1_32_30_r,temp_m1_32_30_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly255 (clk,temp_m1_31_29_r,temp_m1_31_29_i,temp_m1_31_30_r,temp_m1_31_30_i,temp_m1_32_29_r,temp_m1_32_29_i,temp_m1_32_30_r,temp_m1_32_30_i,temp_b1_31_29_r,temp_b1_31_29_i,temp_b1_31_30_r,temp_b1_31_30_i,temp_b1_32_29_r,temp_b1_32_29_i,temp_b1_32_30_r,temp_b1_32_30_i);
MULT MULT256 (clk,in_31_31_r,in_31_31_i,in_31_32_r,in_31_32_i,in_32_31_r,in_32_31_i,in_32_32_r,in_32_32_i,temp_m1_31_31_r,temp_m1_31_31_i,temp_m1_31_32_r,temp_m1_31_32_i,temp_m1_32_31_r,temp_m1_32_31_i,temp_m1_32_32_r,temp_m1_32_32_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly256 (clk,temp_m1_31_31_r,temp_m1_31_31_i,temp_m1_31_32_r,temp_m1_31_32_i,temp_m1_32_31_r,temp_m1_32_31_i,temp_m1_32_32_r,temp_m1_32_32_i,temp_b1_31_31_r,temp_b1_31_31_i,temp_b1_31_32_r,temp_b1_31_32_i,temp_b1_32_31_r,temp_b1_32_31_i,temp_b1_32_32_r,temp_b1_32_32_i);
MULT MULT257 (clk,temp_b1_1_1_r,temp_b1_1_1_i,temp_b1_1_3_r,temp_b1_1_3_i,temp_b1_3_1_r,temp_b1_3_1_i,temp_b1_3_3_r,temp_b1_3_3_i,temp_m2_1_1_r,temp_m2_1_1_i,temp_m2_1_3_r,temp_m2_1_3_i,temp_m2_3_1_r,temp_m2_3_1_i,temp_m2_3_3_r,temp_m2_3_3_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly257 (clk,temp_m2_1_1_r,temp_m2_1_1_i,temp_m2_1_3_r,temp_m2_1_3_i,temp_m2_3_1_r,temp_m2_3_1_i,temp_m2_3_3_r,temp_m2_3_3_i,temp_b2_1_1_r,temp_b2_1_1_i,temp_b2_1_3_r,temp_b2_1_3_i,temp_b2_3_1_r,temp_b2_3_1_i,temp_b2_3_3_r,temp_b2_3_3_i);
MULT MULT258 (clk,temp_b1_1_2_r,temp_b1_1_2_i,temp_b1_1_4_r,temp_b1_1_4_i,temp_b1_3_2_r,temp_b1_3_2_i,temp_b1_3_4_r,temp_b1_3_4_i,temp_m2_1_2_r,temp_m2_1_2_i,temp_m2_1_4_r,temp_m2_1_4_i,temp_m2_3_2_r,temp_m2_3_2_i,temp_m2_3_4_r,temp_m2_3_4_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly258 (clk,temp_m2_1_2_r,temp_m2_1_2_i,temp_m2_1_4_r,temp_m2_1_4_i,temp_m2_3_2_r,temp_m2_3_2_i,temp_m2_3_4_r,temp_m2_3_4_i,temp_b2_1_2_r,temp_b2_1_2_i,temp_b2_1_4_r,temp_b2_1_4_i,temp_b2_3_2_r,temp_b2_3_2_i,temp_b2_3_4_r,temp_b2_3_4_i);
MULT MULT259 (clk,temp_b1_2_1_r,temp_b1_2_1_i,temp_b1_2_3_r,temp_b1_2_3_i,temp_b1_4_1_r,temp_b1_4_1_i,temp_b1_4_3_r,temp_b1_4_3_i,temp_m2_2_1_r,temp_m2_2_1_i,temp_m2_2_3_r,temp_m2_2_3_i,temp_m2_4_1_r,temp_m2_4_1_i,temp_m2_4_3_r,temp_m2_4_3_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly259 (clk,temp_m2_2_1_r,temp_m2_2_1_i,temp_m2_2_3_r,temp_m2_2_3_i,temp_m2_4_1_r,temp_m2_4_1_i,temp_m2_4_3_r,temp_m2_4_3_i,temp_b2_2_1_r,temp_b2_2_1_i,temp_b2_2_3_r,temp_b2_2_3_i,temp_b2_4_1_r,temp_b2_4_1_i,temp_b2_4_3_r,temp_b2_4_3_i);
MULT MULT260 (clk,temp_b1_2_2_r,temp_b1_2_2_i,temp_b1_2_4_r,temp_b1_2_4_i,temp_b1_4_2_r,temp_b1_4_2_i,temp_b1_4_4_r,temp_b1_4_4_i,temp_m2_2_2_r,temp_m2_2_2_i,temp_m2_2_4_r,temp_m2_2_4_i,temp_m2_4_2_r,temp_m2_4_2_i,temp_m2_4_4_r,temp_m2_4_4_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly260 (clk,temp_m2_2_2_r,temp_m2_2_2_i,temp_m2_2_4_r,temp_m2_2_4_i,temp_m2_4_2_r,temp_m2_4_2_i,temp_m2_4_4_r,temp_m2_4_4_i,temp_b2_2_2_r,temp_b2_2_2_i,temp_b2_2_4_r,temp_b2_2_4_i,temp_b2_4_2_r,temp_b2_4_2_i,temp_b2_4_4_r,temp_b2_4_4_i);
MULT MULT261 (clk,temp_b1_1_5_r,temp_b1_1_5_i,temp_b1_1_7_r,temp_b1_1_7_i,temp_b1_3_5_r,temp_b1_3_5_i,temp_b1_3_7_r,temp_b1_3_7_i,temp_m2_1_5_r,temp_m2_1_5_i,temp_m2_1_7_r,temp_m2_1_7_i,temp_m2_3_5_r,temp_m2_3_5_i,temp_m2_3_7_r,temp_m2_3_7_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly261 (clk,temp_m2_1_5_r,temp_m2_1_5_i,temp_m2_1_7_r,temp_m2_1_7_i,temp_m2_3_5_r,temp_m2_3_5_i,temp_m2_3_7_r,temp_m2_3_7_i,temp_b2_1_5_r,temp_b2_1_5_i,temp_b2_1_7_r,temp_b2_1_7_i,temp_b2_3_5_r,temp_b2_3_5_i,temp_b2_3_7_r,temp_b2_3_7_i);
MULT MULT262 (clk,temp_b1_1_6_r,temp_b1_1_6_i,temp_b1_1_8_r,temp_b1_1_8_i,temp_b1_3_6_r,temp_b1_3_6_i,temp_b1_3_8_r,temp_b1_3_8_i,temp_m2_1_6_r,temp_m2_1_6_i,temp_m2_1_8_r,temp_m2_1_8_i,temp_m2_3_6_r,temp_m2_3_6_i,temp_m2_3_8_r,temp_m2_3_8_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly262 (clk,temp_m2_1_6_r,temp_m2_1_6_i,temp_m2_1_8_r,temp_m2_1_8_i,temp_m2_3_6_r,temp_m2_3_6_i,temp_m2_3_8_r,temp_m2_3_8_i,temp_b2_1_6_r,temp_b2_1_6_i,temp_b2_1_8_r,temp_b2_1_8_i,temp_b2_3_6_r,temp_b2_3_6_i,temp_b2_3_8_r,temp_b2_3_8_i);
MULT MULT263 (clk,temp_b1_2_5_r,temp_b1_2_5_i,temp_b1_2_7_r,temp_b1_2_7_i,temp_b1_4_5_r,temp_b1_4_5_i,temp_b1_4_7_r,temp_b1_4_7_i,temp_m2_2_5_r,temp_m2_2_5_i,temp_m2_2_7_r,temp_m2_2_7_i,temp_m2_4_5_r,temp_m2_4_5_i,temp_m2_4_7_r,temp_m2_4_7_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly263 (clk,temp_m2_2_5_r,temp_m2_2_5_i,temp_m2_2_7_r,temp_m2_2_7_i,temp_m2_4_5_r,temp_m2_4_5_i,temp_m2_4_7_r,temp_m2_4_7_i,temp_b2_2_5_r,temp_b2_2_5_i,temp_b2_2_7_r,temp_b2_2_7_i,temp_b2_4_5_r,temp_b2_4_5_i,temp_b2_4_7_r,temp_b2_4_7_i);
MULT MULT264 (clk,temp_b1_2_6_r,temp_b1_2_6_i,temp_b1_2_8_r,temp_b1_2_8_i,temp_b1_4_6_r,temp_b1_4_6_i,temp_b1_4_8_r,temp_b1_4_8_i,temp_m2_2_6_r,temp_m2_2_6_i,temp_m2_2_8_r,temp_m2_2_8_i,temp_m2_4_6_r,temp_m2_4_6_i,temp_m2_4_8_r,temp_m2_4_8_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly264 (clk,temp_m2_2_6_r,temp_m2_2_6_i,temp_m2_2_8_r,temp_m2_2_8_i,temp_m2_4_6_r,temp_m2_4_6_i,temp_m2_4_8_r,temp_m2_4_8_i,temp_b2_2_6_r,temp_b2_2_6_i,temp_b2_2_8_r,temp_b2_2_8_i,temp_b2_4_6_r,temp_b2_4_6_i,temp_b2_4_8_r,temp_b2_4_8_i);
MULT MULT265 (clk,temp_b1_1_9_r,temp_b1_1_9_i,temp_b1_1_11_r,temp_b1_1_11_i,temp_b1_3_9_r,temp_b1_3_9_i,temp_b1_3_11_r,temp_b1_3_11_i,temp_m2_1_9_r,temp_m2_1_9_i,temp_m2_1_11_r,temp_m2_1_11_i,temp_m2_3_9_r,temp_m2_3_9_i,temp_m2_3_11_r,temp_m2_3_11_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly265 (clk,temp_m2_1_9_r,temp_m2_1_9_i,temp_m2_1_11_r,temp_m2_1_11_i,temp_m2_3_9_r,temp_m2_3_9_i,temp_m2_3_11_r,temp_m2_3_11_i,temp_b2_1_9_r,temp_b2_1_9_i,temp_b2_1_11_r,temp_b2_1_11_i,temp_b2_3_9_r,temp_b2_3_9_i,temp_b2_3_11_r,temp_b2_3_11_i);
MULT MULT266 (clk,temp_b1_1_10_r,temp_b1_1_10_i,temp_b1_1_12_r,temp_b1_1_12_i,temp_b1_3_10_r,temp_b1_3_10_i,temp_b1_3_12_r,temp_b1_3_12_i,temp_m2_1_10_r,temp_m2_1_10_i,temp_m2_1_12_r,temp_m2_1_12_i,temp_m2_3_10_r,temp_m2_3_10_i,temp_m2_3_12_r,temp_m2_3_12_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly266 (clk,temp_m2_1_10_r,temp_m2_1_10_i,temp_m2_1_12_r,temp_m2_1_12_i,temp_m2_3_10_r,temp_m2_3_10_i,temp_m2_3_12_r,temp_m2_3_12_i,temp_b2_1_10_r,temp_b2_1_10_i,temp_b2_1_12_r,temp_b2_1_12_i,temp_b2_3_10_r,temp_b2_3_10_i,temp_b2_3_12_r,temp_b2_3_12_i);
MULT MULT267 (clk,temp_b1_2_9_r,temp_b1_2_9_i,temp_b1_2_11_r,temp_b1_2_11_i,temp_b1_4_9_r,temp_b1_4_9_i,temp_b1_4_11_r,temp_b1_4_11_i,temp_m2_2_9_r,temp_m2_2_9_i,temp_m2_2_11_r,temp_m2_2_11_i,temp_m2_4_9_r,temp_m2_4_9_i,temp_m2_4_11_r,temp_m2_4_11_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly267 (clk,temp_m2_2_9_r,temp_m2_2_9_i,temp_m2_2_11_r,temp_m2_2_11_i,temp_m2_4_9_r,temp_m2_4_9_i,temp_m2_4_11_r,temp_m2_4_11_i,temp_b2_2_9_r,temp_b2_2_9_i,temp_b2_2_11_r,temp_b2_2_11_i,temp_b2_4_9_r,temp_b2_4_9_i,temp_b2_4_11_r,temp_b2_4_11_i);
MULT MULT268 (clk,temp_b1_2_10_r,temp_b1_2_10_i,temp_b1_2_12_r,temp_b1_2_12_i,temp_b1_4_10_r,temp_b1_4_10_i,temp_b1_4_12_r,temp_b1_4_12_i,temp_m2_2_10_r,temp_m2_2_10_i,temp_m2_2_12_r,temp_m2_2_12_i,temp_m2_4_10_r,temp_m2_4_10_i,temp_m2_4_12_r,temp_m2_4_12_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly268 (clk,temp_m2_2_10_r,temp_m2_2_10_i,temp_m2_2_12_r,temp_m2_2_12_i,temp_m2_4_10_r,temp_m2_4_10_i,temp_m2_4_12_r,temp_m2_4_12_i,temp_b2_2_10_r,temp_b2_2_10_i,temp_b2_2_12_r,temp_b2_2_12_i,temp_b2_4_10_r,temp_b2_4_10_i,temp_b2_4_12_r,temp_b2_4_12_i);
MULT MULT269 (clk,temp_b1_1_13_r,temp_b1_1_13_i,temp_b1_1_15_r,temp_b1_1_15_i,temp_b1_3_13_r,temp_b1_3_13_i,temp_b1_3_15_r,temp_b1_3_15_i,temp_m2_1_13_r,temp_m2_1_13_i,temp_m2_1_15_r,temp_m2_1_15_i,temp_m2_3_13_r,temp_m2_3_13_i,temp_m2_3_15_r,temp_m2_3_15_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly269 (clk,temp_m2_1_13_r,temp_m2_1_13_i,temp_m2_1_15_r,temp_m2_1_15_i,temp_m2_3_13_r,temp_m2_3_13_i,temp_m2_3_15_r,temp_m2_3_15_i,temp_b2_1_13_r,temp_b2_1_13_i,temp_b2_1_15_r,temp_b2_1_15_i,temp_b2_3_13_r,temp_b2_3_13_i,temp_b2_3_15_r,temp_b2_3_15_i);
MULT MULT270 (clk,temp_b1_1_14_r,temp_b1_1_14_i,temp_b1_1_16_r,temp_b1_1_16_i,temp_b1_3_14_r,temp_b1_3_14_i,temp_b1_3_16_r,temp_b1_3_16_i,temp_m2_1_14_r,temp_m2_1_14_i,temp_m2_1_16_r,temp_m2_1_16_i,temp_m2_3_14_r,temp_m2_3_14_i,temp_m2_3_16_r,temp_m2_3_16_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly270 (clk,temp_m2_1_14_r,temp_m2_1_14_i,temp_m2_1_16_r,temp_m2_1_16_i,temp_m2_3_14_r,temp_m2_3_14_i,temp_m2_3_16_r,temp_m2_3_16_i,temp_b2_1_14_r,temp_b2_1_14_i,temp_b2_1_16_r,temp_b2_1_16_i,temp_b2_3_14_r,temp_b2_3_14_i,temp_b2_3_16_r,temp_b2_3_16_i);
MULT MULT271 (clk,temp_b1_2_13_r,temp_b1_2_13_i,temp_b1_2_15_r,temp_b1_2_15_i,temp_b1_4_13_r,temp_b1_4_13_i,temp_b1_4_15_r,temp_b1_4_15_i,temp_m2_2_13_r,temp_m2_2_13_i,temp_m2_2_15_r,temp_m2_2_15_i,temp_m2_4_13_r,temp_m2_4_13_i,temp_m2_4_15_r,temp_m2_4_15_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly271 (clk,temp_m2_2_13_r,temp_m2_2_13_i,temp_m2_2_15_r,temp_m2_2_15_i,temp_m2_4_13_r,temp_m2_4_13_i,temp_m2_4_15_r,temp_m2_4_15_i,temp_b2_2_13_r,temp_b2_2_13_i,temp_b2_2_15_r,temp_b2_2_15_i,temp_b2_4_13_r,temp_b2_4_13_i,temp_b2_4_15_r,temp_b2_4_15_i);
MULT MULT272 (clk,temp_b1_2_14_r,temp_b1_2_14_i,temp_b1_2_16_r,temp_b1_2_16_i,temp_b1_4_14_r,temp_b1_4_14_i,temp_b1_4_16_r,temp_b1_4_16_i,temp_m2_2_14_r,temp_m2_2_14_i,temp_m2_2_16_r,temp_m2_2_16_i,temp_m2_4_14_r,temp_m2_4_14_i,temp_m2_4_16_r,temp_m2_4_16_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly272 (clk,temp_m2_2_14_r,temp_m2_2_14_i,temp_m2_2_16_r,temp_m2_2_16_i,temp_m2_4_14_r,temp_m2_4_14_i,temp_m2_4_16_r,temp_m2_4_16_i,temp_b2_2_14_r,temp_b2_2_14_i,temp_b2_2_16_r,temp_b2_2_16_i,temp_b2_4_14_r,temp_b2_4_14_i,temp_b2_4_16_r,temp_b2_4_16_i);
MULT MULT273 (clk,temp_b1_1_17_r,temp_b1_1_17_i,temp_b1_1_19_r,temp_b1_1_19_i,temp_b1_3_17_r,temp_b1_3_17_i,temp_b1_3_19_r,temp_b1_3_19_i,temp_m2_1_17_r,temp_m2_1_17_i,temp_m2_1_19_r,temp_m2_1_19_i,temp_m2_3_17_r,temp_m2_3_17_i,temp_m2_3_19_r,temp_m2_3_19_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly273 (clk,temp_m2_1_17_r,temp_m2_1_17_i,temp_m2_1_19_r,temp_m2_1_19_i,temp_m2_3_17_r,temp_m2_3_17_i,temp_m2_3_19_r,temp_m2_3_19_i,temp_b2_1_17_r,temp_b2_1_17_i,temp_b2_1_19_r,temp_b2_1_19_i,temp_b2_3_17_r,temp_b2_3_17_i,temp_b2_3_19_r,temp_b2_3_19_i);
MULT MULT274 (clk,temp_b1_1_18_r,temp_b1_1_18_i,temp_b1_1_20_r,temp_b1_1_20_i,temp_b1_3_18_r,temp_b1_3_18_i,temp_b1_3_20_r,temp_b1_3_20_i,temp_m2_1_18_r,temp_m2_1_18_i,temp_m2_1_20_r,temp_m2_1_20_i,temp_m2_3_18_r,temp_m2_3_18_i,temp_m2_3_20_r,temp_m2_3_20_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly274 (clk,temp_m2_1_18_r,temp_m2_1_18_i,temp_m2_1_20_r,temp_m2_1_20_i,temp_m2_3_18_r,temp_m2_3_18_i,temp_m2_3_20_r,temp_m2_3_20_i,temp_b2_1_18_r,temp_b2_1_18_i,temp_b2_1_20_r,temp_b2_1_20_i,temp_b2_3_18_r,temp_b2_3_18_i,temp_b2_3_20_r,temp_b2_3_20_i);
MULT MULT275 (clk,temp_b1_2_17_r,temp_b1_2_17_i,temp_b1_2_19_r,temp_b1_2_19_i,temp_b1_4_17_r,temp_b1_4_17_i,temp_b1_4_19_r,temp_b1_4_19_i,temp_m2_2_17_r,temp_m2_2_17_i,temp_m2_2_19_r,temp_m2_2_19_i,temp_m2_4_17_r,temp_m2_4_17_i,temp_m2_4_19_r,temp_m2_4_19_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly275 (clk,temp_m2_2_17_r,temp_m2_2_17_i,temp_m2_2_19_r,temp_m2_2_19_i,temp_m2_4_17_r,temp_m2_4_17_i,temp_m2_4_19_r,temp_m2_4_19_i,temp_b2_2_17_r,temp_b2_2_17_i,temp_b2_2_19_r,temp_b2_2_19_i,temp_b2_4_17_r,temp_b2_4_17_i,temp_b2_4_19_r,temp_b2_4_19_i);
MULT MULT276 (clk,temp_b1_2_18_r,temp_b1_2_18_i,temp_b1_2_20_r,temp_b1_2_20_i,temp_b1_4_18_r,temp_b1_4_18_i,temp_b1_4_20_r,temp_b1_4_20_i,temp_m2_2_18_r,temp_m2_2_18_i,temp_m2_2_20_r,temp_m2_2_20_i,temp_m2_4_18_r,temp_m2_4_18_i,temp_m2_4_20_r,temp_m2_4_20_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly276 (clk,temp_m2_2_18_r,temp_m2_2_18_i,temp_m2_2_20_r,temp_m2_2_20_i,temp_m2_4_18_r,temp_m2_4_18_i,temp_m2_4_20_r,temp_m2_4_20_i,temp_b2_2_18_r,temp_b2_2_18_i,temp_b2_2_20_r,temp_b2_2_20_i,temp_b2_4_18_r,temp_b2_4_18_i,temp_b2_4_20_r,temp_b2_4_20_i);
MULT MULT277 (clk,temp_b1_1_21_r,temp_b1_1_21_i,temp_b1_1_23_r,temp_b1_1_23_i,temp_b1_3_21_r,temp_b1_3_21_i,temp_b1_3_23_r,temp_b1_3_23_i,temp_m2_1_21_r,temp_m2_1_21_i,temp_m2_1_23_r,temp_m2_1_23_i,temp_m2_3_21_r,temp_m2_3_21_i,temp_m2_3_23_r,temp_m2_3_23_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly277 (clk,temp_m2_1_21_r,temp_m2_1_21_i,temp_m2_1_23_r,temp_m2_1_23_i,temp_m2_3_21_r,temp_m2_3_21_i,temp_m2_3_23_r,temp_m2_3_23_i,temp_b2_1_21_r,temp_b2_1_21_i,temp_b2_1_23_r,temp_b2_1_23_i,temp_b2_3_21_r,temp_b2_3_21_i,temp_b2_3_23_r,temp_b2_3_23_i);
MULT MULT278 (clk,temp_b1_1_22_r,temp_b1_1_22_i,temp_b1_1_24_r,temp_b1_1_24_i,temp_b1_3_22_r,temp_b1_3_22_i,temp_b1_3_24_r,temp_b1_3_24_i,temp_m2_1_22_r,temp_m2_1_22_i,temp_m2_1_24_r,temp_m2_1_24_i,temp_m2_3_22_r,temp_m2_3_22_i,temp_m2_3_24_r,temp_m2_3_24_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly278 (clk,temp_m2_1_22_r,temp_m2_1_22_i,temp_m2_1_24_r,temp_m2_1_24_i,temp_m2_3_22_r,temp_m2_3_22_i,temp_m2_3_24_r,temp_m2_3_24_i,temp_b2_1_22_r,temp_b2_1_22_i,temp_b2_1_24_r,temp_b2_1_24_i,temp_b2_3_22_r,temp_b2_3_22_i,temp_b2_3_24_r,temp_b2_3_24_i);
MULT MULT279 (clk,temp_b1_2_21_r,temp_b1_2_21_i,temp_b1_2_23_r,temp_b1_2_23_i,temp_b1_4_21_r,temp_b1_4_21_i,temp_b1_4_23_r,temp_b1_4_23_i,temp_m2_2_21_r,temp_m2_2_21_i,temp_m2_2_23_r,temp_m2_2_23_i,temp_m2_4_21_r,temp_m2_4_21_i,temp_m2_4_23_r,temp_m2_4_23_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly279 (clk,temp_m2_2_21_r,temp_m2_2_21_i,temp_m2_2_23_r,temp_m2_2_23_i,temp_m2_4_21_r,temp_m2_4_21_i,temp_m2_4_23_r,temp_m2_4_23_i,temp_b2_2_21_r,temp_b2_2_21_i,temp_b2_2_23_r,temp_b2_2_23_i,temp_b2_4_21_r,temp_b2_4_21_i,temp_b2_4_23_r,temp_b2_4_23_i);
MULT MULT280 (clk,temp_b1_2_22_r,temp_b1_2_22_i,temp_b1_2_24_r,temp_b1_2_24_i,temp_b1_4_22_r,temp_b1_4_22_i,temp_b1_4_24_r,temp_b1_4_24_i,temp_m2_2_22_r,temp_m2_2_22_i,temp_m2_2_24_r,temp_m2_2_24_i,temp_m2_4_22_r,temp_m2_4_22_i,temp_m2_4_24_r,temp_m2_4_24_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly280 (clk,temp_m2_2_22_r,temp_m2_2_22_i,temp_m2_2_24_r,temp_m2_2_24_i,temp_m2_4_22_r,temp_m2_4_22_i,temp_m2_4_24_r,temp_m2_4_24_i,temp_b2_2_22_r,temp_b2_2_22_i,temp_b2_2_24_r,temp_b2_2_24_i,temp_b2_4_22_r,temp_b2_4_22_i,temp_b2_4_24_r,temp_b2_4_24_i);
MULT MULT281 (clk,temp_b1_1_25_r,temp_b1_1_25_i,temp_b1_1_27_r,temp_b1_1_27_i,temp_b1_3_25_r,temp_b1_3_25_i,temp_b1_3_27_r,temp_b1_3_27_i,temp_m2_1_25_r,temp_m2_1_25_i,temp_m2_1_27_r,temp_m2_1_27_i,temp_m2_3_25_r,temp_m2_3_25_i,temp_m2_3_27_r,temp_m2_3_27_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly281 (clk,temp_m2_1_25_r,temp_m2_1_25_i,temp_m2_1_27_r,temp_m2_1_27_i,temp_m2_3_25_r,temp_m2_3_25_i,temp_m2_3_27_r,temp_m2_3_27_i,temp_b2_1_25_r,temp_b2_1_25_i,temp_b2_1_27_r,temp_b2_1_27_i,temp_b2_3_25_r,temp_b2_3_25_i,temp_b2_3_27_r,temp_b2_3_27_i);
MULT MULT282 (clk,temp_b1_1_26_r,temp_b1_1_26_i,temp_b1_1_28_r,temp_b1_1_28_i,temp_b1_3_26_r,temp_b1_3_26_i,temp_b1_3_28_r,temp_b1_3_28_i,temp_m2_1_26_r,temp_m2_1_26_i,temp_m2_1_28_r,temp_m2_1_28_i,temp_m2_3_26_r,temp_m2_3_26_i,temp_m2_3_28_r,temp_m2_3_28_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly282 (clk,temp_m2_1_26_r,temp_m2_1_26_i,temp_m2_1_28_r,temp_m2_1_28_i,temp_m2_3_26_r,temp_m2_3_26_i,temp_m2_3_28_r,temp_m2_3_28_i,temp_b2_1_26_r,temp_b2_1_26_i,temp_b2_1_28_r,temp_b2_1_28_i,temp_b2_3_26_r,temp_b2_3_26_i,temp_b2_3_28_r,temp_b2_3_28_i);
MULT MULT283 (clk,temp_b1_2_25_r,temp_b1_2_25_i,temp_b1_2_27_r,temp_b1_2_27_i,temp_b1_4_25_r,temp_b1_4_25_i,temp_b1_4_27_r,temp_b1_4_27_i,temp_m2_2_25_r,temp_m2_2_25_i,temp_m2_2_27_r,temp_m2_2_27_i,temp_m2_4_25_r,temp_m2_4_25_i,temp_m2_4_27_r,temp_m2_4_27_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly283 (clk,temp_m2_2_25_r,temp_m2_2_25_i,temp_m2_2_27_r,temp_m2_2_27_i,temp_m2_4_25_r,temp_m2_4_25_i,temp_m2_4_27_r,temp_m2_4_27_i,temp_b2_2_25_r,temp_b2_2_25_i,temp_b2_2_27_r,temp_b2_2_27_i,temp_b2_4_25_r,temp_b2_4_25_i,temp_b2_4_27_r,temp_b2_4_27_i);
MULT MULT284 (clk,temp_b1_2_26_r,temp_b1_2_26_i,temp_b1_2_28_r,temp_b1_2_28_i,temp_b1_4_26_r,temp_b1_4_26_i,temp_b1_4_28_r,temp_b1_4_28_i,temp_m2_2_26_r,temp_m2_2_26_i,temp_m2_2_28_r,temp_m2_2_28_i,temp_m2_4_26_r,temp_m2_4_26_i,temp_m2_4_28_r,temp_m2_4_28_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly284 (clk,temp_m2_2_26_r,temp_m2_2_26_i,temp_m2_2_28_r,temp_m2_2_28_i,temp_m2_4_26_r,temp_m2_4_26_i,temp_m2_4_28_r,temp_m2_4_28_i,temp_b2_2_26_r,temp_b2_2_26_i,temp_b2_2_28_r,temp_b2_2_28_i,temp_b2_4_26_r,temp_b2_4_26_i,temp_b2_4_28_r,temp_b2_4_28_i);
MULT MULT285 (clk,temp_b1_1_29_r,temp_b1_1_29_i,temp_b1_1_31_r,temp_b1_1_31_i,temp_b1_3_29_r,temp_b1_3_29_i,temp_b1_3_31_r,temp_b1_3_31_i,temp_m2_1_29_r,temp_m2_1_29_i,temp_m2_1_31_r,temp_m2_1_31_i,temp_m2_3_29_r,temp_m2_3_29_i,temp_m2_3_31_r,temp_m2_3_31_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly285 (clk,temp_m2_1_29_r,temp_m2_1_29_i,temp_m2_1_31_r,temp_m2_1_31_i,temp_m2_3_29_r,temp_m2_3_29_i,temp_m2_3_31_r,temp_m2_3_31_i,temp_b2_1_29_r,temp_b2_1_29_i,temp_b2_1_31_r,temp_b2_1_31_i,temp_b2_3_29_r,temp_b2_3_29_i,temp_b2_3_31_r,temp_b2_3_31_i);
MULT MULT286 (clk,temp_b1_1_30_r,temp_b1_1_30_i,temp_b1_1_32_r,temp_b1_1_32_i,temp_b1_3_30_r,temp_b1_3_30_i,temp_b1_3_32_r,temp_b1_3_32_i,temp_m2_1_30_r,temp_m2_1_30_i,temp_m2_1_32_r,temp_m2_1_32_i,temp_m2_3_30_r,temp_m2_3_30_i,temp_m2_3_32_r,temp_m2_3_32_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly286 (clk,temp_m2_1_30_r,temp_m2_1_30_i,temp_m2_1_32_r,temp_m2_1_32_i,temp_m2_3_30_r,temp_m2_3_30_i,temp_m2_3_32_r,temp_m2_3_32_i,temp_b2_1_30_r,temp_b2_1_30_i,temp_b2_1_32_r,temp_b2_1_32_i,temp_b2_3_30_r,temp_b2_3_30_i,temp_b2_3_32_r,temp_b2_3_32_i);
MULT MULT287 (clk,temp_b1_2_29_r,temp_b1_2_29_i,temp_b1_2_31_r,temp_b1_2_31_i,temp_b1_4_29_r,temp_b1_4_29_i,temp_b1_4_31_r,temp_b1_4_31_i,temp_m2_2_29_r,temp_m2_2_29_i,temp_m2_2_31_r,temp_m2_2_31_i,temp_m2_4_29_r,temp_m2_4_29_i,temp_m2_4_31_r,temp_m2_4_31_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly287 (clk,temp_m2_2_29_r,temp_m2_2_29_i,temp_m2_2_31_r,temp_m2_2_31_i,temp_m2_4_29_r,temp_m2_4_29_i,temp_m2_4_31_r,temp_m2_4_31_i,temp_b2_2_29_r,temp_b2_2_29_i,temp_b2_2_31_r,temp_b2_2_31_i,temp_b2_4_29_r,temp_b2_4_29_i,temp_b2_4_31_r,temp_b2_4_31_i);
MULT MULT288 (clk,temp_b1_2_30_r,temp_b1_2_30_i,temp_b1_2_32_r,temp_b1_2_32_i,temp_b1_4_30_r,temp_b1_4_30_i,temp_b1_4_32_r,temp_b1_4_32_i,temp_m2_2_30_r,temp_m2_2_30_i,temp_m2_2_32_r,temp_m2_2_32_i,temp_m2_4_30_r,temp_m2_4_30_i,temp_m2_4_32_r,temp_m2_4_32_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly288 (clk,temp_m2_2_30_r,temp_m2_2_30_i,temp_m2_2_32_r,temp_m2_2_32_i,temp_m2_4_30_r,temp_m2_4_30_i,temp_m2_4_32_r,temp_m2_4_32_i,temp_b2_2_30_r,temp_b2_2_30_i,temp_b2_2_32_r,temp_b2_2_32_i,temp_b2_4_30_r,temp_b2_4_30_i,temp_b2_4_32_r,temp_b2_4_32_i);
MULT MULT289 (clk,temp_b1_5_1_r,temp_b1_5_1_i,temp_b1_5_3_r,temp_b1_5_3_i,temp_b1_7_1_r,temp_b1_7_1_i,temp_b1_7_3_r,temp_b1_7_3_i,temp_m2_5_1_r,temp_m2_5_1_i,temp_m2_5_3_r,temp_m2_5_3_i,temp_m2_7_1_r,temp_m2_7_1_i,temp_m2_7_3_r,temp_m2_7_3_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly289 (clk,temp_m2_5_1_r,temp_m2_5_1_i,temp_m2_5_3_r,temp_m2_5_3_i,temp_m2_7_1_r,temp_m2_7_1_i,temp_m2_7_3_r,temp_m2_7_3_i,temp_b2_5_1_r,temp_b2_5_1_i,temp_b2_5_3_r,temp_b2_5_3_i,temp_b2_7_1_r,temp_b2_7_1_i,temp_b2_7_3_r,temp_b2_7_3_i);
MULT MULT290 (clk,temp_b1_5_2_r,temp_b1_5_2_i,temp_b1_5_4_r,temp_b1_5_4_i,temp_b1_7_2_r,temp_b1_7_2_i,temp_b1_7_4_r,temp_b1_7_4_i,temp_m2_5_2_r,temp_m2_5_2_i,temp_m2_5_4_r,temp_m2_5_4_i,temp_m2_7_2_r,temp_m2_7_2_i,temp_m2_7_4_r,temp_m2_7_4_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly290 (clk,temp_m2_5_2_r,temp_m2_5_2_i,temp_m2_5_4_r,temp_m2_5_4_i,temp_m2_7_2_r,temp_m2_7_2_i,temp_m2_7_4_r,temp_m2_7_4_i,temp_b2_5_2_r,temp_b2_5_2_i,temp_b2_5_4_r,temp_b2_5_4_i,temp_b2_7_2_r,temp_b2_7_2_i,temp_b2_7_4_r,temp_b2_7_4_i);
MULT MULT291 (clk,temp_b1_6_1_r,temp_b1_6_1_i,temp_b1_6_3_r,temp_b1_6_3_i,temp_b1_8_1_r,temp_b1_8_1_i,temp_b1_8_3_r,temp_b1_8_3_i,temp_m2_6_1_r,temp_m2_6_1_i,temp_m2_6_3_r,temp_m2_6_3_i,temp_m2_8_1_r,temp_m2_8_1_i,temp_m2_8_3_r,temp_m2_8_3_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly291 (clk,temp_m2_6_1_r,temp_m2_6_1_i,temp_m2_6_3_r,temp_m2_6_3_i,temp_m2_8_1_r,temp_m2_8_1_i,temp_m2_8_3_r,temp_m2_8_3_i,temp_b2_6_1_r,temp_b2_6_1_i,temp_b2_6_3_r,temp_b2_6_3_i,temp_b2_8_1_r,temp_b2_8_1_i,temp_b2_8_3_r,temp_b2_8_3_i);
MULT MULT292 (clk,temp_b1_6_2_r,temp_b1_6_2_i,temp_b1_6_4_r,temp_b1_6_4_i,temp_b1_8_2_r,temp_b1_8_2_i,temp_b1_8_4_r,temp_b1_8_4_i,temp_m2_6_2_r,temp_m2_6_2_i,temp_m2_6_4_r,temp_m2_6_4_i,temp_m2_8_2_r,temp_m2_8_2_i,temp_m2_8_4_r,temp_m2_8_4_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly292 (clk,temp_m2_6_2_r,temp_m2_6_2_i,temp_m2_6_4_r,temp_m2_6_4_i,temp_m2_8_2_r,temp_m2_8_2_i,temp_m2_8_4_r,temp_m2_8_4_i,temp_b2_6_2_r,temp_b2_6_2_i,temp_b2_6_4_r,temp_b2_6_4_i,temp_b2_8_2_r,temp_b2_8_2_i,temp_b2_8_4_r,temp_b2_8_4_i);
MULT MULT293 (clk,temp_b1_5_5_r,temp_b1_5_5_i,temp_b1_5_7_r,temp_b1_5_7_i,temp_b1_7_5_r,temp_b1_7_5_i,temp_b1_7_7_r,temp_b1_7_7_i,temp_m2_5_5_r,temp_m2_5_5_i,temp_m2_5_7_r,temp_m2_5_7_i,temp_m2_7_5_r,temp_m2_7_5_i,temp_m2_7_7_r,temp_m2_7_7_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly293 (clk,temp_m2_5_5_r,temp_m2_5_5_i,temp_m2_5_7_r,temp_m2_5_7_i,temp_m2_7_5_r,temp_m2_7_5_i,temp_m2_7_7_r,temp_m2_7_7_i,temp_b2_5_5_r,temp_b2_5_5_i,temp_b2_5_7_r,temp_b2_5_7_i,temp_b2_7_5_r,temp_b2_7_5_i,temp_b2_7_7_r,temp_b2_7_7_i);
MULT MULT294 (clk,temp_b1_5_6_r,temp_b1_5_6_i,temp_b1_5_8_r,temp_b1_5_8_i,temp_b1_7_6_r,temp_b1_7_6_i,temp_b1_7_8_r,temp_b1_7_8_i,temp_m2_5_6_r,temp_m2_5_6_i,temp_m2_5_8_r,temp_m2_5_8_i,temp_m2_7_6_r,temp_m2_7_6_i,temp_m2_7_8_r,temp_m2_7_8_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly294 (clk,temp_m2_5_6_r,temp_m2_5_6_i,temp_m2_5_8_r,temp_m2_5_8_i,temp_m2_7_6_r,temp_m2_7_6_i,temp_m2_7_8_r,temp_m2_7_8_i,temp_b2_5_6_r,temp_b2_5_6_i,temp_b2_5_8_r,temp_b2_5_8_i,temp_b2_7_6_r,temp_b2_7_6_i,temp_b2_7_8_r,temp_b2_7_8_i);
MULT MULT295 (clk,temp_b1_6_5_r,temp_b1_6_5_i,temp_b1_6_7_r,temp_b1_6_7_i,temp_b1_8_5_r,temp_b1_8_5_i,temp_b1_8_7_r,temp_b1_8_7_i,temp_m2_6_5_r,temp_m2_6_5_i,temp_m2_6_7_r,temp_m2_6_7_i,temp_m2_8_5_r,temp_m2_8_5_i,temp_m2_8_7_r,temp_m2_8_7_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly295 (clk,temp_m2_6_5_r,temp_m2_6_5_i,temp_m2_6_7_r,temp_m2_6_7_i,temp_m2_8_5_r,temp_m2_8_5_i,temp_m2_8_7_r,temp_m2_8_7_i,temp_b2_6_5_r,temp_b2_6_5_i,temp_b2_6_7_r,temp_b2_6_7_i,temp_b2_8_5_r,temp_b2_8_5_i,temp_b2_8_7_r,temp_b2_8_7_i);
MULT MULT296 (clk,temp_b1_6_6_r,temp_b1_6_6_i,temp_b1_6_8_r,temp_b1_6_8_i,temp_b1_8_6_r,temp_b1_8_6_i,temp_b1_8_8_r,temp_b1_8_8_i,temp_m2_6_6_r,temp_m2_6_6_i,temp_m2_6_8_r,temp_m2_6_8_i,temp_m2_8_6_r,temp_m2_8_6_i,temp_m2_8_8_r,temp_m2_8_8_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly296 (clk,temp_m2_6_6_r,temp_m2_6_6_i,temp_m2_6_8_r,temp_m2_6_8_i,temp_m2_8_6_r,temp_m2_8_6_i,temp_m2_8_8_r,temp_m2_8_8_i,temp_b2_6_6_r,temp_b2_6_6_i,temp_b2_6_8_r,temp_b2_6_8_i,temp_b2_8_6_r,temp_b2_8_6_i,temp_b2_8_8_r,temp_b2_8_8_i);
MULT MULT297 (clk,temp_b1_5_9_r,temp_b1_5_9_i,temp_b1_5_11_r,temp_b1_5_11_i,temp_b1_7_9_r,temp_b1_7_9_i,temp_b1_7_11_r,temp_b1_7_11_i,temp_m2_5_9_r,temp_m2_5_9_i,temp_m2_5_11_r,temp_m2_5_11_i,temp_m2_7_9_r,temp_m2_7_9_i,temp_m2_7_11_r,temp_m2_7_11_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly297 (clk,temp_m2_5_9_r,temp_m2_5_9_i,temp_m2_5_11_r,temp_m2_5_11_i,temp_m2_7_9_r,temp_m2_7_9_i,temp_m2_7_11_r,temp_m2_7_11_i,temp_b2_5_9_r,temp_b2_5_9_i,temp_b2_5_11_r,temp_b2_5_11_i,temp_b2_7_9_r,temp_b2_7_9_i,temp_b2_7_11_r,temp_b2_7_11_i);
MULT MULT298 (clk,temp_b1_5_10_r,temp_b1_5_10_i,temp_b1_5_12_r,temp_b1_5_12_i,temp_b1_7_10_r,temp_b1_7_10_i,temp_b1_7_12_r,temp_b1_7_12_i,temp_m2_5_10_r,temp_m2_5_10_i,temp_m2_5_12_r,temp_m2_5_12_i,temp_m2_7_10_r,temp_m2_7_10_i,temp_m2_7_12_r,temp_m2_7_12_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly298 (clk,temp_m2_5_10_r,temp_m2_5_10_i,temp_m2_5_12_r,temp_m2_5_12_i,temp_m2_7_10_r,temp_m2_7_10_i,temp_m2_7_12_r,temp_m2_7_12_i,temp_b2_5_10_r,temp_b2_5_10_i,temp_b2_5_12_r,temp_b2_5_12_i,temp_b2_7_10_r,temp_b2_7_10_i,temp_b2_7_12_r,temp_b2_7_12_i);
MULT MULT299 (clk,temp_b1_6_9_r,temp_b1_6_9_i,temp_b1_6_11_r,temp_b1_6_11_i,temp_b1_8_9_r,temp_b1_8_9_i,temp_b1_8_11_r,temp_b1_8_11_i,temp_m2_6_9_r,temp_m2_6_9_i,temp_m2_6_11_r,temp_m2_6_11_i,temp_m2_8_9_r,temp_m2_8_9_i,temp_m2_8_11_r,temp_m2_8_11_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly299 (clk,temp_m2_6_9_r,temp_m2_6_9_i,temp_m2_6_11_r,temp_m2_6_11_i,temp_m2_8_9_r,temp_m2_8_9_i,temp_m2_8_11_r,temp_m2_8_11_i,temp_b2_6_9_r,temp_b2_6_9_i,temp_b2_6_11_r,temp_b2_6_11_i,temp_b2_8_9_r,temp_b2_8_9_i,temp_b2_8_11_r,temp_b2_8_11_i);
MULT MULT300 (clk,temp_b1_6_10_r,temp_b1_6_10_i,temp_b1_6_12_r,temp_b1_6_12_i,temp_b1_8_10_r,temp_b1_8_10_i,temp_b1_8_12_r,temp_b1_8_12_i,temp_m2_6_10_r,temp_m2_6_10_i,temp_m2_6_12_r,temp_m2_6_12_i,temp_m2_8_10_r,temp_m2_8_10_i,temp_m2_8_12_r,temp_m2_8_12_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly300 (clk,temp_m2_6_10_r,temp_m2_6_10_i,temp_m2_6_12_r,temp_m2_6_12_i,temp_m2_8_10_r,temp_m2_8_10_i,temp_m2_8_12_r,temp_m2_8_12_i,temp_b2_6_10_r,temp_b2_6_10_i,temp_b2_6_12_r,temp_b2_6_12_i,temp_b2_8_10_r,temp_b2_8_10_i,temp_b2_8_12_r,temp_b2_8_12_i);
MULT MULT301 (clk,temp_b1_5_13_r,temp_b1_5_13_i,temp_b1_5_15_r,temp_b1_5_15_i,temp_b1_7_13_r,temp_b1_7_13_i,temp_b1_7_15_r,temp_b1_7_15_i,temp_m2_5_13_r,temp_m2_5_13_i,temp_m2_5_15_r,temp_m2_5_15_i,temp_m2_7_13_r,temp_m2_7_13_i,temp_m2_7_15_r,temp_m2_7_15_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly301 (clk,temp_m2_5_13_r,temp_m2_5_13_i,temp_m2_5_15_r,temp_m2_5_15_i,temp_m2_7_13_r,temp_m2_7_13_i,temp_m2_7_15_r,temp_m2_7_15_i,temp_b2_5_13_r,temp_b2_5_13_i,temp_b2_5_15_r,temp_b2_5_15_i,temp_b2_7_13_r,temp_b2_7_13_i,temp_b2_7_15_r,temp_b2_7_15_i);
MULT MULT302 (clk,temp_b1_5_14_r,temp_b1_5_14_i,temp_b1_5_16_r,temp_b1_5_16_i,temp_b1_7_14_r,temp_b1_7_14_i,temp_b1_7_16_r,temp_b1_7_16_i,temp_m2_5_14_r,temp_m2_5_14_i,temp_m2_5_16_r,temp_m2_5_16_i,temp_m2_7_14_r,temp_m2_7_14_i,temp_m2_7_16_r,temp_m2_7_16_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly302 (clk,temp_m2_5_14_r,temp_m2_5_14_i,temp_m2_5_16_r,temp_m2_5_16_i,temp_m2_7_14_r,temp_m2_7_14_i,temp_m2_7_16_r,temp_m2_7_16_i,temp_b2_5_14_r,temp_b2_5_14_i,temp_b2_5_16_r,temp_b2_5_16_i,temp_b2_7_14_r,temp_b2_7_14_i,temp_b2_7_16_r,temp_b2_7_16_i);
MULT MULT303 (clk,temp_b1_6_13_r,temp_b1_6_13_i,temp_b1_6_15_r,temp_b1_6_15_i,temp_b1_8_13_r,temp_b1_8_13_i,temp_b1_8_15_r,temp_b1_8_15_i,temp_m2_6_13_r,temp_m2_6_13_i,temp_m2_6_15_r,temp_m2_6_15_i,temp_m2_8_13_r,temp_m2_8_13_i,temp_m2_8_15_r,temp_m2_8_15_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly303 (clk,temp_m2_6_13_r,temp_m2_6_13_i,temp_m2_6_15_r,temp_m2_6_15_i,temp_m2_8_13_r,temp_m2_8_13_i,temp_m2_8_15_r,temp_m2_8_15_i,temp_b2_6_13_r,temp_b2_6_13_i,temp_b2_6_15_r,temp_b2_6_15_i,temp_b2_8_13_r,temp_b2_8_13_i,temp_b2_8_15_r,temp_b2_8_15_i);
MULT MULT304 (clk,temp_b1_6_14_r,temp_b1_6_14_i,temp_b1_6_16_r,temp_b1_6_16_i,temp_b1_8_14_r,temp_b1_8_14_i,temp_b1_8_16_r,temp_b1_8_16_i,temp_m2_6_14_r,temp_m2_6_14_i,temp_m2_6_16_r,temp_m2_6_16_i,temp_m2_8_14_r,temp_m2_8_14_i,temp_m2_8_16_r,temp_m2_8_16_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly304 (clk,temp_m2_6_14_r,temp_m2_6_14_i,temp_m2_6_16_r,temp_m2_6_16_i,temp_m2_8_14_r,temp_m2_8_14_i,temp_m2_8_16_r,temp_m2_8_16_i,temp_b2_6_14_r,temp_b2_6_14_i,temp_b2_6_16_r,temp_b2_6_16_i,temp_b2_8_14_r,temp_b2_8_14_i,temp_b2_8_16_r,temp_b2_8_16_i);
MULT MULT305 (clk,temp_b1_5_17_r,temp_b1_5_17_i,temp_b1_5_19_r,temp_b1_5_19_i,temp_b1_7_17_r,temp_b1_7_17_i,temp_b1_7_19_r,temp_b1_7_19_i,temp_m2_5_17_r,temp_m2_5_17_i,temp_m2_5_19_r,temp_m2_5_19_i,temp_m2_7_17_r,temp_m2_7_17_i,temp_m2_7_19_r,temp_m2_7_19_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly305 (clk,temp_m2_5_17_r,temp_m2_5_17_i,temp_m2_5_19_r,temp_m2_5_19_i,temp_m2_7_17_r,temp_m2_7_17_i,temp_m2_7_19_r,temp_m2_7_19_i,temp_b2_5_17_r,temp_b2_5_17_i,temp_b2_5_19_r,temp_b2_5_19_i,temp_b2_7_17_r,temp_b2_7_17_i,temp_b2_7_19_r,temp_b2_7_19_i);
MULT MULT306 (clk,temp_b1_5_18_r,temp_b1_5_18_i,temp_b1_5_20_r,temp_b1_5_20_i,temp_b1_7_18_r,temp_b1_7_18_i,temp_b1_7_20_r,temp_b1_7_20_i,temp_m2_5_18_r,temp_m2_5_18_i,temp_m2_5_20_r,temp_m2_5_20_i,temp_m2_7_18_r,temp_m2_7_18_i,temp_m2_7_20_r,temp_m2_7_20_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly306 (clk,temp_m2_5_18_r,temp_m2_5_18_i,temp_m2_5_20_r,temp_m2_5_20_i,temp_m2_7_18_r,temp_m2_7_18_i,temp_m2_7_20_r,temp_m2_7_20_i,temp_b2_5_18_r,temp_b2_5_18_i,temp_b2_5_20_r,temp_b2_5_20_i,temp_b2_7_18_r,temp_b2_7_18_i,temp_b2_7_20_r,temp_b2_7_20_i);
MULT MULT307 (clk,temp_b1_6_17_r,temp_b1_6_17_i,temp_b1_6_19_r,temp_b1_6_19_i,temp_b1_8_17_r,temp_b1_8_17_i,temp_b1_8_19_r,temp_b1_8_19_i,temp_m2_6_17_r,temp_m2_6_17_i,temp_m2_6_19_r,temp_m2_6_19_i,temp_m2_8_17_r,temp_m2_8_17_i,temp_m2_8_19_r,temp_m2_8_19_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly307 (clk,temp_m2_6_17_r,temp_m2_6_17_i,temp_m2_6_19_r,temp_m2_6_19_i,temp_m2_8_17_r,temp_m2_8_17_i,temp_m2_8_19_r,temp_m2_8_19_i,temp_b2_6_17_r,temp_b2_6_17_i,temp_b2_6_19_r,temp_b2_6_19_i,temp_b2_8_17_r,temp_b2_8_17_i,temp_b2_8_19_r,temp_b2_8_19_i);
MULT MULT308 (clk,temp_b1_6_18_r,temp_b1_6_18_i,temp_b1_6_20_r,temp_b1_6_20_i,temp_b1_8_18_r,temp_b1_8_18_i,temp_b1_8_20_r,temp_b1_8_20_i,temp_m2_6_18_r,temp_m2_6_18_i,temp_m2_6_20_r,temp_m2_6_20_i,temp_m2_8_18_r,temp_m2_8_18_i,temp_m2_8_20_r,temp_m2_8_20_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly308 (clk,temp_m2_6_18_r,temp_m2_6_18_i,temp_m2_6_20_r,temp_m2_6_20_i,temp_m2_8_18_r,temp_m2_8_18_i,temp_m2_8_20_r,temp_m2_8_20_i,temp_b2_6_18_r,temp_b2_6_18_i,temp_b2_6_20_r,temp_b2_6_20_i,temp_b2_8_18_r,temp_b2_8_18_i,temp_b2_8_20_r,temp_b2_8_20_i);
MULT MULT309 (clk,temp_b1_5_21_r,temp_b1_5_21_i,temp_b1_5_23_r,temp_b1_5_23_i,temp_b1_7_21_r,temp_b1_7_21_i,temp_b1_7_23_r,temp_b1_7_23_i,temp_m2_5_21_r,temp_m2_5_21_i,temp_m2_5_23_r,temp_m2_5_23_i,temp_m2_7_21_r,temp_m2_7_21_i,temp_m2_7_23_r,temp_m2_7_23_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly309 (clk,temp_m2_5_21_r,temp_m2_5_21_i,temp_m2_5_23_r,temp_m2_5_23_i,temp_m2_7_21_r,temp_m2_7_21_i,temp_m2_7_23_r,temp_m2_7_23_i,temp_b2_5_21_r,temp_b2_5_21_i,temp_b2_5_23_r,temp_b2_5_23_i,temp_b2_7_21_r,temp_b2_7_21_i,temp_b2_7_23_r,temp_b2_7_23_i);
MULT MULT310 (clk,temp_b1_5_22_r,temp_b1_5_22_i,temp_b1_5_24_r,temp_b1_5_24_i,temp_b1_7_22_r,temp_b1_7_22_i,temp_b1_7_24_r,temp_b1_7_24_i,temp_m2_5_22_r,temp_m2_5_22_i,temp_m2_5_24_r,temp_m2_5_24_i,temp_m2_7_22_r,temp_m2_7_22_i,temp_m2_7_24_r,temp_m2_7_24_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly310 (clk,temp_m2_5_22_r,temp_m2_5_22_i,temp_m2_5_24_r,temp_m2_5_24_i,temp_m2_7_22_r,temp_m2_7_22_i,temp_m2_7_24_r,temp_m2_7_24_i,temp_b2_5_22_r,temp_b2_5_22_i,temp_b2_5_24_r,temp_b2_5_24_i,temp_b2_7_22_r,temp_b2_7_22_i,temp_b2_7_24_r,temp_b2_7_24_i);
MULT MULT311 (clk,temp_b1_6_21_r,temp_b1_6_21_i,temp_b1_6_23_r,temp_b1_6_23_i,temp_b1_8_21_r,temp_b1_8_21_i,temp_b1_8_23_r,temp_b1_8_23_i,temp_m2_6_21_r,temp_m2_6_21_i,temp_m2_6_23_r,temp_m2_6_23_i,temp_m2_8_21_r,temp_m2_8_21_i,temp_m2_8_23_r,temp_m2_8_23_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly311 (clk,temp_m2_6_21_r,temp_m2_6_21_i,temp_m2_6_23_r,temp_m2_6_23_i,temp_m2_8_21_r,temp_m2_8_21_i,temp_m2_8_23_r,temp_m2_8_23_i,temp_b2_6_21_r,temp_b2_6_21_i,temp_b2_6_23_r,temp_b2_6_23_i,temp_b2_8_21_r,temp_b2_8_21_i,temp_b2_8_23_r,temp_b2_8_23_i);
MULT MULT312 (clk,temp_b1_6_22_r,temp_b1_6_22_i,temp_b1_6_24_r,temp_b1_6_24_i,temp_b1_8_22_r,temp_b1_8_22_i,temp_b1_8_24_r,temp_b1_8_24_i,temp_m2_6_22_r,temp_m2_6_22_i,temp_m2_6_24_r,temp_m2_6_24_i,temp_m2_8_22_r,temp_m2_8_22_i,temp_m2_8_24_r,temp_m2_8_24_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly312 (clk,temp_m2_6_22_r,temp_m2_6_22_i,temp_m2_6_24_r,temp_m2_6_24_i,temp_m2_8_22_r,temp_m2_8_22_i,temp_m2_8_24_r,temp_m2_8_24_i,temp_b2_6_22_r,temp_b2_6_22_i,temp_b2_6_24_r,temp_b2_6_24_i,temp_b2_8_22_r,temp_b2_8_22_i,temp_b2_8_24_r,temp_b2_8_24_i);
MULT MULT313 (clk,temp_b1_5_25_r,temp_b1_5_25_i,temp_b1_5_27_r,temp_b1_5_27_i,temp_b1_7_25_r,temp_b1_7_25_i,temp_b1_7_27_r,temp_b1_7_27_i,temp_m2_5_25_r,temp_m2_5_25_i,temp_m2_5_27_r,temp_m2_5_27_i,temp_m2_7_25_r,temp_m2_7_25_i,temp_m2_7_27_r,temp_m2_7_27_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly313 (clk,temp_m2_5_25_r,temp_m2_5_25_i,temp_m2_5_27_r,temp_m2_5_27_i,temp_m2_7_25_r,temp_m2_7_25_i,temp_m2_7_27_r,temp_m2_7_27_i,temp_b2_5_25_r,temp_b2_5_25_i,temp_b2_5_27_r,temp_b2_5_27_i,temp_b2_7_25_r,temp_b2_7_25_i,temp_b2_7_27_r,temp_b2_7_27_i);
MULT MULT314 (clk,temp_b1_5_26_r,temp_b1_5_26_i,temp_b1_5_28_r,temp_b1_5_28_i,temp_b1_7_26_r,temp_b1_7_26_i,temp_b1_7_28_r,temp_b1_7_28_i,temp_m2_5_26_r,temp_m2_5_26_i,temp_m2_5_28_r,temp_m2_5_28_i,temp_m2_7_26_r,temp_m2_7_26_i,temp_m2_7_28_r,temp_m2_7_28_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly314 (clk,temp_m2_5_26_r,temp_m2_5_26_i,temp_m2_5_28_r,temp_m2_5_28_i,temp_m2_7_26_r,temp_m2_7_26_i,temp_m2_7_28_r,temp_m2_7_28_i,temp_b2_5_26_r,temp_b2_5_26_i,temp_b2_5_28_r,temp_b2_5_28_i,temp_b2_7_26_r,temp_b2_7_26_i,temp_b2_7_28_r,temp_b2_7_28_i);
MULT MULT315 (clk,temp_b1_6_25_r,temp_b1_6_25_i,temp_b1_6_27_r,temp_b1_6_27_i,temp_b1_8_25_r,temp_b1_8_25_i,temp_b1_8_27_r,temp_b1_8_27_i,temp_m2_6_25_r,temp_m2_6_25_i,temp_m2_6_27_r,temp_m2_6_27_i,temp_m2_8_25_r,temp_m2_8_25_i,temp_m2_8_27_r,temp_m2_8_27_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly315 (clk,temp_m2_6_25_r,temp_m2_6_25_i,temp_m2_6_27_r,temp_m2_6_27_i,temp_m2_8_25_r,temp_m2_8_25_i,temp_m2_8_27_r,temp_m2_8_27_i,temp_b2_6_25_r,temp_b2_6_25_i,temp_b2_6_27_r,temp_b2_6_27_i,temp_b2_8_25_r,temp_b2_8_25_i,temp_b2_8_27_r,temp_b2_8_27_i);
MULT MULT316 (clk,temp_b1_6_26_r,temp_b1_6_26_i,temp_b1_6_28_r,temp_b1_6_28_i,temp_b1_8_26_r,temp_b1_8_26_i,temp_b1_8_28_r,temp_b1_8_28_i,temp_m2_6_26_r,temp_m2_6_26_i,temp_m2_6_28_r,temp_m2_6_28_i,temp_m2_8_26_r,temp_m2_8_26_i,temp_m2_8_28_r,temp_m2_8_28_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly316 (clk,temp_m2_6_26_r,temp_m2_6_26_i,temp_m2_6_28_r,temp_m2_6_28_i,temp_m2_8_26_r,temp_m2_8_26_i,temp_m2_8_28_r,temp_m2_8_28_i,temp_b2_6_26_r,temp_b2_6_26_i,temp_b2_6_28_r,temp_b2_6_28_i,temp_b2_8_26_r,temp_b2_8_26_i,temp_b2_8_28_r,temp_b2_8_28_i);
MULT MULT317 (clk,temp_b1_5_29_r,temp_b1_5_29_i,temp_b1_5_31_r,temp_b1_5_31_i,temp_b1_7_29_r,temp_b1_7_29_i,temp_b1_7_31_r,temp_b1_7_31_i,temp_m2_5_29_r,temp_m2_5_29_i,temp_m2_5_31_r,temp_m2_5_31_i,temp_m2_7_29_r,temp_m2_7_29_i,temp_m2_7_31_r,temp_m2_7_31_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly317 (clk,temp_m2_5_29_r,temp_m2_5_29_i,temp_m2_5_31_r,temp_m2_5_31_i,temp_m2_7_29_r,temp_m2_7_29_i,temp_m2_7_31_r,temp_m2_7_31_i,temp_b2_5_29_r,temp_b2_5_29_i,temp_b2_5_31_r,temp_b2_5_31_i,temp_b2_7_29_r,temp_b2_7_29_i,temp_b2_7_31_r,temp_b2_7_31_i);
MULT MULT318 (clk,temp_b1_5_30_r,temp_b1_5_30_i,temp_b1_5_32_r,temp_b1_5_32_i,temp_b1_7_30_r,temp_b1_7_30_i,temp_b1_7_32_r,temp_b1_7_32_i,temp_m2_5_30_r,temp_m2_5_30_i,temp_m2_5_32_r,temp_m2_5_32_i,temp_m2_7_30_r,temp_m2_7_30_i,temp_m2_7_32_r,temp_m2_7_32_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly318 (clk,temp_m2_5_30_r,temp_m2_5_30_i,temp_m2_5_32_r,temp_m2_5_32_i,temp_m2_7_30_r,temp_m2_7_30_i,temp_m2_7_32_r,temp_m2_7_32_i,temp_b2_5_30_r,temp_b2_5_30_i,temp_b2_5_32_r,temp_b2_5_32_i,temp_b2_7_30_r,temp_b2_7_30_i,temp_b2_7_32_r,temp_b2_7_32_i);
MULT MULT319 (clk,temp_b1_6_29_r,temp_b1_6_29_i,temp_b1_6_31_r,temp_b1_6_31_i,temp_b1_8_29_r,temp_b1_8_29_i,temp_b1_8_31_r,temp_b1_8_31_i,temp_m2_6_29_r,temp_m2_6_29_i,temp_m2_6_31_r,temp_m2_6_31_i,temp_m2_8_29_r,temp_m2_8_29_i,temp_m2_8_31_r,temp_m2_8_31_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly319 (clk,temp_m2_6_29_r,temp_m2_6_29_i,temp_m2_6_31_r,temp_m2_6_31_i,temp_m2_8_29_r,temp_m2_8_29_i,temp_m2_8_31_r,temp_m2_8_31_i,temp_b2_6_29_r,temp_b2_6_29_i,temp_b2_6_31_r,temp_b2_6_31_i,temp_b2_8_29_r,temp_b2_8_29_i,temp_b2_8_31_r,temp_b2_8_31_i);
MULT MULT320 (clk,temp_b1_6_30_r,temp_b1_6_30_i,temp_b1_6_32_r,temp_b1_6_32_i,temp_b1_8_30_r,temp_b1_8_30_i,temp_b1_8_32_r,temp_b1_8_32_i,temp_m2_6_30_r,temp_m2_6_30_i,temp_m2_6_32_r,temp_m2_6_32_i,temp_m2_8_30_r,temp_m2_8_30_i,temp_m2_8_32_r,temp_m2_8_32_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly320 (clk,temp_m2_6_30_r,temp_m2_6_30_i,temp_m2_6_32_r,temp_m2_6_32_i,temp_m2_8_30_r,temp_m2_8_30_i,temp_m2_8_32_r,temp_m2_8_32_i,temp_b2_6_30_r,temp_b2_6_30_i,temp_b2_6_32_r,temp_b2_6_32_i,temp_b2_8_30_r,temp_b2_8_30_i,temp_b2_8_32_r,temp_b2_8_32_i);
MULT MULT321 (clk,temp_b1_9_1_r,temp_b1_9_1_i,temp_b1_9_3_r,temp_b1_9_3_i,temp_b1_11_1_r,temp_b1_11_1_i,temp_b1_11_3_r,temp_b1_11_3_i,temp_m2_9_1_r,temp_m2_9_1_i,temp_m2_9_3_r,temp_m2_9_3_i,temp_m2_11_1_r,temp_m2_11_1_i,temp_m2_11_3_r,temp_m2_11_3_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly321 (clk,temp_m2_9_1_r,temp_m2_9_1_i,temp_m2_9_3_r,temp_m2_9_3_i,temp_m2_11_1_r,temp_m2_11_1_i,temp_m2_11_3_r,temp_m2_11_3_i,temp_b2_9_1_r,temp_b2_9_1_i,temp_b2_9_3_r,temp_b2_9_3_i,temp_b2_11_1_r,temp_b2_11_1_i,temp_b2_11_3_r,temp_b2_11_3_i);
MULT MULT322 (clk,temp_b1_9_2_r,temp_b1_9_2_i,temp_b1_9_4_r,temp_b1_9_4_i,temp_b1_11_2_r,temp_b1_11_2_i,temp_b1_11_4_r,temp_b1_11_4_i,temp_m2_9_2_r,temp_m2_9_2_i,temp_m2_9_4_r,temp_m2_9_4_i,temp_m2_11_2_r,temp_m2_11_2_i,temp_m2_11_4_r,temp_m2_11_4_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly322 (clk,temp_m2_9_2_r,temp_m2_9_2_i,temp_m2_9_4_r,temp_m2_9_4_i,temp_m2_11_2_r,temp_m2_11_2_i,temp_m2_11_4_r,temp_m2_11_4_i,temp_b2_9_2_r,temp_b2_9_2_i,temp_b2_9_4_r,temp_b2_9_4_i,temp_b2_11_2_r,temp_b2_11_2_i,temp_b2_11_4_r,temp_b2_11_4_i);
MULT MULT323 (clk,temp_b1_10_1_r,temp_b1_10_1_i,temp_b1_10_3_r,temp_b1_10_3_i,temp_b1_12_1_r,temp_b1_12_1_i,temp_b1_12_3_r,temp_b1_12_3_i,temp_m2_10_1_r,temp_m2_10_1_i,temp_m2_10_3_r,temp_m2_10_3_i,temp_m2_12_1_r,temp_m2_12_1_i,temp_m2_12_3_r,temp_m2_12_3_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly323 (clk,temp_m2_10_1_r,temp_m2_10_1_i,temp_m2_10_3_r,temp_m2_10_3_i,temp_m2_12_1_r,temp_m2_12_1_i,temp_m2_12_3_r,temp_m2_12_3_i,temp_b2_10_1_r,temp_b2_10_1_i,temp_b2_10_3_r,temp_b2_10_3_i,temp_b2_12_1_r,temp_b2_12_1_i,temp_b2_12_3_r,temp_b2_12_3_i);
MULT MULT324 (clk,temp_b1_10_2_r,temp_b1_10_2_i,temp_b1_10_4_r,temp_b1_10_4_i,temp_b1_12_2_r,temp_b1_12_2_i,temp_b1_12_4_r,temp_b1_12_4_i,temp_m2_10_2_r,temp_m2_10_2_i,temp_m2_10_4_r,temp_m2_10_4_i,temp_m2_12_2_r,temp_m2_12_2_i,temp_m2_12_4_r,temp_m2_12_4_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly324 (clk,temp_m2_10_2_r,temp_m2_10_2_i,temp_m2_10_4_r,temp_m2_10_4_i,temp_m2_12_2_r,temp_m2_12_2_i,temp_m2_12_4_r,temp_m2_12_4_i,temp_b2_10_2_r,temp_b2_10_2_i,temp_b2_10_4_r,temp_b2_10_4_i,temp_b2_12_2_r,temp_b2_12_2_i,temp_b2_12_4_r,temp_b2_12_4_i);
MULT MULT325 (clk,temp_b1_9_5_r,temp_b1_9_5_i,temp_b1_9_7_r,temp_b1_9_7_i,temp_b1_11_5_r,temp_b1_11_5_i,temp_b1_11_7_r,temp_b1_11_7_i,temp_m2_9_5_r,temp_m2_9_5_i,temp_m2_9_7_r,temp_m2_9_7_i,temp_m2_11_5_r,temp_m2_11_5_i,temp_m2_11_7_r,temp_m2_11_7_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly325 (clk,temp_m2_9_5_r,temp_m2_9_5_i,temp_m2_9_7_r,temp_m2_9_7_i,temp_m2_11_5_r,temp_m2_11_5_i,temp_m2_11_7_r,temp_m2_11_7_i,temp_b2_9_5_r,temp_b2_9_5_i,temp_b2_9_7_r,temp_b2_9_7_i,temp_b2_11_5_r,temp_b2_11_5_i,temp_b2_11_7_r,temp_b2_11_7_i);
MULT MULT326 (clk,temp_b1_9_6_r,temp_b1_9_6_i,temp_b1_9_8_r,temp_b1_9_8_i,temp_b1_11_6_r,temp_b1_11_6_i,temp_b1_11_8_r,temp_b1_11_8_i,temp_m2_9_6_r,temp_m2_9_6_i,temp_m2_9_8_r,temp_m2_9_8_i,temp_m2_11_6_r,temp_m2_11_6_i,temp_m2_11_8_r,temp_m2_11_8_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly326 (clk,temp_m2_9_6_r,temp_m2_9_6_i,temp_m2_9_8_r,temp_m2_9_8_i,temp_m2_11_6_r,temp_m2_11_6_i,temp_m2_11_8_r,temp_m2_11_8_i,temp_b2_9_6_r,temp_b2_9_6_i,temp_b2_9_8_r,temp_b2_9_8_i,temp_b2_11_6_r,temp_b2_11_6_i,temp_b2_11_8_r,temp_b2_11_8_i);
MULT MULT327 (clk,temp_b1_10_5_r,temp_b1_10_5_i,temp_b1_10_7_r,temp_b1_10_7_i,temp_b1_12_5_r,temp_b1_12_5_i,temp_b1_12_7_r,temp_b1_12_7_i,temp_m2_10_5_r,temp_m2_10_5_i,temp_m2_10_7_r,temp_m2_10_7_i,temp_m2_12_5_r,temp_m2_12_5_i,temp_m2_12_7_r,temp_m2_12_7_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly327 (clk,temp_m2_10_5_r,temp_m2_10_5_i,temp_m2_10_7_r,temp_m2_10_7_i,temp_m2_12_5_r,temp_m2_12_5_i,temp_m2_12_7_r,temp_m2_12_7_i,temp_b2_10_5_r,temp_b2_10_5_i,temp_b2_10_7_r,temp_b2_10_7_i,temp_b2_12_5_r,temp_b2_12_5_i,temp_b2_12_7_r,temp_b2_12_7_i);
MULT MULT328 (clk,temp_b1_10_6_r,temp_b1_10_6_i,temp_b1_10_8_r,temp_b1_10_8_i,temp_b1_12_6_r,temp_b1_12_6_i,temp_b1_12_8_r,temp_b1_12_8_i,temp_m2_10_6_r,temp_m2_10_6_i,temp_m2_10_8_r,temp_m2_10_8_i,temp_m2_12_6_r,temp_m2_12_6_i,temp_m2_12_8_r,temp_m2_12_8_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly328 (clk,temp_m2_10_6_r,temp_m2_10_6_i,temp_m2_10_8_r,temp_m2_10_8_i,temp_m2_12_6_r,temp_m2_12_6_i,temp_m2_12_8_r,temp_m2_12_8_i,temp_b2_10_6_r,temp_b2_10_6_i,temp_b2_10_8_r,temp_b2_10_8_i,temp_b2_12_6_r,temp_b2_12_6_i,temp_b2_12_8_r,temp_b2_12_8_i);
MULT MULT329 (clk,temp_b1_9_9_r,temp_b1_9_9_i,temp_b1_9_11_r,temp_b1_9_11_i,temp_b1_11_9_r,temp_b1_11_9_i,temp_b1_11_11_r,temp_b1_11_11_i,temp_m2_9_9_r,temp_m2_9_9_i,temp_m2_9_11_r,temp_m2_9_11_i,temp_m2_11_9_r,temp_m2_11_9_i,temp_m2_11_11_r,temp_m2_11_11_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly329 (clk,temp_m2_9_9_r,temp_m2_9_9_i,temp_m2_9_11_r,temp_m2_9_11_i,temp_m2_11_9_r,temp_m2_11_9_i,temp_m2_11_11_r,temp_m2_11_11_i,temp_b2_9_9_r,temp_b2_9_9_i,temp_b2_9_11_r,temp_b2_9_11_i,temp_b2_11_9_r,temp_b2_11_9_i,temp_b2_11_11_r,temp_b2_11_11_i);
MULT MULT330 (clk,temp_b1_9_10_r,temp_b1_9_10_i,temp_b1_9_12_r,temp_b1_9_12_i,temp_b1_11_10_r,temp_b1_11_10_i,temp_b1_11_12_r,temp_b1_11_12_i,temp_m2_9_10_r,temp_m2_9_10_i,temp_m2_9_12_r,temp_m2_9_12_i,temp_m2_11_10_r,temp_m2_11_10_i,temp_m2_11_12_r,temp_m2_11_12_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly330 (clk,temp_m2_9_10_r,temp_m2_9_10_i,temp_m2_9_12_r,temp_m2_9_12_i,temp_m2_11_10_r,temp_m2_11_10_i,temp_m2_11_12_r,temp_m2_11_12_i,temp_b2_9_10_r,temp_b2_9_10_i,temp_b2_9_12_r,temp_b2_9_12_i,temp_b2_11_10_r,temp_b2_11_10_i,temp_b2_11_12_r,temp_b2_11_12_i);
MULT MULT331 (clk,temp_b1_10_9_r,temp_b1_10_9_i,temp_b1_10_11_r,temp_b1_10_11_i,temp_b1_12_9_r,temp_b1_12_9_i,temp_b1_12_11_r,temp_b1_12_11_i,temp_m2_10_9_r,temp_m2_10_9_i,temp_m2_10_11_r,temp_m2_10_11_i,temp_m2_12_9_r,temp_m2_12_9_i,temp_m2_12_11_r,temp_m2_12_11_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly331 (clk,temp_m2_10_9_r,temp_m2_10_9_i,temp_m2_10_11_r,temp_m2_10_11_i,temp_m2_12_9_r,temp_m2_12_9_i,temp_m2_12_11_r,temp_m2_12_11_i,temp_b2_10_9_r,temp_b2_10_9_i,temp_b2_10_11_r,temp_b2_10_11_i,temp_b2_12_9_r,temp_b2_12_9_i,temp_b2_12_11_r,temp_b2_12_11_i);
MULT MULT332 (clk,temp_b1_10_10_r,temp_b1_10_10_i,temp_b1_10_12_r,temp_b1_10_12_i,temp_b1_12_10_r,temp_b1_12_10_i,temp_b1_12_12_r,temp_b1_12_12_i,temp_m2_10_10_r,temp_m2_10_10_i,temp_m2_10_12_r,temp_m2_10_12_i,temp_m2_12_10_r,temp_m2_12_10_i,temp_m2_12_12_r,temp_m2_12_12_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly332 (clk,temp_m2_10_10_r,temp_m2_10_10_i,temp_m2_10_12_r,temp_m2_10_12_i,temp_m2_12_10_r,temp_m2_12_10_i,temp_m2_12_12_r,temp_m2_12_12_i,temp_b2_10_10_r,temp_b2_10_10_i,temp_b2_10_12_r,temp_b2_10_12_i,temp_b2_12_10_r,temp_b2_12_10_i,temp_b2_12_12_r,temp_b2_12_12_i);
MULT MULT333 (clk,temp_b1_9_13_r,temp_b1_9_13_i,temp_b1_9_15_r,temp_b1_9_15_i,temp_b1_11_13_r,temp_b1_11_13_i,temp_b1_11_15_r,temp_b1_11_15_i,temp_m2_9_13_r,temp_m2_9_13_i,temp_m2_9_15_r,temp_m2_9_15_i,temp_m2_11_13_r,temp_m2_11_13_i,temp_m2_11_15_r,temp_m2_11_15_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly333 (clk,temp_m2_9_13_r,temp_m2_9_13_i,temp_m2_9_15_r,temp_m2_9_15_i,temp_m2_11_13_r,temp_m2_11_13_i,temp_m2_11_15_r,temp_m2_11_15_i,temp_b2_9_13_r,temp_b2_9_13_i,temp_b2_9_15_r,temp_b2_9_15_i,temp_b2_11_13_r,temp_b2_11_13_i,temp_b2_11_15_r,temp_b2_11_15_i);
MULT MULT334 (clk,temp_b1_9_14_r,temp_b1_9_14_i,temp_b1_9_16_r,temp_b1_9_16_i,temp_b1_11_14_r,temp_b1_11_14_i,temp_b1_11_16_r,temp_b1_11_16_i,temp_m2_9_14_r,temp_m2_9_14_i,temp_m2_9_16_r,temp_m2_9_16_i,temp_m2_11_14_r,temp_m2_11_14_i,temp_m2_11_16_r,temp_m2_11_16_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly334 (clk,temp_m2_9_14_r,temp_m2_9_14_i,temp_m2_9_16_r,temp_m2_9_16_i,temp_m2_11_14_r,temp_m2_11_14_i,temp_m2_11_16_r,temp_m2_11_16_i,temp_b2_9_14_r,temp_b2_9_14_i,temp_b2_9_16_r,temp_b2_9_16_i,temp_b2_11_14_r,temp_b2_11_14_i,temp_b2_11_16_r,temp_b2_11_16_i);
MULT MULT335 (clk,temp_b1_10_13_r,temp_b1_10_13_i,temp_b1_10_15_r,temp_b1_10_15_i,temp_b1_12_13_r,temp_b1_12_13_i,temp_b1_12_15_r,temp_b1_12_15_i,temp_m2_10_13_r,temp_m2_10_13_i,temp_m2_10_15_r,temp_m2_10_15_i,temp_m2_12_13_r,temp_m2_12_13_i,temp_m2_12_15_r,temp_m2_12_15_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly335 (clk,temp_m2_10_13_r,temp_m2_10_13_i,temp_m2_10_15_r,temp_m2_10_15_i,temp_m2_12_13_r,temp_m2_12_13_i,temp_m2_12_15_r,temp_m2_12_15_i,temp_b2_10_13_r,temp_b2_10_13_i,temp_b2_10_15_r,temp_b2_10_15_i,temp_b2_12_13_r,temp_b2_12_13_i,temp_b2_12_15_r,temp_b2_12_15_i);
MULT MULT336 (clk,temp_b1_10_14_r,temp_b1_10_14_i,temp_b1_10_16_r,temp_b1_10_16_i,temp_b1_12_14_r,temp_b1_12_14_i,temp_b1_12_16_r,temp_b1_12_16_i,temp_m2_10_14_r,temp_m2_10_14_i,temp_m2_10_16_r,temp_m2_10_16_i,temp_m2_12_14_r,temp_m2_12_14_i,temp_m2_12_16_r,temp_m2_12_16_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly336 (clk,temp_m2_10_14_r,temp_m2_10_14_i,temp_m2_10_16_r,temp_m2_10_16_i,temp_m2_12_14_r,temp_m2_12_14_i,temp_m2_12_16_r,temp_m2_12_16_i,temp_b2_10_14_r,temp_b2_10_14_i,temp_b2_10_16_r,temp_b2_10_16_i,temp_b2_12_14_r,temp_b2_12_14_i,temp_b2_12_16_r,temp_b2_12_16_i);
MULT MULT337 (clk,temp_b1_9_17_r,temp_b1_9_17_i,temp_b1_9_19_r,temp_b1_9_19_i,temp_b1_11_17_r,temp_b1_11_17_i,temp_b1_11_19_r,temp_b1_11_19_i,temp_m2_9_17_r,temp_m2_9_17_i,temp_m2_9_19_r,temp_m2_9_19_i,temp_m2_11_17_r,temp_m2_11_17_i,temp_m2_11_19_r,temp_m2_11_19_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly337 (clk,temp_m2_9_17_r,temp_m2_9_17_i,temp_m2_9_19_r,temp_m2_9_19_i,temp_m2_11_17_r,temp_m2_11_17_i,temp_m2_11_19_r,temp_m2_11_19_i,temp_b2_9_17_r,temp_b2_9_17_i,temp_b2_9_19_r,temp_b2_9_19_i,temp_b2_11_17_r,temp_b2_11_17_i,temp_b2_11_19_r,temp_b2_11_19_i);
MULT MULT338 (clk,temp_b1_9_18_r,temp_b1_9_18_i,temp_b1_9_20_r,temp_b1_9_20_i,temp_b1_11_18_r,temp_b1_11_18_i,temp_b1_11_20_r,temp_b1_11_20_i,temp_m2_9_18_r,temp_m2_9_18_i,temp_m2_9_20_r,temp_m2_9_20_i,temp_m2_11_18_r,temp_m2_11_18_i,temp_m2_11_20_r,temp_m2_11_20_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly338 (clk,temp_m2_9_18_r,temp_m2_9_18_i,temp_m2_9_20_r,temp_m2_9_20_i,temp_m2_11_18_r,temp_m2_11_18_i,temp_m2_11_20_r,temp_m2_11_20_i,temp_b2_9_18_r,temp_b2_9_18_i,temp_b2_9_20_r,temp_b2_9_20_i,temp_b2_11_18_r,temp_b2_11_18_i,temp_b2_11_20_r,temp_b2_11_20_i);
MULT MULT339 (clk,temp_b1_10_17_r,temp_b1_10_17_i,temp_b1_10_19_r,temp_b1_10_19_i,temp_b1_12_17_r,temp_b1_12_17_i,temp_b1_12_19_r,temp_b1_12_19_i,temp_m2_10_17_r,temp_m2_10_17_i,temp_m2_10_19_r,temp_m2_10_19_i,temp_m2_12_17_r,temp_m2_12_17_i,temp_m2_12_19_r,temp_m2_12_19_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly339 (clk,temp_m2_10_17_r,temp_m2_10_17_i,temp_m2_10_19_r,temp_m2_10_19_i,temp_m2_12_17_r,temp_m2_12_17_i,temp_m2_12_19_r,temp_m2_12_19_i,temp_b2_10_17_r,temp_b2_10_17_i,temp_b2_10_19_r,temp_b2_10_19_i,temp_b2_12_17_r,temp_b2_12_17_i,temp_b2_12_19_r,temp_b2_12_19_i);
MULT MULT340 (clk,temp_b1_10_18_r,temp_b1_10_18_i,temp_b1_10_20_r,temp_b1_10_20_i,temp_b1_12_18_r,temp_b1_12_18_i,temp_b1_12_20_r,temp_b1_12_20_i,temp_m2_10_18_r,temp_m2_10_18_i,temp_m2_10_20_r,temp_m2_10_20_i,temp_m2_12_18_r,temp_m2_12_18_i,temp_m2_12_20_r,temp_m2_12_20_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly340 (clk,temp_m2_10_18_r,temp_m2_10_18_i,temp_m2_10_20_r,temp_m2_10_20_i,temp_m2_12_18_r,temp_m2_12_18_i,temp_m2_12_20_r,temp_m2_12_20_i,temp_b2_10_18_r,temp_b2_10_18_i,temp_b2_10_20_r,temp_b2_10_20_i,temp_b2_12_18_r,temp_b2_12_18_i,temp_b2_12_20_r,temp_b2_12_20_i);
MULT MULT341 (clk,temp_b1_9_21_r,temp_b1_9_21_i,temp_b1_9_23_r,temp_b1_9_23_i,temp_b1_11_21_r,temp_b1_11_21_i,temp_b1_11_23_r,temp_b1_11_23_i,temp_m2_9_21_r,temp_m2_9_21_i,temp_m2_9_23_r,temp_m2_9_23_i,temp_m2_11_21_r,temp_m2_11_21_i,temp_m2_11_23_r,temp_m2_11_23_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly341 (clk,temp_m2_9_21_r,temp_m2_9_21_i,temp_m2_9_23_r,temp_m2_9_23_i,temp_m2_11_21_r,temp_m2_11_21_i,temp_m2_11_23_r,temp_m2_11_23_i,temp_b2_9_21_r,temp_b2_9_21_i,temp_b2_9_23_r,temp_b2_9_23_i,temp_b2_11_21_r,temp_b2_11_21_i,temp_b2_11_23_r,temp_b2_11_23_i);
MULT MULT342 (clk,temp_b1_9_22_r,temp_b1_9_22_i,temp_b1_9_24_r,temp_b1_9_24_i,temp_b1_11_22_r,temp_b1_11_22_i,temp_b1_11_24_r,temp_b1_11_24_i,temp_m2_9_22_r,temp_m2_9_22_i,temp_m2_9_24_r,temp_m2_9_24_i,temp_m2_11_22_r,temp_m2_11_22_i,temp_m2_11_24_r,temp_m2_11_24_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly342 (clk,temp_m2_9_22_r,temp_m2_9_22_i,temp_m2_9_24_r,temp_m2_9_24_i,temp_m2_11_22_r,temp_m2_11_22_i,temp_m2_11_24_r,temp_m2_11_24_i,temp_b2_9_22_r,temp_b2_9_22_i,temp_b2_9_24_r,temp_b2_9_24_i,temp_b2_11_22_r,temp_b2_11_22_i,temp_b2_11_24_r,temp_b2_11_24_i);
MULT MULT343 (clk,temp_b1_10_21_r,temp_b1_10_21_i,temp_b1_10_23_r,temp_b1_10_23_i,temp_b1_12_21_r,temp_b1_12_21_i,temp_b1_12_23_r,temp_b1_12_23_i,temp_m2_10_21_r,temp_m2_10_21_i,temp_m2_10_23_r,temp_m2_10_23_i,temp_m2_12_21_r,temp_m2_12_21_i,temp_m2_12_23_r,temp_m2_12_23_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly343 (clk,temp_m2_10_21_r,temp_m2_10_21_i,temp_m2_10_23_r,temp_m2_10_23_i,temp_m2_12_21_r,temp_m2_12_21_i,temp_m2_12_23_r,temp_m2_12_23_i,temp_b2_10_21_r,temp_b2_10_21_i,temp_b2_10_23_r,temp_b2_10_23_i,temp_b2_12_21_r,temp_b2_12_21_i,temp_b2_12_23_r,temp_b2_12_23_i);
MULT MULT344 (clk,temp_b1_10_22_r,temp_b1_10_22_i,temp_b1_10_24_r,temp_b1_10_24_i,temp_b1_12_22_r,temp_b1_12_22_i,temp_b1_12_24_r,temp_b1_12_24_i,temp_m2_10_22_r,temp_m2_10_22_i,temp_m2_10_24_r,temp_m2_10_24_i,temp_m2_12_22_r,temp_m2_12_22_i,temp_m2_12_24_r,temp_m2_12_24_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly344 (clk,temp_m2_10_22_r,temp_m2_10_22_i,temp_m2_10_24_r,temp_m2_10_24_i,temp_m2_12_22_r,temp_m2_12_22_i,temp_m2_12_24_r,temp_m2_12_24_i,temp_b2_10_22_r,temp_b2_10_22_i,temp_b2_10_24_r,temp_b2_10_24_i,temp_b2_12_22_r,temp_b2_12_22_i,temp_b2_12_24_r,temp_b2_12_24_i);
MULT MULT345 (clk,temp_b1_9_25_r,temp_b1_9_25_i,temp_b1_9_27_r,temp_b1_9_27_i,temp_b1_11_25_r,temp_b1_11_25_i,temp_b1_11_27_r,temp_b1_11_27_i,temp_m2_9_25_r,temp_m2_9_25_i,temp_m2_9_27_r,temp_m2_9_27_i,temp_m2_11_25_r,temp_m2_11_25_i,temp_m2_11_27_r,temp_m2_11_27_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly345 (clk,temp_m2_9_25_r,temp_m2_9_25_i,temp_m2_9_27_r,temp_m2_9_27_i,temp_m2_11_25_r,temp_m2_11_25_i,temp_m2_11_27_r,temp_m2_11_27_i,temp_b2_9_25_r,temp_b2_9_25_i,temp_b2_9_27_r,temp_b2_9_27_i,temp_b2_11_25_r,temp_b2_11_25_i,temp_b2_11_27_r,temp_b2_11_27_i);
MULT MULT346 (clk,temp_b1_9_26_r,temp_b1_9_26_i,temp_b1_9_28_r,temp_b1_9_28_i,temp_b1_11_26_r,temp_b1_11_26_i,temp_b1_11_28_r,temp_b1_11_28_i,temp_m2_9_26_r,temp_m2_9_26_i,temp_m2_9_28_r,temp_m2_9_28_i,temp_m2_11_26_r,temp_m2_11_26_i,temp_m2_11_28_r,temp_m2_11_28_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly346 (clk,temp_m2_9_26_r,temp_m2_9_26_i,temp_m2_9_28_r,temp_m2_9_28_i,temp_m2_11_26_r,temp_m2_11_26_i,temp_m2_11_28_r,temp_m2_11_28_i,temp_b2_9_26_r,temp_b2_9_26_i,temp_b2_9_28_r,temp_b2_9_28_i,temp_b2_11_26_r,temp_b2_11_26_i,temp_b2_11_28_r,temp_b2_11_28_i);
MULT MULT347 (clk,temp_b1_10_25_r,temp_b1_10_25_i,temp_b1_10_27_r,temp_b1_10_27_i,temp_b1_12_25_r,temp_b1_12_25_i,temp_b1_12_27_r,temp_b1_12_27_i,temp_m2_10_25_r,temp_m2_10_25_i,temp_m2_10_27_r,temp_m2_10_27_i,temp_m2_12_25_r,temp_m2_12_25_i,temp_m2_12_27_r,temp_m2_12_27_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly347 (clk,temp_m2_10_25_r,temp_m2_10_25_i,temp_m2_10_27_r,temp_m2_10_27_i,temp_m2_12_25_r,temp_m2_12_25_i,temp_m2_12_27_r,temp_m2_12_27_i,temp_b2_10_25_r,temp_b2_10_25_i,temp_b2_10_27_r,temp_b2_10_27_i,temp_b2_12_25_r,temp_b2_12_25_i,temp_b2_12_27_r,temp_b2_12_27_i);
MULT MULT348 (clk,temp_b1_10_26_r,temp_b1_10_26_i,temp_b1_10_28_r,temp_b1_10_28_i,temp_b1_12_26_r,temp_b1_12_26_i,temp_b1_12_28_r,temp_b1_12_28_i,temp_m2_10_26_r,temp_m2_10_26_i,temp_m2_10_28_r,temp_m2_10_28_i,temp_m2_12_26_r,temp_m2_12_26_i,temp_m2_12_28_r,temp_m2_12_28_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly348 (clk,temp_m2_10_26_r,temp_m2_10_26_i,temp_m2_10_28_r,temp_m2_10_28_i,temp_m2_12_26_r,temp_m2_12_26_i,temp_m2_12_28_r,temp_m2_12_28_i,temp_b2_10_26_r,temp_b2_10_26_i,temp_b2_10_28_r,temp_b2_10_28_i,temp_b2_12_26_r,temp_b2_12_26_i,temp_b2_12_28_r,temp_b2_12_28_i);
MULT MULT349 (clk,temp_b1_9_29_r,temp_b1_9_29_i,temp_b1_9_31_r,temp_b1_9_31_i,temp_b1_11_29_r,temp_b1_11_29_i,temp_b1_11_31_r,temp_b1_11_31_i,temp_m2_9_29_r,temp_m2_9_29_i,temp_m2_9_31_r,temp_m2_9_31_i,temp_m2_11_29_r,temp_m2_11_29_i,temp_m2_11_31_r,temp_m2_11_31_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly349 (clk,temp_m2_9_29_r,temp_m2_9_29_i,temp_m2_9_31_r,temp_m2_9_31_i,temp_m2_11_29_r,temp_m2_11_29_i,temp_m2_11_31_r,temp_m2_11_31_i,temp_b2_9_29_r,temp_b2_9_29_i,temp_b2_9_31_r,temp_b2_9_31_i,temp_b2_11_29_r,temp_b2_11_29_i,temp_b2_11_31_r,temp_b2_11_31_i);
MULT MULT350 (clk,temp_b1_9_30_r,temp_b1_9_30_i,temp_b1_9_32_r,temp_b1_9_32_i,temp_b1_11_30_r,temp_b1_11_30_i,temp_b1_11_32_r,temp_b1_11_32_i,temp_m2_9_30_r,temp_m2_9_30_i,temp_m2_9_32_r,temp_m2_9_32_i,temp_m2_11_30_r,temp_m2_11_30_i,temp_m2_11_32_r,temp_m2_11_32_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly350 (clk,temp_m2_9_30_r,temp_m2_9_30_i,temp_m2_9_32_r,temp_m2_9_32_i,temp_m2_11_30_r,temp_m2_11_30_i,temp_m2_11_32_r,temp_m2_11_32_i,temp_b2_9_30_r,temp_b2_9_30_i,temp_b2_9_32_r,temp_b2_9_32_i,temp_b2_11_30_r,temp_b2_11_30_i,temp_b2_11_32_r,temp_b2_11_32_i);
MULT MULT351 (clk,temp_b1_10_29_r,temp_b1_10_29_i,temp_b1_10_31_r,temp_b1_10_31_i,temp_b1_12_29_r,temp_b1_12_29_i,temp_b1_12_31_r,temp_b1_12_31_i,temp_m2_10_29_r,temp_m2_10_29_i,temp_m2_10_31_r,temp_m2_10_31_i,temp_m2_12_29_r,temp_m2_12_29_i,temp_m2_12_31_r,temp_m2_12_31_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly351 (clk,temp_m2_10_29_r,temp_m2_10_29_i,temp_m2_10_31_r,temp_m2_10_31_i,temp_m2_12_29_r,temp_m2_12_29_i,temp_m2_12_31_r,temp_m2_12_31_i,temp_b2_10_29_r,temp_b2_10_29_i,temp_b2_10_31_r,temp_b2_10_31_i,temp_b2_12_29_r,temp_b2_12_29_i,temp_b2_12_31_r,temp_b2_12_31_i);
MULT MULT352 (clk,temp_b1_10_30_r,temp_b1_10_30_i,temp_b1_10_32_r,temp_b1_10_32_i,temp_b1_12_30_r,temp_b1_12_30_i,temp_b1_12_32_r,temp_b1_12_32_i,temp_m2_10_30_r,temp_m2_10_30_i,temp_m2_10_32_r,temp_m2_10_32_i,temp_m2_12_30_r,temp_m2_12_30_i,temp_m2_12_32_r,temp_m2_12_32_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly352 (clk,temp_m2_10_30_r,temp_m2_10_30_i,temp_m2_10_32_r,temp_m2_10_32_i,temp_m2_12_30_r,temp_m2_12_30_i,temp_m2_12_32_r,temp_m2_12_32_i,temp_b2_10_30_r,temp_b2_10_30_i,temp_b2_10_32_r,temp_b2_10_32_i,temp_b2_12_30_r,temp_b2_12_30_i,temp_b2_12_32_r,temp_b2_12_32_i);
MULT MULT353 (clk,temp_b1_13_1_r,temp_b1_13_1_i,temp_b1_13_3_r,temp_b1_13_3_i,temp_b1_15_1_r,temp_b1_15_1_i,temp_b1_15_3_r,temp_b1_15_3_i,temp_m2_13_1_r,temp_m2_13_1_i,temp_m2_13_3_r,temp_m2_13_3_i,temp_m2_15_1_r,temp_m2_15_1_i,temp_m2_15_3_r,temp_m2_15_3_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly353 (clk,temp_m2_13_1_r,temp_m2_13_1_i,temp_m2_13_3_r,temp_m2_13_3_i,temp_m2_15_1_r,temp_m2_15_1_i,temp_m2_15_3_r,temp_m2_15_3_i,temp_b2_13_1_r,temp_b2_13_1_i,temp_b2_13_3_r,temp_b2_13_3_i,temp_b2_15_1_r,temp_b2_15_1_i,temp_b2_15_3_r,temp_b2_15_3_i);
MULT MULT354 (clk,temp_b1_13_2_r,temp_b1_13_2_i,temp_b1_13_4_r,temp_b1_13_4_i,temp_b1_15_2_r,temp_b1_15_2_i,temp_b1_15_4_r,temp_b1_15_4_i,temp_m2_13_2_r,temp_m2_13_2_i,temp_m2_13_4_r,temp_m2_13_4_i,temp_m2_15_2_r,temp_m2_15_2_i,temp_m2_15_4_r,temp_m2_15_4_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly354 (clk,temp_m2_13_2_r,temp_m2_13_2_i,temp_m2_13_4_r,temp_m2_13_4_i,temp_m2_15_2_r,temp_m2_15_2_i,temp_m2_15_4_r,temp_m2_15_4_i,temp_b2_13_2_r,temp_b2_13_2_i,temp_b2_13_4_r,temp_b2_13_4_i,temp_b2_15_2_r,temp_b2_15_2_i,temp_b2_15_4_r,temp_b2_15_4_i);
MULT MULT355 (clk,temp_b1_14_1_r,temp_b1_14_1_i,temp_b1_14_3_r,temp_b1_14_3_i,temp_b1_16_1_r,temp_b1_16_1_i,temp_b1_16_3_r,temp_b1_16_3_i,temp_m2_14_1_r,temp_m2_14_1_i,temp_m2_14_3_r,temp_m2_14_3_i,temp_m2_16_1_r,temp_m2_16_1_i,temp_m2_16_3_r,temp_m2_16_3_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly355 (clk,temp_m2_14_1_r,temp_m2_14_1_i,temp_m2_14_3_r,temp_m2_14_3_i,temp_m2_16_1_r,temp_m2_16_1_i,temp_m2_16_3_r,temp_m2_16_3_i,temp_b2_14_1_r,temp_b2_14_1_i,temp_b2_14_3_r,temp_b2_14_3_i,temp_b2_16_1_r,temp_b2_16_1_i,temp_b2_16_3_r,temp_b2_16_3_i);
MULT MULT356 (clk,temp_b1_14_2_r,temp_b1_14_2_i,temp_b1_14_4_r,temp_b1_14_4_i,temp_b1_16_2_r,temp_b1_16_2_i,temp_b1_16_4_r,temp_b1_16_4_i,temp_m2_14_2_r,temp_m2_14_2_i,temp_m2_14_4_r,temp_m2_14_4_i,temp_m2_16_2_r,temp_m2_16_2_i,temp_m2_16_4_r,temp_m2_16_4_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly356 (clk,temp_m2_14_2_r,temp_m2_14_2_i,temp_m2_14_4_r,temp_m2_14_4_i,temp_m2_16_2_r,temp_m2_16_2_i,temp_m2_16_4_r,temp_m2_16_4_i,temp_b2_14_2_r,temp_b2_14_2_i,temp_b2_14_4_r,temp_b2_14_4_i,temp_b2_16_2_r,temp_b2_16_2_i,temp_b2_16_4_r,temp_b2_16_4_i);
MULT MULT357 (clk,temp_b1_13_5_r,temp_b1_13_5_i,temp_b1_13_7_r,temp_b1_13_7_i,temp_b1_15_5_r,temp_b1_15_5_i,temp_b1_15_7_r,temp_b1_15_7_i,temp_m2_13_5_r,temp_m2_13_5_i,temp_m2_13_7_r,temp_m2_13_7_i,temp_m2_15_5_r,temp_m2_15_5_i,temp_m2_15_7_r,temp_m2_15_7_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly357 (clk,temp_m2_13_5_r,temp_m2_13_5_i,temp_m2_13_7_r,temp_m2_13_7_i,temp_m2_15_5_r,temp_m2_15_5_i,temp_m2_15_7_r,temp_m2_15_7_i,temp_b2_13_5_r,temp_b2_13_5_i,temp_b2_13_7_r,temp_b2_13_7_i,temp_b2_15_5_r,temp_b2_15_5_i,temp_b2_15_7_r,temp_b2_15_7_i);
MULT MULT358 (clk,temp_b1_13_6_r,temp_b1_13_6_i,temp_b1_13_8_r,temp_b1_13_8_i,temp_b1_15_6_r,temp_b1_15_6_i,temp_b1_15_8_r,temp_b1_15_8_i,temp_m2_13_6_r,temp_m2_13_6_i,temp_m2_13_8_r,temp_m2_13_8_i,temp_m2_15_6_r,temp_m2_15_6_i,temp_m2_15_8_r,temp_m2_15_8_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly358 (clk,temp_m2_13_6_r,temp_m2_13_6_i,temp_m2_13_8_r,temp_m2_13_8_i,temp_m2_15_6_r,temp_m2_15_6_i,temp_m2_15_8_r,temp_m2_15_8_i,temp_b2_13_6_r,temp_b2_13_6_i,temp_b2_13_8_r,temp_b2_13_8_i,temp_b2_15_6_r,temp_b2_15_6_i,temp_b2_15_8_r,temp_b2_15_8_i);
MULT MULT359 (clk,temp_b1_14_5_r,temp_b1_14_5_i,temp_b1_14_7_r,temp_b1_14_7_i,temp_b1_16_5_r,temp_b1_16_5_i,temp_b1_16_7_r,temp_b1_16_7_i,temp_m2_14_5_r,temp_m2_14_5_i,temp_m2_14_7_r,temp_m2_14_7_i,temp_m2_16_5_r,temp_m2_16_5_i,temp_m2_16_7_r,temp_m2_16_7_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly359 (clk,temp_m2_14_5_r,temp_m2_14_5_i,temp_m2_14_7_r,temp_m2_14_7_i,temp_m2_16_5_r,temp_m2_16_5_i,temp_m2_16_7_r,temp_m2_16_7_i,temp_b2_14_5_r,temp_b2_14_5_i,temp_b2_14_7_r,temp_b2_14_7_i,temp_b2_16_5_r,temp_b2_16_5_i,temp_b2_16_7_r,temp_b2_16_7_i);
MULT MULT360 (clk,temp_b1_14_6_r,temp_b1_14_6_i,temp_b1_14_8_r,temp_b1_14_8_i,temp_b1_16_6_r,temp_b1_16_6_i,temp_b1_16_8_r,temp_b1_16_8_i,temp_m2_14_6_r,temp_m2_14_6_i,temp_m2_14_8_r,temp_m2_14_8_i,temp_m2_16_6_r,temp_m2_16_6_i,temp_m2_16_8_r,temp_m2_16_8_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly360 (clk,temp_m2_14_6_r,temp_m2_14_6_i,temp_m2_14_8_r,temp_m2_14_8_i,temp_m2_16_6_r,temp_m2_16_6_i,temp_m2_16_8_r,temp_m2_16_8_i,temp_b2_14_6_r,temp_b2_14_6_i,temp_b2_14_8_r,temp_b2_14_8_i,temp_b2_16_6_r,temp_b2_16_6_i,temp_b2_16_8_r,temp_b2_16_8_i);
MULT MULT361 (clk,temp_b1_13_9_r,temp_b1_13_9_i,temp_b1_13_11_r,temp_b1_13_11_i,temp_b1_15_9_r,temp_b1_15_9_i,temp_b1_15_11_r,temp_b1_15_11_i,temp_m2_13_9_r,temp_m2_13_9_i,temp_m2_13_11_r,temp_m2_13_11_i,temp_m2_15_9_r,temp_m2_15_9_i,temp_m2_15_11_r,temp_m2_15_11_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly361 (clk,temp_m2_13_9_r,temp_m2_13_9_i,temp_m2_13_11_r,temp_m2_13_11_i,temp_m2_15_9_r,temp_m2_15_9_i,temp_m2_15_11_r,temp_m2_15_11_i,temp_b2_13_9_r,temp_b2_13_9_i,temp_b2_13_11_r,temp_b2_13_11_i,temp_b2_15_9_r,temp_b2_15_9_i,temp_b2_15_11_r,temp_b2_15_11_i);
MULT MULT362 (clk,temp_b1_13_10_r,temp_b1_13_10_i,temp_b1_13_12_r,temp_b1_13_12_i,temp_b1_15_10_r,temp_b1_15_10_i,temp_b1_15_12_r,temp_b1_15_12_i,temp_m2_13_10_r,temp_m2_13_10_i,temp_m2_13_12_r,temp_m2_13_12_i,temp_m2_15_10_r,temp_m2_15_10_i,temp_m2_15_12_r,temp_m2_15_12_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly362 (clk,temp_m2_13_10_r,temp_m2_13_10_i,temp_m2_13_12_r,temp_m2_13_12_i,temp_m2_15_10_r,temp_m2_15_10_i,temp_m2_15_12_r,temp_m2_15_12_i,temp_b2_13_10_r,temp_b2_13_10_i,temp_b2_13_12_r,temp_b2_13_12_i,temp_b2_15_10_r,temp_b2_15_10_i,temp_b2_15_12_r,temp_b2_15_12_i);
MULT MULT363 (clk,temp_b1_14_9_r,temp_b1_14_9_i,temp_b1_14_11_r,temp_b1_14_11_i,temp_b1_16_9_r,temp_b1_16_9_i,temp_b1_16_11_r,temp_b1_16_11_i,temp_m2_14_9_r,temp_m2_14_9_i,temp_m2_14_11_r,temp_m2_14_11_i,temp_m2_16_9_r,temp_m2_16_9_i,temp_m2_16_11_r,temp_m2_16_11_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly363 (clk,temp_m2_14_9_r,temp_m2_14_9_i,temp_m2_14_11_r,temp_m2_14_11_i,temp_m2_16_9_r,temp_m2_16_9_i,temp_m2_16_11_r,temp_m2_16_11_i,temp_b2_14_9_r,temp_b2_14_9_i,temp_b2_14_11_r,temp_b2_14_11_i,temp_b2_16_9_r,temp_b2_16_9_i,temp_b2_16_11_r,temp_b2_16_11_i);
MULT MULT364 (clk,temp_b1_14_10_r,temp_b1_14_10_i,temp_b1_14_12_r,temp_b1_14_12_i,temp_b1_16_10_r,temp_b1_16_10_i,temp_b1_16_12_r,temp_b1_16_12_i,temp_m2_14_10_r,temp_m2_14_10_i,temp_m2_14_12_r,temp_m2_14_12_i,temp_m2_16_10_r,temp_m2_16_10_i,temp_m2_16_12_r,temp_m2_16_12_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly364 (clk,temp_m2_14_10_r,temp_m2_14_10_i,temp_m2_14_12_r,temp_m2_14_12_i,temp_m2_16_10_r,temp_m2_16_10_i,temp_m2_16_12_r,temp_m2_16_12_i,temp_b2_14_10_r,temp_b2_14_10_i,temp_b2_14_12_r,temp_b2_14_12_i,temp_b2_16_10_r,temp_b2_16_10_i,temp_b2_16_12_r,temp_b2_16_12_i);
MULT MULT365 (clk,temp_b1_13_13_r,temp_b1_13_13_i,temp_b1_13_15_r,temp_b1_13_15_i,temp_b1_15_13_r,temp_b1_15_13_i,temp_b1_15_15_r,temp_b1_15_15_i,temp_m2_13_13_r,temp_m2_13_13_i,temp_m2_13_15_r,temp_m2_13_15_i,temp_m2_15_13_r,temp_m2_15_13_i,temp_m2_15_15_r,temp_m2_15_15_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly365 (clk,temp_m2_13_13_r,temp_m2_13_13_i,temp_m2_13_15_r,temp_m2_13_15_i,temp_m2_15_13_r,temp_m2_15_13_i,temp_m2_15_15_r,temp_m2_15_15_i,temp_b2_13_13_r,temp_b2_13_13_i,temp_b2_13_15_r,temp_b2_13_15_i,temp_b2_15_13_r,temp_b2_15_13_i,temp_b2_15_15_r,temp_b2_15_15_i);
MULT MULT366 (clk,temp_b1_13_14_r,temp_b1_13_14_i,temp_b1_13_16_r,temp_b1_13_16_i,temp_b1_15_14_r,temp_b1_15_14_i,temp_b1_15_16_r,temp_b1_15_16_i,temp_m2_13_14_r,temp_m2_13_14_i,temp_m2_13_16_r,temp_m2_13_16_i,temp_m2_15_14_r,temp_m2_15_14_i,temp_m2_15_16_r,temp_m2_15_16_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly366 (clk,temp_m2_13_14_r,temp_m2_13_14_i,temp_m2_13_16_r,temp_m2_13_16_i,temp_m2_15_14_r,temp_m2_15_14_i,temp_m2_15_16_r,temp_m2_15_16_i,temp_b2_13_14_r,temp_b2_13_14_i,temp_b2_13_16_r,temp_b2_13_16_i,temp_b2_15_14_r,temp_b2_15_14_i,temp_b2_15_16_r,temp_b2_15_16_i);
MULT MULT367 (clk,temp_b1_14_13_r,temp_b1_14_13_i,temp_b1_14_15_r,temp_b1_14_15_i,temp_b1_16_13_r,temp_b1_16_13_i,temp_b1_16_15_r,temp_b1_16_15_i,temp_m2_14_13_r,temp_m2_14_13_i,temp_m2_14_15_r,temp_m2_14_15_i,temp_m2_16_13_r,temp_m2_16_13_i,temp_m2_16_15_r,temp_m2_16_15_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly367 (clk,temp_m2_14_13_r,temp_m2_14_13_i,temp_m2_14_15_r,temp_m2_14_15_i,temp_m2_16_13_r,temp_m2_16_13_i,temp_m2_16_15_r,temp_m2_16_15_i,temp_b2_14_13_r,temp_b2_14_13_i,temp_b2_14_15_r,temp_b2_14_15_i,temp_b2_16_13_r,temp_b2_16_13_i,temp_b2_16_15_r,temp_b2_16_15_i);
MULT MULT368 (clk,temp_b1_14_14_r,temp_b1_14_14_i,temp_b1_14_16_r,temp_b1_14_16_i,temp_b1_16_14_r,temp_b1_16_14_i,temp_b1_16_16_r,temp_b1_16_16_i,temp_m2_14_14_r,temp_m2_14_14_i,temp_m2_14_16_r,temp_m2_14_16_i,temp_m2_16_14_r,temp_m2_16_14_i,temp_m2_16_16_r,temp_m2_16_16_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly368 (clk,temp_m2_14_14_r,temp_m2_14_14_i,temp_m2_14_16_r,temp_m2_14_16_i,temp_m2_16_14_r,temp_m2_16_14_i,temp_m2_16_16_r,temp_m2_16_16_i,temp_b2_14_14_r,temp_b2_14_14_i,temp_b2_14_16_r,temp_b2_14_16_i,temp_b2_16_14_r,temp_b2_16_14_i,temp_b2_16_16_r,temp_b2_16_16_i);
MULT MULT369 (clk,temp_b1_13_17_r,temp_b1_13_17_i,temp_b1_13_19_r,temp_b1_13_19_i,temp_b1_15_17_r,temp_b1_15_17_i,temp_b1_15_19_r,temp_b1_15_19_i,temp_m2_13_17_r,temp_m2_13_17_i,temp_m2_13_19_r,temp_m2_13_19_i,temp_m2_15_17_r,temp_m2_15_17_i,temp_m2_15_19_r,temp_m2_15_19_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly369 (clk,temp_m2_13_17_r,temp_m2_13_17_i,temp_m2_13_19_r,temp_m2_13_19_i,temp_m2_15_17_r,temp_m2_15_17_i,temp_m2_15_19_r,temp_m2_15_19_i,temp_b2_13_17_r,temp_b2_13_17_i,temp_b2_13_19_r,temp_b2_13_19_i,temp_b2_15_17_r,temp_b2_15_17_i,temp_b2_15_19_r,temp_b2_15_19_i);
MULT MULT370 (clk,temp_b1_13_18_r,temp_b1_13_18_i,temp_b1_13_20_r,temp_b1_13_20_i,temp_b1_15_18_r,temp_b1_15_18_i,temp_b1_15_20_r,temp_b1_15_20_i,temp_m2_13_18_r,temp_m2_13_18_i,temp_m2_13_20_r,temp_m2_13_20_i,temp_m2_15_18_r,temp_m2_15_18_i,temp_m2_15_20_r,temp_m2_15_20_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly370 (clk,temp_m2_13_18_r,temp_m2_13_18_i,temp_m2_13_20_r,temp_m2_13_20_i,temp_m2_15_18_r,temp_m2_15_18_i,temp_m2_15_20_r,temp_m2_15_20_i,temp_b2_13_18_r,temp_b2_13_18_i,temp_b2_13_20_r,temp_b2_13_20_i,temp_b2_15_18_r,temp_b2_15_18_i,temp_b2_15_20_r,temp_b2_15_20_i);
MULT MULT371 (clk,temp_b1_14_17_r,temp_b1_14_17_i,temp_b1_14_19_r,temp_b1_14_19_i,temp_b1_16_17_r,temp_b1_16_17_i,temp_b1_16_19_r,temp_b1_16_19_i,temp_m2_14_17_r,temp_m2_14_17_i,temp_m2_14_19_r,temp_m2_14_19_i,temp_m2_16_17_r,temp_m2_16_17_i,temp_m2_16_19_r,temp_m2_16_19_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly371 (clk,temp_m2_14_17_r,temp_m2_14_17_i,temp_m2_14_19_r,temp_m2_14_19_i,temp_m2_16_17_r,temp_m2_16_17_i,temp_m2_16_19_r,temp_m2_16_19_i,temp_b2_14_17_r,temp_b2_14_17_i,temp_b2_14_19_r,temp_b2_14_19_i,temp_b2_16_17_r,temp_b2_16_17_i,temp_b2_16_19_r,temp_b2_16_19_i);
MULT MULT372 (clk,temp_b1_14_18_r,temp_b1_14_18_i,temp_b1_14_20_r,temp_b1_14_20_i,temp_b1_16_18_r,temp_b1_16_18_i,temp_b1_16_20_r,temp_b1_16_20_i,temp_m2_14_18_r,temp_m2_14_18_i,temp_m2_14_20_r,temp_m2_14_20_i,temp_m2_16_18_r,temp_m2_16_18_i,temp_m2_16_20_r,temp_m2_16_20_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly372 (clk,temp_m2_14_18_r,temp_m2_14_18_i,temp_m2_14_20_r,temp_m2_14_20_i,temp_m2_16_18_r,temp_m2_16_18_i,temp_m2_16_20_r,temp_m2_16_20_i,temp_b2_14_18_r,temp_b2_14_18_i,temp_b2_14_20_r,temp_b2_14_20_i,temp_b2_16_18_r,temp_b2_16_18_i,temp_b2_16_20_r,temp_b2_16_20_i);
MULT MULT373 (clk,temp_b1_13_21_r,temp_b1_13_21_i,temp_b1_13_23_r,temp_b1_13_23_i,temp_b1_15_21_r,temp_b1_15_21_i,temp_b1_15_23_r,temp_b1_15_23_i,temp_m2_13_21_r,temp_m2_13_21_i,temp_m2_13_23_r,temp_m2_13_23_i,temp_m2_15_21_r,temp_m2_15_21_i,temp_m2_15_23_r,temp_m2_15_23_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly373 (clk,temp_m2_13_21_r,temp_m2_13_21_i,temp_m2_13_23_r,temp_m2_13_23_i,temp_m2_15_21_r,temp_m2_15_21_i,temp_m2_15_23_r,temp_m2_15_23_i,temp_b2_13_21_r,temp_b2_13_21_i,temp_b2_13_23_r,temp_b2_13_23_i,temp_b2_15_21_r,temp_b2_15_21_i,temp_b2_15_23_r,temp_b2_15_23_i);
MULT MULT374 (clk,temp_b1_13_22_r,temp_b1_13_22_i,temp_b1_13_24_r,temp_b1_13_24_i,temp_b1_15_22_r,temp_b1_15_22_i,temp_b1_15_24_r,temp_b1_15_24_i,temp_m2_13_22_r,temp_m2_13_22_i,temp_m2_13_24_r,temp_m2_13_24_i,temp_m2_15_22_r,temp_m2_15_22_i,temp_m2_15_24_r,temp_m2_15_24_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly374 (clk,temp_m2_13_22_r,temp_m2_13_22_i,temp_m2_13_24_r,temp_m2_13_24_i,temp_m2_15_22_r,temp_m2_15_22_i,temp_m2_15_24_r,temp_m2_15_24_i,temp_b2_13_22_r,temp_b2_13_22_i,temp_b2_13_24_r,temp_b2_13_24_i,temp_b2_15_22_r,temp_b2_15_22_i,temp_b2_15_24_r,temp_b2_15_24_i);
MULT MULT375 (clk,temp_b1_14_21_r,temp_b1_14_21_i,temp_b1_14_23_r,temp_b1_14_23_i,temp_b1_16_21_r,temp_b1_16_21_i,temp_b1_16_23_r,temp_b1_16_23_i,temp_m2_14_21_r,temp_m2_14_21_i,temp_m2_14_23_r,temp_m2_14_23_i,temp_m2_16_21_r,temp_m2_16_21_i,temp_m2_16_23_r,temp_m2_16_23_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly375 (clk,temp_m2_14_21_r,temp_m2_14_21_i,temp_m2_14_23_r,temp_m2_14_23_i,temp_m2_16_21_r,temp_m2_16_21_i,temp_m2_16_23_r,temp_m2_16_23_i,temp_b2_14_21_r,temp_b2_14_21_i,temp_b2_14_23_r,temp_b2_14_23_i,temp_b2_16_21_r,temp_b2_16_21_i,temp_b2_16_23_r,temp_b2_16_23_i);
MULT MULT376 (clk,temp_b1_14_22_r,temp_b1_14_22_i,temp_b1_14_24_r,temp_b1_14_24_i,temp_b1_16_22_r,temp_b1_16_22_i,temp_b1_16_24_r,temp_b1_16_24_i,temp_m2_14_22_r,temp_m2_14_22_i,temp_m2_14_24_r,temp_m2_14_24_i,temp_m2_16_22_r,temp_m2_16_22_i,temp_m2_16_24_r,temp_m2_16_24_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly376 (clk,temp_m2_14_22_r,temp_m2_14_22_i,temp_m2_14_24_r,temp_m2_14_24_i,temp_m2_16_22_r,temp_m2_16_22_i,temp_m2_16_24_r,temp_m2_16_24_i,temp_b2_14_22_r,temp_b2_14_22_i,temp_b2_14_24_r,temp_b2_14_24_i,temp_b2_16_22_r,temp_b2_16_22_i,temp_b2_16_24_r,temp_b2_16_24_i);
MULT MULT377 (clk,temp_b1_13_25_r,temp_b1_13_25_i,temp_b1_13_27_r,temp_b1_13_27_i,temp_b1_15_25_r,temp_b1_15_25_i,temp_b1_15_27_r,temp_b1_15_27_i,temp_m2_13_25_r,temp_m2_13_25_i,temp_m2_13_27_r,temp_m2_13_27_i,temp_m2_15_25_r,temp_m2_15_25_i,temp_m2_15_27_r,temp_m2_15_27_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly377 (clk,temp_m2_13_25_r,temp_m2_13_25_i,temp_m2_13_27_r,temp_m2_13_27_i,temp_m2_15_25_r,temp_m2_15_25_i,temp_m2_15_27_r,temp_m2_15_27_i,temp_b2_13_25_r,temp_b2_13_25_i,temp_b2_13_27_r,temp_b2_13_27_i,temp_b2_15_25_r,temp_b2_15_25_i,temp_b2_15_27_r,temp_b2_15_27_i);
MULT MULT378 (clk,temp_b1_13_26_r,temp_b1_13_26_i,temp_b1_13_28_r,temp_b1_13_28_i,temp_b1_15_26_r,temp_b1_15_26_i,temp_b1_15_28_r,temp_b1_15_28_i,temp_m2_13_26_r,temp_m2_13_26_i,temp_m2_13_28_r,temp_m2_13_28_i,temp_m2_15_26_r,temp_m2_15_26_i,temp_m2_15_28_r,temp_m2_15_28_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly378 (clk,temp_m2_13_26_r,temp_m2_13_26_i,temp_m2_13_28_r,temp_m2_13_28_i,temp_m2_15_26_r,temp_m2_15_26_i,temp_m2_15_28_r,temp_m2_15_28_i,temp_b2_13_26_r,temp_b2_13_26_i,temp_b2_13_28_r,temp_b2_13_28_i,temp_b2_15_26_r,temp_b2_15_26_i,temp_b2_15_28_r,temp_b2_15_28_i);
MULT MULT379 (clk,temp_b1_14_25_r,temp_b1_14_25_i,temp_b1_14_27_r,temp_b1_14_27_i,temp_b1_16_25_r,temp_b1_16_25_i,temp_b1_16_27_r,temp_b1_16_27_i,temp_m2_14_25_r,temp_m2_14_25_i,temp_m2_14_27_r,temp_m2_14_27_i,temp_m2_16_25_r,temp_m2_16_25_i,temp_m2_16_27_r,temp_m2_16_27_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly379 (clk,temp_m2_14_25_r,temp_m2_14_25_i,temp_m2_14_27_r,temp_m2_14_27_i,temp_m2_16_25_r,temp_m2_16_25_i,temp_m2_16_27_r,temp_m2_16_27_i,temp_b2_14_25_r,temp_b2_14_25_i,temp_b2_14_27_r,temp_b2_14_27_i,temp_b2_16_25_r,temp_b2_16_25_i,temp_b2_16_27_r,temp_b2_16_27_i);
MULT MULT380 (clk,temp_b1_14_26_r,temp_b1_14_26_i,temp_b1_14_28_r,temp_b1_14_28_i,temp_b1_16_26_r,temp_b1_16_26_i,temp_b1_16_28_r,temp_b1_16_28_i,temp_m2_14_26_r,temp_m2_14_26_i,temp_m2_14_28_r,temp_m2_14_28_i,temp_m2_16_26_r,temp_m2_16_26_i,temp_m2_16_28_r,temp_m2_16_28_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly380 (clk,temp_m2_14_26_r,temp_m2_14_26_i,temp_m2_14_28_r,temp_m2_14_28_i,temp_m2_16_26_r,temp_m2_16_26_i,temp_m2_16_28_r,temp_m2_16_28_i,temp_b2_14_26_r,temp_b2_14_26_i,temp_b2_14_28_r,temp_b2_14_28_i,temp_b2_16_26_r,temp_b2_16_26_i,temp_b2_16_28_r,temp_b2_16_28_i);
MULT MULT381 (clk,temp_b1_13_29_r,temp_b1_13_29_i,temp_b1_13_31_r,temp_b1_13_31_i,temp_b1_15_29_r,temp_b1_15_29_i,temp_b1_15_31_r,temp_b1_15_31_i,temp_m2_13_29_r,temp_m2_13_29_i,temp_m2_13_31_r,temp_m2_13_31_i,temp_m2_15_29_r,temp_m2_15_29_i,temp_m2_15_31_r,temp_m2_15_31_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly381 (clk,temp_m2_13_29_r,temp_m2_13_29_i,temp_m2_13_31_r,temp_m2_13_31_i,temp_m2_15_29_r,temp_m2_15_29_i,temp_m2_15_31_r,temp_m2_15_31_i,temp_b2_13_29_r,temp_b2_13_29_i,temp_b2_13_31_r,temp_b2_13_31_i,temp_b2_15_29_r,temp_b2_15_29_i,temp_b2_15_31_r,temp_b2_15_31_i);
MULT MULT382 (clk,temp_b1_13_30_r,temp_b1_13_30_i,temp_b1_13_32_r,temp_b1_13_32_i,temp_b1_15_30_r,temp_b1_15_30_i,temp_b1_15_32_r,temp_b1_15_32_i,temp_m2_13_30_r,temp_m2_13_30_i,temp_m2_13_32_r,temp_m2_13_32_i,temp_m2_15_30_r,temp_m2_15_30_i,temp_m2_15_32_r,temp_m2_15_32_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly382 (clk,temp_m2_13_30_r,temp_m2_13_30_i,temp_m2_13_32_r,temp_m2_13_32_i,temp_m2_15_30_r,temp_m2_15_30_i,temp_m2_15_32_r,temp_m2_15_32_i,temp_b2_13_30_r,temp_b2_13_30_i,temp_b2_13_32_r,temp_b2_13_32_i,temp_b2_15_30_r,temp_b2_15_30_i,temp_b2_15_32_r,temp_b2_15_32_i);
MULT MULT383 (clk,temp_b1_14_29_r,temp_b1_14_29_i,temp_b1_14_31_r,temp_b1_14_31_i,temp_b1_16_29_r,temp_b1_16_29_i,temp_b1_16_31_r,temp_b1_16_31_i,temp_m2_14_29_r,temp_m2_14_29_i,temp_m2_14_31_r,temp_m2_14_31_i,temp_m2_16_29_r,temp_m2_16_29_i,temp_m2_16_31_r,temp_m2_16_31_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly383 (clk,temp_m2_14_29_r,temp_m2_14_29_i,temp_m2_14_31_r,temp_m2_14_31_i,temp_m2_16_29_r,temp_m2_16_29_i,temp_m2_16_31_r,temp_m2_16_31_i,temp_b2_14_29_r,temp_b2_14_29_i,temp_b2_14_31_r,temp_b2_14_31_i,temp_b2_16_29_r,temp_b2_16_29_i,temp_b2_16_31_r,temp_b2_16_31_i);
MULT MULT384 (clk,temp_b1_14_30_r,temp_b1_14_30_i,temp_b1_14_32_r,temp_b1_14_32_i,temp_b1_16_30_r,temp_b1_16_30_i,temp_b1_16_32_r,temp_b1_16_32_i,temp_m2_14_30_r,temp_m2_14_30_i,temp_m2_14_32_r,temp_m2_14_32_i,temp_m2_16_30_r,temp_m2_16_30_i,temp_m2_16_32_r,temp_m2_16_32_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly384 (clk,temp_m2_14_30_r,temp_m2_14_30_i,temp_m2_14_32_r,temp_m2_14_32_i,temp_m2_16_30_r,temp_m2_16_30_i,temp_m2_16_32_r,temp_m2_16_32_i,temp_b2_14_30_r,temp_b2_14_30_i,temp_b2_14_32_r,temp_b2_14_32_i,temp_b2_16_30_r,temp_b2_16_30_i,temp_b2_16_32_r,temp_b2_16_32_i);
MULT MULT385 (clk,temp_b1_17_1_r,temp_b1_17_1_i,temp_b1_17_3_r,temp_b1_17_3_i,temp_b1_19_1_r,temp_b1_19_1_i,temp_b1_19_3_r,temp_b1_19_3_i,temp_m2_17_1_r,temp_m2_17_1_i,temp_m2_17_3_r,temp_m2_17_3_i,temp_m2_19_1_r,temp_m2_19_1_i,temp_m2_19_3_r,temp_m2_19_3_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly385 (clk,temp_m2_17_1_r,temp_m2_17_1_i,temp_m2_17_3_r,temp_m2_17_3_i,temp_m2_19_1_r,temp_m2_19_1_i,temp_m2_19_3_r,temp_m2_19_3_i,temp_b2_17_1_r,temp_b2_17_1_i,temp_b2_17_3_r,temp_b2_17_3_i,temp_b2_19_1_r,temp_b2_19_1_i,temp_b2_19_3_r,temp_b2_19_3_i);
MULT MULT386 (clk,temp_b1_17_2_r,temp_b1_17_2_i,temp_b1_17_4_r,temp_b1_17_4_i,temp_b1_19_2_r,temp_b1_19_2_i,temp_b1_19_4_r,temp_b1_19_4_i,temp_m2_17_2_r,temp_m2_17_2_i,temp_m2_17_4_r,temp_m2_17_4_i,temp_m2_19_2_r,temp_m2_19_2_i,temp_m2_19_4_r,temp_m2_19_4_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly386 (clk,temp_m2_17_2_r,temp_m2_17_2_i,temp_m2_17_4_r,temp_m2_17_4_i,temp_m2_19_2_r,temp_m2_19_2_i,temp_m2_19_4_r,temp_m2_19_4_i,temp_b2_17_2_r,temp_b2_17_2_i,temp_b2_17_4_r,temp_b2_17_4_i,temp_b2_19_2_r,temp_b2_19_2_i,temp_b2_19_4_r,temp_b2_19_4_i);
MULT MULT387 (clk,temp_b1_18_1_r,temp_b1_18_1_i,temp_b1_18_3_r,temp_b1_18_3_i,temp_b1_20_1_r,temp_b1_20_1_i,temp_b1_20_3_r,temp_b1_20_3_i,temp_m2_18_1_r,temp_m2_18_1_i,temp_m2_18_3_r,temp_m2_18_3_i,temp_m2_20_1_r,temp_m2_20_1_i,temp_m2_20_3_r,temp_m2_20_3_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly387 (clk,temp_m2_18_1_r,temp_m2_18_1_i,temp_m2_18_3_r,temp_m2_18_3_i,temp_m2_20_1_r,temp_m2_20_1_i,temp_m2_20_3_r,temp_m2_20_3_i,temp_b2_18_1_r,temp_b2_18_1_i,temp_b2_18_3_r,temp_b2_18_3_i,temp_b2_20_1_r,temp_b2_20_1_i,temp_b2_20_3_r,temp_b2_20_3_i);
MULT MULT388 (clk,temp_b1_18_2_r,temp_b1_18_2_i,temp_b1_18_4_r,temp_b1_18_4_i,temp_b1_20_2_r,temp_b1_20_2_i,temp_b1_20_4_r,temp_b1_20_4_i,temp_m2_18_2_r,temp_m2_18_2_i,temp_m2_18_4_r,temp_m2_18_4_i,temp_m2_20_2_r,temp_m2_20_2_i,temp_m2_20_4_r,temp_m2_20_4_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly388 (clk,temp_m2_18_2_r,temp_m2_18_2_i,temp_m2_18_4_r,temp_m2_18_4_i,temp_m2_20_2_r,temp_m2_20_2_i,temp_m2_20_4_r,temp_m2_20_4_i,temp_b2_18_2_r,temp_b2_18_2_i,temp_b2_18_4_r,temp_b2_18_4_i,temp_b2_20_2_r,temp_b2_20_2_i,temp_b2_20_4_r,temp_b2_20_4_i);
MULT MULT389 (clk,temp_b1_17_5_r,temp_b1_17_5_i,temp_b1_17_7_r,temp_b1_17_7_i,temp_b1_19_5_r,temp_b1_19_5_i,temp_b1_19_7_r,temp_b1_19_7_i,temp_m2_17_5_r,temp_m2_17_5_i,temp_m2_17_7_r,temp_m2_17_7_i,temp_m2_19_5_r,temp_m2_19_5_i,temp_m2_19_7_r,temp_m2_19_7_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly389 (clk,temp_m2_17_5_r,temp_m2_17_5_i,temp_m2_17_7_r,temp_m2_17_7_i,temp_m2_19_5_r,temp_m2_19_5_i,temp_m2_19_7_r,temp_m2_19_7_i,temp_b2_17_5_r,temp_b2_17_5_i,temp_b2_17_7_r,temp_b2_17_7_i,temp_b2_19_5_r,temp_b2_19_5_i,temp_b2_19_7_r,temp_b2_19_7_i);
MULT MULT390 (clk,temp_b1_17_6_r,temp_b1_17_6_i,temp_b1_17_8_r,temp_b1_17_8_i,temp_b1_19_6_r,temp_b1_19_6_i,temp_b1_19_8_r,temp_b1_19_8_i,temp_m2_17_6_r,temp_m2_17_6_i,temp_m2_17_8_r,temp_m2_17_8_i,temp_m2_19_6_r,temp_m2_19_6_i,temp_m2_19_8_r,temp_m2_19_8_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly390 (clk,temp_m2_17_6_r,temp_m2_17_6_i,temp_m2_17_8_r,temp_m2_17_8_i,temp_m2_19_6_r,temp_m2_19_6_i,temp_m2_19_8_r,temp_m2_19_8_i,temp_b2_17_6_r,temp_b2_17_6_i,temp_b2_17_8_r,temp_b2_17_8_i,temp_b2_19_6_r,temp_b2_19_6_i,temp_b2_19_8_r,temp_b2_19_8_i);
MULT MULT391 (clk,temp_b1_18_5_r,temp_b1_18_5_i,temp_b1_18_7_r,temp_b1_18_7_i,temp_b1_20_5_r,temp_b1_20_5_i,temp_b1_20_7_r,temp_b1_20_7_i,temp_m2_18_5_r,temp_m2_18_5_i,temp_m2_18_7_r,temp_m2_18_7_i,temp_m2_20_5_r,temp_m2_20_5_i,temp_m2_20_7_r,temp_m2_20_7_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly391 (clk,temp_m2_18_5_r,temp_m2_18_5_i,temp_m2_18_7_r,temp_m2_18_7_i,temp_m2_20_5_r,temp_m2_20_5_i,temp_m2_20_7_r,temp_m2_20_7_i,temp_b2_18_5_r,temp_b2_18_5_i,temp_b2_18_7_r,temp_b2_18_7_i,temp_b2_20_5_r,temp_b2_20_5_i,temp_b2_20_7_r,temp_b2_20_7_i);
MULT MULT392 (clk,temp_b1_18_6_r,temp_b1_18_6_i,temp_b1_18_8_r,temp_b1_18_8_i,temp_b1_20_6_r,temp_b1_20_6_i,temp_b1_20_8_r,temp_b1_20_8_i,temp_m2_18_6_r,temp_m2_18_6_i,temp_m2_18_8_r,temp_m2_18_8_i,temp_m2_20_6_r,temp_m2_20_6_i,temp_m2_20_8_r,temp_m2_20_8_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly392 (clk,temp_m2_18_6_r,temp_m2_18_6_i,temp_m2_18_8_r,temp_m2_18_8_i,temp_m2_20_6_r,temp_m2_20_6_i,temp_m2_20_8_r,temp_m2_20_8_i,temp_b2_18_6_r,temp_b2_18_6_i,temp_b2_18_8_r,temp_b2_18_8_i,temp_b2_20_6_r,temp_b2_20_6_i,temp_b2_20_8_r,temp_b2_20_8_i);
MULT MULT393 (clk,temp_b1_17_9_r,temp_b1_17_9_i,temp_b1_17_11_r,temp_b1_17_11_i,temp_b1_19_9_r,temp_b1_19_9_i,temp_b1_19_11_r,temp_b1_19_11_i,temp_m2_17_9_r,temp_m2_17_9_i,temp_m2_17_11_r,temp_m2_17_11_i,temp_m2_19_9_r,temp_m2_19_9_i,temp_m2_19_11_r,temp_m2_19_11_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly393 (clk,temp_m2_17_9_r,temp_m2_17_9_i,temp_m2_17_11_r,temp_m2_17_11_i,temp_m2_19_9_r,temp_m2_19_9_i,temp_m2_19_11_r,temp_m2_19_11_i,temp_b2_17_9_r,temp_b2_17_9_i,temp_b2_17_11_r,temp_b2_17_11_i,temp_b2_19_9_r,temp_b2_19_9_i,temp_b2_19_11_r,temp_b2_19_11_i);
MULT MULT394 (clk,temp_b1_17_10_r,temp_b1_17_10_i,temp_b1_17_12_r,temp_b1_17_12_i,temp_b1_19_10_r,temp_b1_19_10_i,temp_b1_19_12_r,temp_b1_19_12_i,temp_m2_17_10_r,temp_m2_17_10_i,temp_m2_17_12_r,temp_m2_17_12_i,temp_m2_19_10_r,temp_m2_19_10_i,temp_m2_19_12_r,temp_m2_19_12_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly394 (clk,temp_m2_17_10_r,temp_m2_17_10_i,temp_m2_17_12_r,temp_m2_17_12_i,temp_m2_19_10_r,temp_m2_19_10_i,temp_m2_19_12_r,temp_m2_19_12_i,temp_b2_17_10_r,temp_b2_17_10_i,temp_b2_17_12_r,temp_b2_17_12_i,temp_b2_19_10_r,temp_b2_19_10_i,temp_b2_19_12_r,temp_b2_19_12_i);
MULT MULT395 (clk,temp_b1_18_9_r,temp_b1_18_9_i,temp_b1_18_11_r,temp_b1_18_11_i,temp_b1_20_9_r,temp_b1_20_9_i,temp_b1_20_11_r,temp_b1_20_11_i,temp_m2_18_9_r,temp_m2_18_9_i,temp_m2_18_11_r,temp_m2_18_11_i,temp_m2_20_9_r,temp_m2_20_9_i,temp_m2_20_11_r,temp_m2_20_11_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly395 (clk,temp_m2_18_9_r,temp_m2_18_9_i,temp_m2_18_11_r,temp_m2_18_11_i,temp_m2_20_9_r,temp_m2_20_9_i,temp_m2_20_11_r,temp_m2_20_11_i,temp_b2_18_9_r,temp_b2_18_9_i,temp_b2_18_11_r,temp_b2_18_11_i,temp_b2_20_9_r,temp_b2_20_9_i,temp_b2_20_11_r,temp_b2_20_11_i);
MULT MULT396 (clk,temp_b1_18_10_r,temp_b1_18_10_i,temp_b1_18_12_r,temp_b1_18_12_i,temp_b1_20_10_r,temp_b1_20_10_i,temp_b1_20_12_r,temp_b1_20_12_i,temp_m2_18_10_r,temp_m2_18_10_i,temp_m2_18_12_r,temp_m2_18_12_i,temp_m2_20_10_r,temp_m2_20_10_i,temp_m2_20_12_r,temp_m2_20_12_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly396 (clk,temp_m2_18_10_r,temp_m2_18_10_i,temp_m2_18_12_r,temp_m2_18_12_i,temp_m2_20_10_r,temp_m2_20_10_i,temp_m2_20_12_r,temp_m2_20_12_i,temp_b2_18_10_r,temp_b2_18_10_i,temp_b2_18_12_r,temp_b2_18_12_i,temp_b2_20_10_r,temp_b2_20_10_i,temp_b2_20_12_r,temp_b2_20_12_i);
MULT MULT397 (clk,temp_b1_17_13_r,temp_b1_17_13_i,temp_b1_17_15_r,temp_b1_17_15_i,temp_b1_19_13_r,temp_b1_19_13_i,temp_b1_19_15_r,temp_b1_19_15_i,temp_m2_17_13_r,temp_m2_17_13_i,temp_m2_17_15_r,temp_m2_17_15_i,temp_m2_19_13_r,temp_m2_19_13_i,temp_m2_19_15_r,temp_m2_19_15_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly397 (clk,temp_m2_17_13_r,temp_m2_17_13_i,temp_m2_17_15_r,temp_m2_17_15_i,temp_m2_19_13_r,temp_m2_19_13_i,temp_m2_19_15_r,temp_m2_19_15_i,temp_b2_17_13_r,temp_b2_17_13_i,temp_b2_17_15_r,temp_b2_17_15_i,temp_b2_19_13_r,temp_b2_19_13_i,temp_b2_19_15_r,temp_b2_19_15_i);
MULT MULT398 (clk,temp_b1_17_14_r,temp_b1_17_14_i,temp_b1_17_16_r,temp_b1_17_16_i,temp_b1_19_14_r,temp_b1_19_14_i,temp_b1_19_16_r,temp_b1_19_16_i,temp_m2_17_14_r,temp_m2_17_14_i,temp_m2_17_16_r,temp_m2_17_16_i,temp_m2_19_14_r,temp_m2_19_14_i,temp_m2_19_16_r,temp_m2_19_16_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly398 (clk,temp_m2_17_14_r,temp_m2_17_14_i,temp_m2_17_16_r,temp_m2_17_16_i,temp_m2_19_14_r,temp_m2_19_14_i,temp_m2_19_16_r,temp_m2_19_16_i,temp_b2_17_14_r,temp_b2_17_14_i,temp_b2_17_16_r,temp_b2_17_16_i,temp_b2_19_14_r,temp_b2_19_14_i,temp_b2_19_16_r,temp_b2_19_16_i);
MULT MULT399 (clk,temp_b1_18_13_r,temp_b1_18_13_i,temp_b1_18_15_r,temp_b1_18_15_i,temp_b1_20_13_r,temp_b1_20_13_i,temp_b1_20_15_r,temp_b1_20_15_i,temp_m2_18_13_r,temp_m2_18_13_i,temp_m2_18_15_r,temp_m2_18_15_i,temp_m2_20_13_r,temp_m2_20_13_i,temp_m2_20_15_r,temp_m2_20_15_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly399 (clk,temp_m2_18_13_r,temp_m2_18_13_i,temp_m2_18_15_r,temp_m2_18_15_i,temp_m2_20_13_r,temp_m2_20_13_i,temp_m2_20_15_r,temp_m2_20_15_i,temp_b2_18_13_r,temp_b2_18_13_i,temp_b2_18_15_r,temp_b2_18_15_i,temp_b2_20_13_r,temp_b2_20_13_i,temp_b2_20_15_r,temp_b2_20_15_i);
MULT MULT400 (clk,temp_b1_18_14_r,temp_b1_18_14_i,temp_b1_18_16_r,temp_b1_18_16_i,temp_b1_20_14_r,temp_b1_20_14_i,temp_b1_20_16_r,temp_b1_20_16_i,temp_m2_18_14_r,temp_m2_18_14_i,temp_m2_18_16_r,temp_m2_18_16_i,temp_m2_20_14_r,temp_m2_20_14_i,temp_m2_20_16_r,temp_m2_20_16_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly400 (clk,temp_m2_18_14_r,temp_m2_18_14_i,temp_m2_18_16_r,temp_m2_18_16_i,temp_m2_20_14_r,temp_m2_20_14_i,temp_m2_20_16_r,temp_m2_20_16_i,temp_b2_18_14_r,temp_b2_18_14_i,temp_b2_18_16_r,temp_b2_18_16_i,temp_b2_20_14_r,temp_b2_20_14_i,temp_b2_20_16_r,temp_b2_20_16_i);
MULT MULT401 (clk,temp_b1_17_17_r,temp_b1_17_17_i,temp_b1_17_19_r,temp_b1_17_19_i,temp_b1_19_17_r,temp_b1_19_17_i,temp_b1_19_19_r,temp_b1_19_19_i,temp_m2_17_17_r,temp_m2_17_17_i,temp_m2_17_19_r,temp_m2_17_19_i,temp_m2_19_17_r,temp_m2_19_17_i,temp_m2_19_19_r,temp_m2_19_19_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly401 (clk,temp_m2_17_17_r,temp_m2_17_17_i,temp_m2_17_19_r,temp_m2_17_19_i,temp_m2_19_17_r,temp_m2_19_17_i,temp_m2_19_19_r,temp_m2_19_19_i,temp_b2_17_17_r,temp_b2_17_17_i,temp_b2_17_19_r,temp_b2_17_19_i,temp_b2_19_17_r,temp_b2_19_17_i,temp_b2_19_19_r,temp_b2_19_19_i);
MULT MULT402 (clk,temp_b1_17_18_r,temp_b1_17_18_i,temp_b1_17_20_r,temp_b1_17_20_i,temp_b1_19_18_r,temp_b1_19_18_i,temp_b1_19_20_r,temp_b1_19_20_i,temp_m2_17_18_r,temp_m2_17_18_i,temp_m2_17_20_r,temp_m2_17_20_i,temp_m2_19_18_r,temp_m2_19_18_i,temp_m2_19_20_r,temp_m2_19_20_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly402 (clk,temp_m2_17_18_r,temp_m2_17_18_i,temp_m2_17_20_r,temp_m2_17_20_i,temp_m2_19_18_r,temp_m2_19_18_i,temp_m2_19_20_r,temp_m2_19_20_i,temp_b2_17_18_r,temp_b2_17_18_i,temp_b2_17_20_r,temp_b2_17_20_i,temp_b2_19_18_r,temp_b2_19_18_i,temp_b2_19_20_r,temp_b2_19_20_i);
MULT MULT403 (clk,temp_b1_18_17_r,temp_b1_18_17_i,temp_b1_18_19_r,temp_b1_18_19_i,temp_b1_20_17_r,temp_b1_20_17_i,temp_b1_20_19_r,temp_b1_20_19_i,temp_m2_18_17_r,temp_m2_18_17_i,temp_m2_18_19_r,temp_m2_18_19_i,temp_m2_20_17_r,temp_m2_20_17_i,temp_m2_20_19_r,temp_m2_20_19_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly403 (clk,temp_m2_18_17_r,temp_m2_18_17_i,temp_m2_18_19_r,temp_m2_18_19_i,temp_m2_20_17_r,temp_m2_20_17_i,temp_m2_20_19_r,temp_m2_20_19_i,temp_b2_18_17_r,temp_b2_18_17_i,temp_b2_18_19_r,temp_b2_18_19_i,temp_b2_20_17_r,temp_b2_20_17_i,temp_b2_20_19_r,temp_b2_20_19_i);
MULT MULT404 (clk,temp_b1_18_18_r,temp_b1_18_18_i,temp_b1_18_20_r,temp_b1_18_20_i,temp_b1_20_18_r,temp_b1_20_18_i,temp_b1_20_20_r,temp_b1_20_20_i,temp_m2_18_18_r,temp_m2_18_18_i,temp_m2_18_20_r,temp_m2_18_20_i,temp_m2_20_18_r,temp_m2_20_18_i,temp_m2_20_20_r,temp_m2_20_20_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly404 (clk,temp_m2_18_18_r,temp_m2_18_18_i,temp_m2_18_20_r,temp_m2_18_20_i,temp_m2_20_18_r,temp_m2_20_18_i,temp_m2_20_20_r,temp_m2_20_20_i,temp_b2_18_18_r,temp_b2_18_18_i,temp_b2_18_20_r,temp_b2_18_20_i,temp_b2_20_18_r,temp_b2_20_18_i,temp_b2_20_20_r,temp_b2_20_20_i);
MULT MULT405 (clk,temp_b1_17_21_r,temp_b1_17_21_i,temp_b1_17_23_r,temp_b1_17_23_i,temp_b1_19_21_r,temp_b1_19_21_i,temp_b1_19_23_r,temp_b1_19_23_i,temp_m2_17_21_r,temp_m2_17_21_i,temp_m2_17_23_r,temp_m2_17_23_i,temp_m2_19_21_r,temp_m2_19_21_i,temp_m2_19_23_r,temp_m2_19_23_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly405 (clk,temp_m2_17_21_r,temp_m2_17_21_i,temp_m2_17_23_r,temp_m2_17_23_i,temp_m2_19_21_r,temp_m2_19_21_i,temp_m2_19_23_r,temp_m2_19_23_i,temp_b2_17_21_r,temp_b2_17_21_i,temp_b2_17_23_r,temp_b2_17_23_i,temp_b2_19_21_r,temp_b2_19_21_i,temp_b2_19_23_r,temp_b2_19_23_i);
MULT MULT406 (clk,temp_b1_17_22_r,temp_b1_17_22_i,temp_b1_17_24_r,temp_b1_17_24_i,temp_b1_19_22_r,temp_b1_19_22_i,temp_b1_19_24_r,temp_b1_19_24_i,temp_m2_17_22_r,temp_m2_17_22_i,temp_m2_17_24_r,temp_m2_17_24_i,temp_m2_19_22_r,temp_m2_19_22_i,temp_m2_19_24_r,temp_m2_19_24_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly406 (clk,temp_m2_17_22_r,temp_m2_17_22_i,temp_m2_17_24_r,temp_m2_17_24_i,temp_m2_19_22_r,temp_m2_19_22_i,temp_m2_19_24_r,temp_m2_19_24_i,temp_b2_17_22_r,temp_b2_17_22_i,temp_b2_17_24_r,temp_b2_17_24_i,temp_b2_19_22_r,temp_b2_19_22_i,temp_b2_19_24_r,temp_b2_19_24_i);
MULT MULT407 (clk,temp_b1_18_21_r,temp_b1_18_21_i,temp_b1_18_23_r,temp_b1_18_23_i,temp_b1_20_21_r,temp_b1_20_21_i,temp_b1_20_23_r,temp_b1_20_23_i,temp_m2_18_21_r,temp_m2_18_21_i,temp_m2_18_23_r,temp_m2_18_23_i,temp_m2_20_21_r,temp_m2_20_21_i,temp_m2_20_23_r,temp_m2_20_23_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly407 (clk,temp_m2_18_21_r,temp_m2_18_21_i,temp_m2_18_23_r,temp_m2_18_23_i,temp_m2_20_21_r,temp_m2_20_21_i,temp_m2_20_23_r,temp_m2_20_23_i,temp_b2_18_21_r,temp_b2_18_21_i,temp_b2_18_23_r,temp_b2_18_23_i,temp_b2_20_21_r,temp_b2_20_21_i,temp_b2_20_23_r,temp_b2_20_23_i);
MULT MULT408 (clk,temp_b1_18_22_r,temp_b1_18_22_i,temp_b1_18_24_r,temp_b1_18_24_i,temp_b1_20_22_r,temp_b1_20_22_i,temp_b1_20_24_r,temp_b1_20_24_i,temp_m2_18_22_r,temp_m2_18_22_i,temp_m2_18_24_r,temp_m2_18_24_i,temp_m2_20_22_r,temp_m2_20_22_i,temp_m2_20_24_r,temp_m2_20_24_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly408 (clk,temp_m2_18_22_r,temp_m2_18_22_i,temp_m2_18_24_r,temp_m2_18_24_i,temp_m2_20_22_r,temp_m2_20_22_i,temp_m2_20_24_r,temp_m2_20_24_i,temp_b2_18_22_r,temp_b2_18_22_i,temp_b2_18_24_r,temp_b2_18_24_i,temp_b2_20_22_r,temp_b2_20_22_i,temp_b2_20_24_r,temp_b2_20_24_i);
MULT MULT409 (clk,temp_b1_17_25_r,temp_b1_17_25_i,temp_b1_17_27_r,temp_b1_17_27_i,temp_b1_19_25_r,temp_b1_19_25_i,temp_b1_19_27_r,temp_b1_19_27_i,temp_m2_17_25_r,temp_m2_17_25_i,temp_m2_17_27_r,temp_m2_17_27_i,temp_m2_19_25_r,temp_m2_19_25_i,temp_m2_19_27_r,temp_m2_19_27_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly409 (clk,temp_m2_17_25_r,temp_m2_17_25_i,temp_m2_17_27_r,temp_m2_17_27_i,temp_m2_19_25_r,temp_m2_19_25_i,temp_m2_19_27_r,temp_m2_19_27_i,temp_b2_17_25_r,temp_b2_17_25_i,temp_b2_17_27_r,temp_b2_17_27_i,temp_b2_19_25_r,temp_b2_19_25_i,temp_b2_19_27_r,temp_b2_19_27_i);
MULT MULT410 (clk,temp_b1_17_26_r,temp_b1_17_26_i,temp_b1_17_28_r,temp_b1_17_28_i,temp_b1_19_26_r,temp_b1_19_26_i,temp_b1_19_28_r,temp_b1_19_28_i,temp_m2_17_26_r,temp_m2_17_26_i,temp_m2_17_28_r,temp_m2_17_28_i,temp_m2_19_26_r,temp_m2_19_26_i,temp_m2_19_28_r,temp_m2_19_28_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly410 (clk,temp_m2_17_26_r,temp_m2_17_26_i,temp_m2_17_28_r,temp_m2_17_28_i,temp_m2_19_26_r,temp_m2_19_26_i,temp_m2_19_28_r,temp_m2_19_28_i,temp_b2_17_26_r,temp_b2_17_26_i,temp_b2_17_28_r,temp_b2_17_28_i,temp_b2_19_26_r,temp_b2_19_26_i,temp_b2_19_28_r,temp_b2_19_28_i);
MULT MULT411 (clk,temp_b1_18_25_r,temp_b1_18_25_i,temp_b1_18_27_r,temp_b1_18_27_i,temp_b1_20_25_r,temp_b1_20_25_i,temp_b1_20_27_r,temp_b1_20_27_i,temp_m2_18_25_r,temp_m2_18_25_i,temp_m2_18_27_r,temp_m2_18_27_i,temp_m2_20_25_r,temp_m2_20_25_i,temp_m2_20_27_r,temp_m2_20_27_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly411 (clk,temp_m2_18_25_r,temp_m2_18_25_i,temp_m2_18_27_r,temp_m2_18_27_i,temp_m2_20_25_r,temp_m2_20_25_i,temp_m2_20_27_r,temp_m2_20_27_i,temp_b2_18_25_r,temp_b2_18_25_i,temp_b2_18_27_r,temp_b2_18_27_i,temp_b2_20_25_r,temp_b2_20_25_i,temp_b2_20_27_r,temp_b2_20_27_i);
MULT MULT412 (clk,temp_b1_18_26_r,temp_b1_18_26_i,temp_b1_18_28_r,temp_b1_18_28_i,temp_b1_20_26_r,temp_b1_20_26_i,temp_b1_20_28_r,temp_b1_20_28_i,temp_m2_18_26_r,temp_m2_18_26_i,temp_m2_18_28_r,temp_m2_18_28_i,temp_m2_20_26_r,temp_m2_20_26_i,temp_m2_20_28_r,temp_m2_20_28_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly412 (clk,temp_m2_18_26_r,temp_m2_18_26_i,temp_m2_18_28_r,temp_m2_18_28_i,temp_m2_20_26_r,temp_m2_20_26_i,temp_m2_20_28_r,temp_m2_20_28_i,temp_b2_18_26_r,temp_b2_18_26_i,temp_b2_18_28_r,temp_b2_18_28_i,temp_b2_20_26_r,temp_b2_20_26_i,temp_b2_20_28_r,temp_b2_20_28_i);
MULT MULT413 (clk,temp_b1_17_29_r,temp_b1_17_29_i,temp_b1_17_31_r,temp_b1_17_31_i,temp_b1_19_29_r,temp_b1_19_29_i,temp_b1_19_31_r,temp_b1_19_31_i,temp_m2_17_29_r,temp_m2_17_29_i,temp_m2_17_31_r,temp_m2_17_31_i,temp_m2_19_29_r,temp_m2_19_29_i,temp_m2_19_31_r,temp_m2_19_31_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly413 (clk,temp_m2_17_29_r,temp_m2_17_29_i,temp_m2_17_31_r,temp_m2_17_31_i,temp_m2_19_29_r,temp_m2_19_29_i,temp_m2_19_31_r,temp_m2_19_31_i,temp_b2_17_29_r,temp_b2_17_29_i,temp_b2_17_31_r,temp_b2_17_31_i,temp_b2_19_29_r,temp_b2_19_29_i,temp_b2_19_31_r,temp_b2_19_31_i);
MULT MULT414 (clk,temp_b1_17_30_r,temp_b1_17_30_i,temp_b1_17_32_r,temp_b1_17_32_i,temp_b1_19_30_r,temp_b1_19_30_i,temp_b1_19_32_r,temp_b1_19_32_i,temp_m2_17_30_r,temp_m2_17_30_i,temp_m2_17_32_r,temp_m2_17_32_i,temp_m2_19_30_r,temp_m2_19_30_i,temp_m2_19_32_r,temp_m2_19_32_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly414 (clk,temp_m2_17_30_r,temp_m2_17_30_i,temp_m2_17_32_r,temp_m2_17_32_i,temp_m2_19_30_r,temp_m2_19_30_i,temp_m2_19_32_r,temp_m2_19_32_i,temp_b2_17_30_r,temp_b2_17_30_i,temp_b2_17_32_r,temp_b2_17_32_i,temp_b2_19_30_r,temp_b2_19_30_i,temp_b2_19_32_r,temp_b2_19_32_i);
MULT MULT415 (clk,temp_b1_18_29_r,temp_b1_18_29_i,temp_b1_18_31_r,temp_b1_18_31_i,temp_b1_20_29_r,temp_b1_20_29_i,temp_b1_20_31_r,temp_b1_20_31_i,temp_m2_18_29_r,temp_m2_18_29_i,temp_m2_18_31_r,temp_m2_18_31_i,temp_m2_20_29_r,temp_m2_20_29_i,temp_m2_20_31_r,temp_m2_20_31_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly415 (clk,temp_m2_18_29_r,temp_m2_18_29_i,temp_m2_18_31_r,temp_m2_18_31_i,temp_m2_20_29_r,temp_m2_20_29_i,temp_m2_20_31_r,temp_m2_20_31_i,temp_b2_18_29_r,temp_b2_18_29_i,temp_b2_18_31_r,temp_b2_18_31_i,temp_b2_20_29_r,temp_b2_20_29_i,temp_b2_20_31_r,temp_b2_20_31_i);
MULT MULT416 (clk,temp_b1_18_30_r,temp_b1_18_30_i,temp_b1_18_32_r,temp_b1_18_32_i,temp_b1_20_30_r,temp_b1_20_30_i,temp_b1_20_32_r,temp_b1_20_32_i,temp_m2_18_30_r,temp_m2_18_30_i,temp_m2_18_32_r,temp_m2_18_32_i,temp_m2_20_30_r,temp_m2_20_30_i,temp_m2_20_32_r,temp_m2_20_32_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly416 (clk,temp_m2_18_30_r,temp_m2_18_30_i,temp_m2_18_32_r,temp_m2_18_32_i,temp_m2_20_30_r,temp_m2_20_30_i,temp_m2_20_32_r,temp_m2_20_32_i,temp_b2_18_30_r,temp_b2_18_30_i,temp_b2_18_32_r,temp_b2_18_32_i,temp_b2_20_30_r,temp_b2_20_30_i,temp_b2_20_32_r,temp_b2_20_32_i);
MULT MULT417 (clk,temp_b1_21_1_r,temp_b1_21_1_i,temp_b1_21_3_r,temp_b1_21_3_i,temp_b1_23_1_r,temp_b1_23_1_i,temp_b1_23_3_r,temp_b1_23_3_i,temp_m2_21_1_r,temp_m2_21_1_i,temp_m2_21_3_r,temp_m2_21_3_i,temp_m2_23_1_r,temp_m2_23_1_i,temp_m2_23_3_r,temp_m2_23_3_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly417 (clk,temp_m2_21_1_r,temp_m2_21_1_i,temp_m2_21_3_r,temp_m2_21_3_i,temp_m2_23_1_r,temp_m2_23_1_i,temp_m2_23_3_r,temp_m2_23_3_i,temp_b2_21_1_r,temp_b2_21_1_i,temp_b2_21_3_r,temp_b2_21_3_i,temp_b2_23_1_r,temp_b2_23_1_i,temp_b2_23_3_r,temp_b2_23_3_i);
MULT MULT418 (clk,temp_b1_21_2_r,temp_b1_21_2_i,temp_b1_21_4_r,temp_b1_21_4_i,temp_b1_23_2_r,temp_b1_23_2_i,temp_b1_23_4_r,temp_b1_23_4_i,temp_m2_21_2_r,temp_m2_21_2_i,temp_m2_21_4_r,temp_m2_21_4_i,temp_m2_23_2_r,temp_m2_23_2_i,temp_m2_23_4_r,temp_m2_23_4_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly418 (clk,temp_m2_21_2_r,temp_m2_21_2_i,temp_m2_21_4_r,temp_m2_21_4_i,temp_m2_23_2_r,temp_m2_23_2_i,temp_m2_23_4_r,temp_m2_23_4_i,temp_b2_21_2_r,temp_b2_21_2_i,temp_b2_21_4_r,temp_b2_21_4_i,temp_b2_23_2_r,temp_b2_23_2_i,temp_b2_23_4_r,temp_b2_23_4_i);
MULT MULT419 (clk,temp_b1_22_1_r,temp_b1_22_1_i,temp_b1_22_3_r,temp_b1_22_3_i,temp_b1_24_1_r,temp_b1_24_1_i,temp_b1_24_3_r,temp_b1_24_3_i,temp_m2_22_1_r,temp_m2_22_1_i,temp_m2_22_3_r,temp_m2_22_3_i,temp_m2_24_1_r,temp_m2_24_1_i,temp_m2_24_3_r,temp_m2_24_3_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly419 (clk,temp_m2_22_1_r,temp_m2_22_1_i,temp_m2_22_3_r,temp_m2_22_3_i,temp_m2_24_1_r,temp_m2_24_1_i,temp_m2_24_3_r,temp_m2_24_3_i,temp_b2_22_1_r,temp_b2_22_1_i,temp_b2_22_3_r,temp_b2_22_3_i,temp_b2_24_1_r,temp_b2_24_1_i,temp_b2_24_3_r,temp_b2_24_3_i);
MULT MULT420 (clk,temp_b1_22_2_r,temp_b1_22_2_i,temp_b1_22_4_r,temp_b1_22_4_i,temp_b1_24_2_r,temp_b1_24_2_i,temp_b1_24_4_r,temp_b1_24_4_i,temp_m2_22_2_r,temp_m2_22_2_i,temp_m2_22_4_r,temp_m2_22_4_i,temp_m2_24_2_r,temp_m2_24_2_i,temp_m2_24_4_r,temp_m2_24_4_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly420 (clk,temp_m2_22_2_r,temp_m2_22_2_i,temp_m2_22_4_r,temp_m2_22_4_i,temp_m2_24_2_r,temp_m2_24_2_i,temp_m2_24_4_r,temp_m2_24_4_i,temp_b2_22_2_r,temp_b2_22_2_i,temp_b2_22_4_r,temp_b2_22_4_i,temp_b2_24_2_r,temp_b2_24_2_i,temp_b2_24_4_r,temp_b2_24_4_i);
MULT MULT421 (clk,temp_b1_21_5_r,temp_b1_21_5_i,temp_b1_21_7_r,temp_b1_21_7_i,temp_b1_23_5_r,temp_b1_23_5_i,temp_b1_23_7_r,temp_b1_23_7_i,temp_m2_21_5_r,temp_m2_21_5_i,temp_m2_21_7_r,temp_m2_21_7_i,temp_m2_23_5_r,temp_m2_23_5_i,temp_m2_23_7_r,temp_m2_23_7_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly421 (clk,temp_m2_21_5_r,temp_m2_21_5_i,temp_m2_21_7_r,temp_m2_21_7_i,temp_m2_23_5_r,temp_m2_23_5_i,temp_m2_23_7_r,temp_m2_23_7_i,temp_b2_21_5_r,temp_b2_21_5_i,temp_b2_21_7_r,temp_b2_21_7_i,temp_b2_23_5_r,temp_b2_23_5_i,temp_b2_23_7_r,temp_b2_23_7_i);
MULT MULT422 (clk,temp_b1_21_6_r,temp_b1_21_6_i,temp_b1_21_8_r,temp_b1_21_8_i,temp_b1_23_6_r,temp_b1_23_6_i,temp_b1_23_8_r,temp_b1_23_8_i,temp_m2_21_6_r,temp_m2_21_6_i,temp_m2_21_8_r,temp_m2_21_8_i,temp_m2_23_6_r,temp_m2_23_6_i,temp_m2_23_8_r,temp_m2_23_8_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly422 (clk,temp_m2_21_6_r,temp_m2_21_6_i,temp_m2_21_8_r,temp_m2_21_8_i,temp_m2_23_6_r,temp_m2_23_6_i,temp_m2_23_8_r,temp_m2_23_8_i,temp_b2_21_6_r,temp_b2_21_6_i,temp_b2_21_8_r,temp_b2_21_8_i,temp_b2_23_6_r,temp_b2_23_6_i,temp_b2_23_8_r,temp_b2_23_8_i);
MULT MULT423 (clk,temp_b1_22_5_r,temp_b1_22_5_i,temp_b1_22_7_r,temp_b1_22_7_i,temp_b1_24_5_r,temp_b1_24_5_i,temp_b1_24_7_r,temp_b1_24_7_i,temp_m2_22_5_r,temp_m2_22_5_i,temp_m2_22_7_r,temp_m2_22_7_i,temp_m2_24_5_r,temp_m2_24_5_i,temp_m2_24_7_r,temp_m2_24_7_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly423 (clk,temp_m2_22_5_r,temp_m2_22_5_i,temp_m2_22_7_r,temp_m2_22_7_i,temp_m2_24_5_r,temp_m2_24_5_i,temp_m2_24_7_r,temp_m2_24_7_i,temp_b2_22_5_r,temp_b2_22_5_i,temp_b2_22_7_r,temp_b2_22_7_i,temp_b2_24_5_r,temp_b2_24_5_i,temp_b2_24_7_r,temp_b2_24_7_i);
MULT MULT424 (clk,temp_b1_22_6_r,temp_b1_22_6_i,temp_b1_22_8_r,temp_b1_22_8_i,temp_b1_24_6_r,temp_b1_24_6_i,temp_b1_24_8_r,temp_b1_24_8_i,temp_m2_22_6_r,temp_m2_22_6_i,temp_m2_22_8_r,temp_m2_22_8_i,temp_m2_24_6_r,temp_m2_24_6_i,temp_m2_24_8_r,temp_m2_24_8_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly424 (clk,temp_m2_22_6_r,temp_m2_22_6_i,temp_m2_22_8_r,temp_m2_22_8_i,temp_m2_24_6_r,temp_m2_24_6_i,temp_m2_24_8_r,temp_m2_24_8_i,temp_b2_22_6_r,temp_b2_22_6_i,temp_b2_22_8_r,temp_b2_22_8_i,temp_b2_24_6_r,temp_b2_24_6_i,temp_b2_24_8_r,temp_b2_24_8_i);
MULT MULT425 (clk,temp_b1_21_9_r,temp_b1_21_9_i,temp_b1_21_11_r,temp_b1_21_11_i,temp_b1_23_9_r,temp_b1_23_9_i,temp_b1_23_11_r,temp_b1_23_11_i,temp_m2_21_9_r,temp_m2_21_9_i,temp_m2_21_11_r,temp_m2_21_11_i,temp_m2_23_9_r,temp_m2_23_9_i,temp_m2_23_11_r,temp_m2_23_11_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly425 (clk,temp_m2_21_9_r,temp_m2_21_9_i,temp_m2_21_11_r,temp_m2_21_11_i,temp_m2_23_9_r,temp_m2_23_9_i,temp_m2_23_11_r,temp_m2_23_11_i,temp_b2_21_9_r,temp_b2_21_9_i,temp_b2_21_11_r,temp_b2_21_11_i,temp_b2_23_9_r,temp_b2_23_9_i,temp_b2_23_11_r,temp_b2_23_11_i);
MULT MULT426 (clk,temp_b1_21_10_r,temp_b1_21_10_i,temp_b1_21_12_r,temp_b1_21_12_i,temp_b1_23_10_r,temp_b1_23_10_i,temp_b1_23_12_r,temp_b1_23_12_i,temp_m2_21_10_r,temp_m2_21_10_i,temp_m2_21_12_r,temp_m2_21_12_i,temp_m2_23_10_r,temp_m2_23_10_i,temp_m2_23_12_r,temp_m2_23_12_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly426 (clk,temp_m2_21_10_r,temp_m2_21_10_i,temp_m2_21_12_r,temp_m2_21_12_i,temp_m2_23_10_r,temp_m2_23_10_i,temp_m2_23_12_r,temp_m2_23_12_i,temp_b2_21_10_r,temp_b2_21_10_i,temp_b2_21_12_r,temp_b2_21_12_i,temp_b2_23_10_r,temp_b2_23_10_i,temp_b2_23_12_r,temp_b2_23_12_i);
MULT MULT427 (clk,temp_b1_22_9_r,temp_b1_22_9_i,temp_b1_22_11_r,temp_b1_22_11_i,temp_b1_24_9_r,temp_b1_24_9_i,temp_b1_24_11_r,temp_b1_24_11_i,temp_m2_22_9_r,temp_m2_22_9_i,temp_m2_22_11_r,temp_m2_22_11_i,temp_m2_24_9_r,temp_m2_24_9_i,temp_m2_24_11_r,temp_m2_24_11_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly427 (clk,temp_m2_22_9_r,temp_m2_22_9_i,temp_m2_22_11_r,temp_m2_22_11_i,temp_m2_24_9_r,temp_m2_24_9_i,temp_m2_24_11_r,temp_m2_24_11_i,temp_b2_22_9_r,temp_b2_22_9_i,temp_b2_22_11_r,temp_b2_22_11_i,temp_b2_24_9_r,temp_b2_24_9_i,temp_b2_24_11_r,temp_b2_24_11_i);
MULT MULT428 (clk,temp_b1_22_10_r,temp_b1_22_10_i,temp_b1_22_12_r,temp_b1_22_12_i,temp_b1_24_10_r,temp_b1_24_10_i,temp_b1_24_12_r,temp_b1_24_12_i,temp_m2_22_10_r,temp_m2_22_10_i,temp_m2_22_12_r,temp_m2_22_12_i,temp_m2_24_10_r,temp_m2_24_10_i,temp_m2_24_12_r,temp_m2_24_12_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly428 (clk,temp_m2_22_10_r,temp_m2_22_10_i,temp_m2_22_12_r,temp_m2_22_12_i,temp_m2_24_10_r,temp_m2_24_10_i,temp_m2_24_12_r,temp_m2_24_12_i,temp_b2_22_10_r,temp_b2_22_10_i,temp_b2_22_12_r,temp_b2_22_12_i,temp_b2_24_10_r,temp_b2_24_10_i,temp_b2_24_12_r,temp_b2_24_12_i);
MULT MULT429 (clk,temp_b1_21_13_r,temp_b1_21_13_i,temp_b1_21_15_r,temp_b1_21_15_i,temp_b1_23_13_r,temp_b1_23_13_i,temp_b1_23_15_r,temp_b1_23_15_i,temp_m2_21_13_r,temp_m2_21_13_i,temp_m2_21_15_r,temp_m2_21_15_i,temp_m2_23_13_r,temp_m2_23_13_i,temp_m2_23_15_r,temp_m2_23_15_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly429 (clk,temp_m2_21_13_r,temp_m2_21_13_i,temp_m2_21_15_r,temp_m2_21_15_i,temp_m2_23_13_r,temp_m2_23_13_i,temp_m2_23_15_r,temp_m2_23_15_i,temp_b2_21_13_r,temp_b2_21_13_i,temp_b2_21_15_r,temp_b2_21_15_i,temp_b2_23_13_r,temp_b2_23_13_i,temp_b2_23_15_r,temp_b2_23_15_i);
MULT MULT430 (clk,temp_b1_21_14_r,temp_b1_21_14_i,temp_b1_21_16_r,temp_b1_21_16_i,temp_b1_23_14_r,temp_b1_23_14_i,temp_b1_23_16_r,temp_b1_23_16_i,temp_m2_21_14_r,temp_m2_21_14_i,temp_m2_21_16_r,temp_m2_21_16_i,temp_m2_23_14_r,temp_m2_23_14_i,temp_m2_23_16_r,temp_m2_23_16_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly430 (clk,temp_m2_21_14_r,temp_m2_21_14_i,temp_m2_21_16_r,temp_m2_21_16_i,temp_m2_23_14_r,temp_m2_23_14_i,temp_m2_23_16_r,temp_m2_23_16_i,temp_b2_21_14_r,temp_b2_21_14_i,temp_b2_21_16_r,temp_b2_21_16_i,temp_b2_23_14_r,temp_b2_23_14_i,temp_b2_23_16_r,temp_b2_23_16_i);
MULT MULT431 (clk,temp_b1_22_13_r,temp_b1_22_13_i,temp_b1_22_15_r,temp_b1_22_15_i,temp_b1_24_13_r,temp_b1_24_13_i,temp_b1_24_15_r,temp_b1_24_15_i,temp_m2_22_13_r,temp_m2_22_13_i,temp_m2_22_15_r,temp_m2_22_15_i,temp_m2_24_13_r,temp_m2_24_13_i,temp_m2_24_15_r,temp_m2_24_15_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly431 (clk,temp_m2_22_13_r,temp_m2_22_13_i,temp_m2_22_15_r,temp_m2_22_15_i,temp_m2_24_13_r,temp_m2_24_13_i,temp_m2_24_15_r,temp_m2_24_15_i,temp_b2_22_13_r,temp_b2_22_13_i,temp_b2_22_15_r,temp_b2_22_15_i,temp_b2_24_13_r,temp_b2_24_13_i,temp_b2_24_15_r,temp_b2_24_15_i);
MULT MULT432 (clk,temp_b1_22_14_r,temp_b1_22_14_i,temp_b1_22_16_r,temp_b1_22_16_i,temp_b1_24_14_r,temp_b1_24_14_i,temp_b1_24_16_r,temp_b1_24_16_i,temp_m2_22_14_r,temp_m2_22_14_i,temp_m2_22_16_r,temp_m2_22_16_i,temp_m2_24_14_r,temp_m2_24_14_i,temp_m2_24_16_r,temp_m2_24_16_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly432 (clk,temp_m2_22_14_r,temp_m2_22_14_i,temp_m2_22_16_r,temp_m2_22_16_i,temp_m2_24_14_r,temp_m2_24_14_i,temp_m2_24_16_r,temp_m2_24_16_i,temp_b2_22_14_r,temp_b2_22_14_i,temp_b2_22_16_r,temp_b2_22_16_i,temp_b2_24_14_r,temp_b2_24_14_i,temp_b2_24_16_r,temp_b2_24_16_i);
MULT MULT433 (clk,temp_b1_21_17_r,temp_b1_21_17_i,temp_b1_21_19_r,temp_b1_21_19_i,temp_b1_23_17_r,temp_b1_23_17_i,temp_b1_23_19_r,temp_b1_23_19_i,temp_m2_21_17_r,temp_m2_21_17_i,temp_m2_21_19_r,temp_m2_21_19_i,temp_m2_23_17_r,temp_m2_23_17_i,temp_m2_23_19_r,temp_m2_23_19_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly433 (clk,temp_m2_21_17_r,temp_m2_21_17_i,temp_m2_21_19_r,temp_m2_21_19_i,temp_m2_23_17_r,temp_m2_23_17_i,temp_m2_23_19_r,temp_m2_23_19_i,temp_b2_21_17_r,temp_b2_21_17_i,temp_b2_21_19_r,temp_b2_21_19_i,temp_b2_23_17_r,temp_b2_23_17_i,temp_b2_23_19_r,temp_b2_23_19_i);
MULT MULT434 (clk,temp_b1_21_18_r,temp_b1_21_18_i,temp_b1_21_20_r,temp_b1_21_20_i,temp_b1_23_18_r,temp_b1_23_18_i,temp_b1_23_20_r,temp_b1_23_20_i,temp_m2_21_18_r,temp_m2_21_18_i,temp_m2_21_20_r,temp_m2_21_20_i,temp_m2_23_18_r,temp_m2_23_18_i,temp_m2_23_20_r,temp_m2_23_20_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly434 (clk,temp_m2_21_18_r,temp_m2_21_18_i,temp_m2_21_20_r,temp_m2_21_20_i,temp_m2_23_18_r,temp_m2_23_18_i,temp_m2_23_20_r,temp_m2_23_20_i,temp_b2_21_18_r,temp_b2_21_18_i,temp_b2_21_20_r,temp_b2_21_20_i,temp_b2_23_18_r,temp_b2_23_18_i,temp_b2_23_20_r,temp_b2_23_20_i);
MULT MULT435 (clk,temp_b1_22_17_r,temp_b1_22_17_i,temp_b1_22_19_r,temp_b1_22_19_i,temp_b1_24_17_r,temp_b1_24_17_i,temp_b1_24_19_r,temp_b1_24_19_i,temp_m2_22_17_r,temp_m2_22_17_i,temp_m2_22_19_r,temp_m2_22_19_i,temp_m2_24_17_r,temp_m2_24_17_i,temp_m2_24_19_r,temp_m2_24_19_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly435 (clk,temp_m2_22_17_r,temp_m2_22_17_i,temp_m2_22_19_r,temp_m2_22_19_i,temp_m2_24_17_r,temp_m2_24_17_i,temp_m2_24_19_r,temp_m2_24_19_i,temp_b2_22_17_r,temp_b2_22_17_i,temp_b2_22_19_r,temp_b2_22_19_i,temp_b2_24_17_r,temp_b2_24_17_i,temp_b2_24_19_r,temp_b2_24_19_i);
MULT MULT436 (clk,temp_b1_22_18_r,temp_b1_22_18_i,temp_b1_22_20_r,temp_b1_22_20_i,temp_b1_24_18_r,temp_b1_24_18_i,temp_b1_24_20_r,temp_b1_24_20_i,temp_m2_22_18_r,temp_m2_22_18_i,temp_m2_22_20_r,temp_m2_22_20_i,temp_m2_24_18_r,temp_m2_24_18_i,temp_m2_24_20_r,temp_m2_24_20_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly436 (clk,temp_m2_22_18_r,temp_m2_22_18_i,temp_m2_22_20_r,temp_m2_22_20_i,temp_m2_24_18_r,temp_m2_24_18_i,temp_m2_24_20_r,temp_m2_24_20_i,temp_b2_22_18_r,temp_b2_22_18_i,temp_b2_22_20_r,temp_b2_22_20_i,temp_b2_24_18_r,temp_b2_24_18_i,temp_b2_24_20_r,temp_b2_24_20_i);
MULT MULT437 (clk,temp_b1_21_21_r,temp_b1_21_21_i,temp_b1_21_23_r,temp_b1_21_23_i,temp_b1_23_21_r,temp_b1_23_21_i,temp_b1_23_23_r,temp_b1_23_23_i,temp_m2_21_21_r,temp_m2_21_21_i,temp_m2_21_23_r,temp_m2_21_23_i,temp_m2_23_21_r,temp_m2_23_21_i,temp_m2_23_23_r,temp_m2_23_23_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly437 (clk,temp_m2_21_21_r,temp_m2_21_21_i,temp_m2_21_23_r,temp_m2_21_23_i,temp_m2_23_21_r,temp_m2_23_21_i,temp_m2_23_23_r,temp_m2_23_23_i,temp_b2_21_21_r,temp_b2_21_21_i,temp_b2_21_23_r,temp_b2_21_23_i,temp_b2_23_21_r,temp_b2_23_21_i,temp_b2_23_23_r,temp_b2_23_23_i);
MULT MULT438 (clk,temp_b1_21_22_r,temp_b1_21_22_i,temp_b1_21_24_r,temp_b1_21_24_i,temp_b1_23_22_r,temp_b1_23_22_i,temp_b1_23_24_r,temp_b1_23_24_i,temp_m2_21_22_r,temp_m2_21_22_i,temp_m2_21_24_r,temp_m2_21_24_i,temp_m2_23_22_r,temp_m2_23_22_i,temp_m2_23_24_r,temp_m2_23_24_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly438 (clk,temp_m2_21_22_r,temp_m2_21_22_i,temp_m2_21_24_r,temp_m2_21_24_i,temp_m2_23_22_r,temp_m2_23_22_i,temp_m2_23_24_r,temp_m2_23_24_i,temp_b2_21_22_r,temp_b2_21_22_i,temp_b2_21_24_r,temp_b2_21_24_i,temp_b2_23_22_r,temp_b2_23_22_i,temp_b2_23_24_r,temp_b2_23_24_i);
MULT MULT439 (clk,temp_b1_22_21_r,temp_b1_22_21_i,temp_b1_22_23_r,temp_b1_22_23_i,temp_b1_24_21_r,temp_b1_24_21_i,temp_b1_24_23_r,temp_b1_24_23_i,temp_m2_22_21_r,temp_m2_22_21_i,temp_m2_22_23_r,temp_m2_22_23_i,temp_m2_24_21_r,temp_m2_24_21_i,temp_m2_24_23_r,temp_m2_24_23_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly439 (clk,temp_m2_22_21_r,temp_m2_22_21_i,temp_m2_22_23_r,temp_m2_22_23_i,temp_m2_24_21_r,temp_m2_24_21_i,temp_m2_24_23_r,temp_m2_24_23_i,temp_b2_22_21_r,temp_b2_22_21_i,temp_b2_22_23_r,temp_b2_22_23_i,temp_b2_24_21_r,temp_b2_24_21_i,temp_b2_24_23_r,temp_b2_24_23_i);
MULT MULT440 (clk,temp_b1_22_22_r,temp_b1_22_22_i,temp_b1_22_24_r,temp_b1_22_24_i,temp_b1_24_22_r,temp_b1_24_22_i,temp_b1_24_24_r,temp_b1_24_24_i,temp_m2_22_22_r,temp_m2_22_22_i,temp_m2_22_24_r,temp_m2_22_24_i,temp_m2_24_22_r,temp_m2_24_22_i,temp_m2_24_24_r,temp_m2_24_24_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly440 (clk,temp_m2_22_22_r,temp_m2_22_22_i,temp_m2_22_24_r,temp_m2_22_24_i,temp_m2_24_22_r,temp_m2_24_22_i,temp_m2_24_24_r,temp_m2_24_24_i,temp_b2_22_22_r,temp_b2_22_22_i,temp_b2_22_24_r,temp_b2_22_24_i,temp_b2_24_22_r,temp_b2_24_22_i,temp_b2_24_24_r,temp_b2_24_24_i);
MULT MULT441 (clk,temp_b1_21_25_r,temp_b1_21_25_i,temp_b1_21_27_r,temp_b1_21_27_i,temp_b1_23_25_r,temp_b1_23_25_i,temp_b1_23_27_r,temp_b1_23_27_i,temp_m2_21_25_r,temp_m2_21_25_i,temp_m2_21_27_r,temp_m2_21_27_i,temp_m2_23_25_r,temp_m2_23_25_i,temp_m2_23_27_r,temp_m2_23_27_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly441 (clk,temp_m2_21_25_r,temp_m2_21_25_i,temp_m2_21_27_r,temp_m2_21_27_i,temp_m2_23_25_r,temp_m2_23_25_i,temp_m2_23_27_r,temp_m2_23_27_i,temp_b2_21_25_r,temp_b2_21_25_i,temp_b2_21_27_r,temp_b2_21_27_i,temp_b2_23_25_r,temp_b2_23_25_i,temp_b2_23_27_r,temp_b2_23_27_i);
MULT MULT442 (clk,temp_b1_21_26_r,temp_b1_21_26_i,temp_b1_21_28_r,temp_b1_21_28_i,temp_b1_23_26_r,temp_b1_23_26_i,temp_b1_23_28_r,temp_b1_23_28_i,temp_m2_21_26_r,temp_m2_21_26_i,temp_m2_21_28_r,temp_m2_21_28_i,temp_m2_23_26_r,temp_m2_23_26_i,temp_m2_23_28_r,temp_m2_23_28_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly442 (clk,temp_m2_21_26_r,temp_m2_21_26_i,temp_m2_21_28_r,temp_m2_21_28_i,temp_m2_23_26_r,temp_m2_23_26_i,temp_m2_23_28_r,temp_m2_23_28_i,temp_b2_21_26_r,temp_b2_21_26_i,temp_b2_21_28_r,temp_b2_21_28_i,temp_b2_23_26_r,temp_b2_23_26_i,temp_b2_23_28_r,temp_b2_23_28_i);
MULT MULT443 (clk,temp_b1_22_25_r,temp_b1_22_25_i,temp_b1_22_27_r,temp_b1_22_27_i,temp_b1_24_25_r,temp_b1_24_25_i,temp_b1_24_27_r,temp_b1_24_27_i,temp_m2_22_25_r,temp_m2_22_25_i,temp_m2_22_27_r,temp_m2_22_27_i,temp_m2_24_25_r,temp_m2_24_25_i,temp_m2_24_27_r,temp_m2_24_27_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly443 (clk,temp_m2_22_25_r,temp_m2_22_25_i,temp_m2_22_27_r,temp_m2_22_27_i,temp_m2_24_25_r,temp_m2_24_25_i,temp_m2_24_27_r,temp_m2_24_27_i,temp_b2_22_25_r,temp_b2_22_25_i,temp_b2_22_27_r,temp_b2_22_27_i,temp_b2_24_25_r,temp_b2_24_25_i,temp_b2_24_27_r,temp_b2_24_27_i);
MULT MULT444 (clk,temp_b1_22_26_r,temp_b1_22_26_i,temp_b1_22_28_r,temp_b1_22_28_i,temp_b1_24_26_r,temp_b1_24_26_i,temp_b1_24_28_r,temp_b1_24_28_i,temp_m2_22_26_r,temp_m2_22_26_i,temp_m2_22_28_r,temp_m2_22_28_i,temp_m2_24_26_r,temp_m2_24_26_i,temp_m2_24_28_r,temp_m2_24_28_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly444 (clk,temp_m2_22_26_r,temp_m2_22_26_i,temp_m2_22_28_r,temp_m2_22_28_i,temp_m2_24_26_r,temp_m2_24_26_i,temp_m2_24_28_r,temp_m2_24_28_i,temp_b2_22_26_r,temp_b2_22_26_i,temp_b2_22_28_r,temp_b2_22_28_i,temp_b2_24_26_r,temp_b2_24_26_i,temp_b2_24_28_r,temp_b2_24_28_i);
MULT MULT445 (clk,temp_b1_21_29_r,temp_b1_21_29_i,temp_b1_21_31_r,temp_b1_21_31_i,temp_b1_23_29_r,temp_b1_23_29_i,temp_b1_23_31_r,temp_b1_23_31_i,temp_m2_21_29_r,temp_m2_21_29_i,temp_m2_21_31_r,temp_m2_21_31_i,temp_m2_23_29_r,temp_m2_23_29_i,temp_m2_23_31_r,temp_m2_23_31_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly445 (clk,temp_m2_21_29_r,temp_m2_21_29_i,temp_m2_21_31_r,temp_m2_21_31_i,temp_m2_23_29_r,temp_m2_23_29_i,temp_m2_23_31_r,temp_m2_23_31_i,temp_b2_21_29_r,temp_b2_21_29_i,temp_b2_21_31_r,temp_b2_21_31_i,temp_b2_23_29_r,temp_b2_23_29_i,temp_b2_23_31_r,temp_b2_23_31_i);
MULT MULT446 (clk,temp_b1_21_30_r,temp_b1_21_30_i,temp_b1_21_32_r,temp_b1_21_32_i,temp_b1_23_30_r,temp_b1_23_30_i,temp_b1_23_32_r,temp_b1_23_32_i,temp_m2_21_30_r,temp_m2_21_30_i,temp_m2_21_32_r,temp_m2_21_32_i,temp_m2_23_30_r,temp_m2_23_30_i,temp_m2_23_32_r,temp_m2_23_32_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly446 (clk,temp_m2_21_30_r,temp_m2_21_30_i,temp_m2_21_32_r,temp_m2_21_32_i,temp_m2_23_30_r,temp_m2_23_30_i,temp_m2_23_32_r,temp_m2_23_32_i,temp_b2_21_30_r,temp_b2_21_30_i,temp_b2_21_32_r,temp_b2_21_32_i,temp_b2_23_30_r,temp_b2_23_30_i,temp_b2_23_32_r,temp_b2_23_32_i);
MULT MULT447 (clk,temp_b1_22_29_r,temp_b1_22_29_i,temp_b1_22_31_r,temp_b1_22_31_i,temp_b1_24_29_r,temp_b1_24_29_i,temp_b1_24_31_r,temp_b1_24_31_i,temp_m2_22_29_r,temp_m2_22_29_i,temp_m2_22_31_r,temp_m2_22_31_i,temp_m2_24_29_r,temp_m2_24_29_i,temp_m2_24_31_r,temp_m2_24_31_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly447 (clk,temp_m2_22_29_r,temp_m2_22_29_i,temp_m2_22_31_r,temp_m2_22_31_i,temp_m2_24_29_r,temp_m2_24_29_i,temp_m2_24_31_r,temp_m2_24_31_i,temp_b2_22_29_r,temp_b2_22_29_i,temp_b2_22_31_r,temp_b2_22_31_i,temp_b2_24_29_r,temp_b2_24_29_i,temp_b2_24_31_r,temp_b2_24_31_i);
MULT MULT448 (clk,temp_b1_22_30_r,temp_b1_22_30_i,temp_b1_22_32_r,temp_b1_22_32_i,temp_b1_24_30_r,temp_b1_24_30_i,temp_b1_24_32_r,temp_b1_24_32_i,temp_m2_22_30_r,temp_m2_22_30_i,temp_m2_22_32_r,temp_m2_22_32_i,temp_m2_24_30_r,temp_m2_24_30_i,temp_m2_24_32_r,temp_m2_24_32_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly448 (clk,temp_m2_22_30_r,temp_m2_22_30_i,temp_m2_22_32_r,temp_m2_22_32_i,temp_m2_24_30_r,temp_m2_24_30_i,temp_m2_24_32_r,temp_m2_24_32_i,temp_b2_22_30_r,temp_b2_22_30_i,temp_b2_22_32_r,temp_b2_22_32_i,temp_b2_24_30_r,temp_b2_24_30_i,temp_b2_24_32_r,temp_b2_24_32_i);
MULT MULT449 (clk,temp_b1_25_1_r,temp_b1_25_1_i,temp_b1_25_3_r,temp_b1_25_3_i,temp_b1_27_1_r,temp_b1_27_1_i,temp_b1_27_3_r,temp_b1_27_3_i,temp_m2_25_1_r,temp_m2_25_1_i,temp_m2_25_3_r,temp_m2_25_3_i,temp_m2_27_1_r,temp_m2_27_1_i,temp_m2_27_3_r,temp_m2_27_3_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly449 (clk,temp_m2_25_1_r,temp_m2_25_1_i,temp_m2_25_3_r,temp_m2_25_3_i,temp_m2_27_1_r,temp_m2_27_1_i,temp_m2_27_3_r,temp_m2_27_3_i,temp_b2_25_1_r,temp_b2_25_1_i,temp_b2_25_3_r,temp_b2_25_3_i,temp_b2_27_1_r,temp_b2_27_1_i,temp_b2_27_3_r,temp_b2_27_3_i);
MULT MULT450 (clk,temp_b1_25_2_r,temp_b1_25_2_i,temp_b1_25_4_r,temp_b1_25_4_i,temp_b1_27_2_r,temp_b1_27_2_i,temp_b1_27_4_r,temp_b1_27_4_i,temp_m2_25_2_r,temp_m2_25_2_i,temp_m2_25_4_r,temp_m2_25_4_i,temp_m2_27_2_r,temp_m2_27_2_i,temp_m2_27_4_r,temp_m2_27_4_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly450 (clk,temp_m2_25_2_r,temp_m2_25_2_i,temp_m2_25_4_r,temp_m2_25_4_i,temp_m2_27_2_r,temp_m2_27_2_i,temp_m2_27_4_r,temp_m2_27_4_i,temp_b2_25_2_r,temp_b2_25_2_i,temp_b2_25_4_r,temp_b2_25_4_i,temp_b2_27_2_r,temp_b2_27_2_i,temp_b2_27_4_r,temp_b2_27_4_i);
MULT MULT451 (clk,temp_b1_26_1_r,temp_b1_26_1_i,temp_b1_26_3_r,temp_b1_26_3_i,temp_b1_28_1_r,temp_b1_28_1_i,temp_b1_28_3_r,temp_b1_28_3_i,temp_m2_26_1_r,temp_m2_26_1_i,temp_m2_26_3_r,temp_m2_26_3_i,temp_m2_28_1_r,temp_m2_28_1_i,temp_m2_28_3_r,temp_m2_28_3_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly451 (clk,temp_m2_26_1_r,temp_m2_26_1_i,temp_m2_26_3_r,temp_m2_26_3_i,temp_m2_28_1_r,temp_m2_28_1_i,temp_m2_28_3_r,temp_m2_28_3_i,temp_b2_26_1_r,temp_b2_26_1_i,temp_b2_26_3_r,temp_b2_26_3_i,temp_b2_28_1_r,temp_b2_28_1_i,temp_b2_28_3_r,temp_b2_28_3_i);
MULT MULT452 (clk,temp_b1_26_2_r,temp_b1_26_2_i,temp_b1_26_4_r,temp_b1_26_4_i,temp_b1_28_2_r,temp_b1_28_2_i,temp_b1_28_4_r,temp_b1_28_4_i,temp_m2_26_2_r,temp_m2_26_2_i,temp_m2_26_4_r,temp_m2_26_4_i,temp_m2_28_2_r,temp_m2_28_2_i,temp_m2_28_4_r,temp_m2_28_4_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly452 (clk,temp_m2_26_2_r,temp_m2_26_2_i,temp_m2_26_4_r,temp_m2_26_4_i,temp_m2_28_2_r,temp_m2_28_2_i,temp_m2_28_4_r,temp_m2_28_4_i,temp_b2_26_2_r,temp_b2_26_2_i,temp_b2_26_4_r,temp_b2_26_4_i,temp_b2_28_2_r,temp_b2_28_2_i,temp_b2_28_4_r,temp_b2_28_4_i);
MULT MULT453 (clk,temp_b1_25_5_r,temp_b1_25_5_i,temp_b1_25_7_r,temp_b1_25_7_i,temp_b1_27_5_r,temp_b1_27_5_i,temp_b1_27_7_r,temp_b1_27_7_i,temp_m2_25_5_r,temp_m2_25_5_i,temp_m2_25_7_r,temp_m2_25_7_i,temp_m2_27_5_r,temp_m2_27_5_i,temp_m2_27_7_r,temp_m2_27_7_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly453 (clk,temp_m2_25_5_r,temp_m2_25_5_i,temp_m2_25_7_r,temp_m2_25_7_i,temp_m2_27_5_r,temp_m2_27_5_i,temp_m2_27_7_r,temp_m2_27_7_i,temp_b2_25_5_r,temp_b2_25_5_i,temp_b2_25_7_r,temp_b2_25_7_i,temp_b2_27_5_r,temp_b2_27_5_i,temp_b2_27_7_r,temp_b2_27_7_i);
MULT MULT454 (clk,temp_b1_25_6_r,temp_b1_25_6_i,temp_b1_25_8_r,temp_b1_25_8_i,temp_b1_27_6_r,temp_b1_27_6_i,temp_b1_27_8_r,temp_b1_27_8_i,temp_m2_25_6_r,temp_m2_25_6_i,temp_m2_25_8_r,temp_m2_25_8_i,temp_m2_27_6_r,temp_m2_27_6_i,temp_m2_27_8_r,temp_m2_27_8_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly454 (clk,temp_m2_25_6_r,temp_m2_25_6_i,temp_m2_25_8_r,temp_m2_25_8_i,temp_m2_27_6_r,temp_m2_27_6_i,temp_m2_27_8_r,temp_m2_27_8_i,temp_b2_25_6_r,temp_b2_25_6_i,temp_b2_25_8_r,temp_b2_25_8_i,temp_b2_27_6_r,temp_b2_27_6_i,temp_b2_27_8_r,temp_b2_27_8_i);
MULT MULT455 (clk,temp_b1_26_5_r,temp_b1_26_5_i,temp_b1_26_7_r,temp_b1_26_7_i,temp_b1_28_5_r,temp_b1_28_5_i,temp_b1_28_7_r,temp_b1_28_7_i,temp_m2_26_5_r,temp_m2_26_5_i,temp_m2_26_7_r,temp_m2_26_7_i,temp_m2_28_5_r,temp_m2_28_5_i,temp_m2_28_7_r,temp_m2_28_7_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly455 (clk,temp_m2_26_5_r,temp_m2_26_5_i,temp_m2_26_7_r,temp_m2_26_7_i,temp_m2_28_5_r,temp_m2_28_5_i,temp_m2_28_7_r,temp_m2_28_7_i,temp_b2_26_5_r,temp_b2_26_5_i,temp_b2_26_7_r,temp_b2_26_7_i,temp_b2_28_5_r,temp_b2_28_5_i,temp_b2_28_7_r,temp_b2_28_7_i);
MULT MULT456 (clk,temp_b1_26_6_r,temp_b1_26_6_i,temp_b1_26_8_r,temp_b1_26_8_i,temp_b1_28_6_r,temp_b1_28_6_i,temp_b1_28_8_r,temp_b1_28_8_i,temp_m2_26_6_r,temp_m2_26_6_i,temp_m2_26_8_r,temp_m2_26_8_i,temp_m2_28_6_r,temp_m2_28_6_i,temp_m2_28_8_r,temp_m2_28_8_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly456 (clk,temp_m2_26_6_r,temp_m2_26_6_i,temp_m2_26_8_r,temp_m2_26_8_i,temp_m2_28_6_r,temp_m2_28_6_i,temp_m2_28_8_r,temp_m2_28_8_i,temp_b2_26_6_r,temp_b2_26_6_i,temp_b2_26_8_r,temp_b2_26_8_i,temp_b2_28_6_r,temp_b2_28_6_i,temp_b2_28_8_r,temp_b2_28_8_i);
MULT MULT457 (clk,temp_b1_25_9_r,temp_b1_25_9_i,temp_b1_25_11_r,temp_b1_25_11_i,temp_b1_27_9_r,temp_b1_27_9_i,temp_b1_27_11_r,temp_b1_27_11_i,temp_m2_25_9_r,temp_m2_25_9_i,temp_m2_25_11_r,temp_m2_25_11_i,temp_m2_27_9_r,temp_m2_27_9_i,temp_m2_27_11_r,temp_m2_27_11_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly457 (clk,temp_m2_25_9_r,temp_m2_25_9_i,temp_m2_25_11_r,temp_m2_25_11_i,temp_m2_27_9_r,temp_m2_27_9_i,temp_m2_27_11_r,temp_m2_27_11_i,temp_b2_25_9_r,temp_b2_25_9_i,temp_b2_25_11_r,temp_b2_25_11_i,temp_b2_27_9_r,temp_b2_27_9_i,temp_b2_27_11_r,temp_b2_27_11_i);
MULT MULT458 (clk,temp_b1_25_10_r,temp_b1_25_10_i,temp_b1_25_12_r,temp_b1_25_12_i,temp_b1_27_10_r,temp_b1_27_10_i,temp_b1_27_12_r,temp_b1_27_12_i,temp_m2_25_10_r,temp_m2_25_10_i,temp_m2_25_12_r,temp_m2_25_12_i,temp_m2_27_10_r,temp_m2_27_10_i,temp_m2_27_12_r,temp_m2_27_12_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly458 (clk,temp_m2_25_10_r,temp_m2_25_10_i,temp_m2_25_12_r,temp_m2_25_12_i,temp_m2_27_10_r,temp_m2_27_10_i,temp_m2_27_12_r,temp_m2_27_12_i,temp_b2_25_10_r,temp_b2_25_10_i,temp_b2_25_12_r,temp_b2_25_12_i,temp_b2_27_10_r,temp_b2_27_10_i,temp_b2_27_12_r,temp_b2_27_12_i);
MULT MULT459 (clk,temp_b1_26_9_r,temp_b1_26_9_i,temp_b1_26_11_r,temp_b1_26_11_i,temp_b1_28_9_r,temp_b1_28_9_i,temp_b1_28_11_r,temp_b1_28_11_i,temp_m2_26_9_r,temp_m2_26_9_i,temp_m2_26_11_r,temp_m2_26_11_i,temp_m2_28_9_r,temp_m2_28_9_i,temp_m2_28_11_r,temp_m2_28_11_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly459 (clk,temp_m2_26_9_r,temp_m2_26_9_i,temp_m2_26_11_r,temp_m2_26_11_i,temp_m2_28_9_r,temp_m2_28_9_i,temp_m2_28_11_r,temp_m2_28_11_i,temp_b2_26_9_r,temp_b2_26_9_i,temp_b2_26_11_r,temp_b2_26_11_i,temp_b2_28_9_r,temp_b2_28_9_i,temp_b2_28_11_r,temp_b2_28_11_i);
MULT MULT460 (clk,temp_b1_26_10_r,temp_b1_26_10_i,temp_b1_26_12_r,temp_b1_26_12_i,temp_b1_28_10_r,temp_b1_28_10_i,temp_b1_28_12_r,temp_b1_28_12_i,temp_m2_26_10_r,temp_m2_26_10_i,temp_m2_26_12_r,temp_m2_26_12_i,temp_m2_28_10_r,temp_m2_28_10_i,temp_m2_28_12_r,temp_m2_28_12_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly460 (clk,temp_m2_26_10_r,temp_m2_26_10_i,temp_m2_26_12_r,temp_m2_26_12_i,temp_m2_28_10_r,temp_m2_28_10_i,temp_m2_28_12_r,temp_m2_28_12_i,temp_b2_26_10_r,temp_b2_26_10_i,temp_b2_26_12_r,temp_b2_26_12_i,temp_b2_28_10_r,temp_b2_28_10_i,temp_b2_28_12_r,temp_b2_28_12_i);
MULT MULT461 (clk,temp_b1_25_13_r,temp_b1_25_13_i,temp_b1_25_15_r,temp_b1_25_15_i,temp_b1_27_13_r,temp_b1_27_13_i,temp_b1_27_15_r,temp_b1_27_15_i,temp_m2_25_13_r,temp_m2_25_13_i,temp_m2_25_15_r,temp_m2_25_15_i,temp_m2_27_13_r,temp_m2_27_13_i,temp_m2_27_15_r,temp_m2_27_15_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly461 (clk,temp_m2_25_13_r,temp_m2_25_13_i,temp_m2_25_15_r,temp_m2_25_15_i,temp_m2_27_13_r,temp_m2_27_13_i,temp_m2_27_15_r,temp_m2_27_15_i,temp_b2_25_13_r,temp_b2_25_13_i,temp_b2_25_15_r,temp_b2_25_15_i,temp_b2_27_13_r,temp_b2_27_13_i,temp_b2_27_15_r,temp_b2_27_15_i);
MULT MULT462 (clk,temp_b1_25_14_r,temp_b1_25_14_i,temp_b1_25_16_r,temp_b1_25_16_i,temp_b1_27_14_r,temp_b1_27_14_i,temp_b1_27_16_r,temp_b1_27_16_i,temp_m2_25_14_r,temp_m2_25_14_i,temp_m2_25_16_r,temp_m2_25_16_i,temp_m2_27_14_r,temp_m2_27_14_i,temp_m2_27_16_r,temp_m2_27_16_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly462 (clk,temp_m2_25_14_r,temp_m2_25_14_i,temp_m2_25_16_r,temp_m2_25_16_i,temp_m2_27_14_r,temp_m2_27_14_i,temp_m2_27_16_r,temp_m2_27_16_i,temp_b2_25_14_r,temp_b2_25_14_i,temp_b2_25_16_r,temp_b2_25_16_i,temp_b2_27_14_r,temp_b2_27_14_i,temp_b2_27_16_r,temp_b2_27_16_i);
MULT MULT463 (clk,temp_b1_26_13_r,temp_b1_26_13_i,temp_b1_26_15_r,temp_b1_26_15_i,temp_b1_28_13_r,temp_b1_28_13_i,temp_b1_28_15_r,temp_b1_28_15_i,temp_m2_26_13_r,temp_m2_26_13_i,temp_m2_26_15_r,temp_m2_26_15_i,temp_m2_28_13_r,temp_m2_28_13_i,temp_m2_28_15_r,temp_m2_28_15_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly463 (clk,temp_m2_26_13_r,temp_m2_26_13_i,temp_m2_26_15_r,temp_m2_26_15_i,temp_m2_28_13_r,temp_m2_28_13_i,temp_m2_28_15_r,temp_m2_28_15_i,temp_b2_26_13_r,temp_b2_26_13_i,temp_b2_26_15_r,temp_b2_26_15_i,temp_b2_28_13_r,temp_b2_28_13_i,temp_b2_28_15_r,temp_b2_28_15_i);
MULT MULT464 (clk,temp_b1_26_14_r,temp_b1_26_14_i,temp_b1_26_16_r,temp_b1_26_16_i,temp_b1_28_14_r,temp_b1_28_14_i,temp_b1_28_16_r,temp_b1_28_16_i,temp_m2_26_14_r,temp_m2_26_14_i,temp_m2_26_16_r,temp_m2_26_16_i,temp_m2_28_14_r,temp_m2_28_14_i,temp_m2_28_16_r,temp_m2_28_16_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly464 (clk,temp_m2_26_14_r,temp_m2_26_14_i,temp_m2_26_16_r,temp_m2_26_16_i,temp_m2_28_14_r,temp_m2_28_14_i,temp_m2_28_16_r,temp_m2_28_16_i,temp_b2_26_14_r,temp_b2_26_14_i,temp_b2_26_16_r,temp_b2_26_16_i,temp_b2_28_14_r,temp_b2_28_14_i,temp_b2_28_16_r,temp_b2_28_16_i);
MULT MULT465 (clk,temp_b1_25_17_r,temp_b1_25_17_i,temp_b1_25_19_r,temp_b1_25_19_i,temp_b1_27_17_r,temp_b1_27_17_i,temp_b1_27_19_r,temp_b1_27_19_i,temp_m2_25_17_r,temp_m2_25_17_i,temp_m2_25_19_r,temp_m2_25_19_i,temp_m2_27_17_r,temp_m2_27_17_i,temp_m2_27_19_r,temp_m2_27_19_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly465 (clk,temp_m2_25_17_r,temp_m2_25_17_i,temp_m2_25_19_r,temp_m2_25_19_i,temp_m2_27_17_r,temp_m2_27_17_i,temp_m2_27_19_r,temp_m2_27_19_i,temp_b2_25_17_r,temp_b2_25_17_i,temp_b2_25_19_r,temp_b2_25_19_i,temp_b2_27_17_r,temp_b2_27_17_i,temp_b2_27_19_r,temp_b2_27_19_i);
MULT MULT466 (clk,temp_b1_25_18_r,temp_b1_25_18_i,temp_b1_25_20_r,temp_b1_25_20_i,temp_b1_27_18_r,temp_b1_27_18_i,temp_b1_27_20_r,temp_b1_27_20_i,temp_m2_25_18_r,temp_m2_25_18_i,temp_m2_25_20_r,temp_m2_25_20_i,temp_m2_27_18_r,temp_m2_27_18_i,temp_m2_27_20_r,temp_m2_27_20_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly466 (clk,temp_m2_25_18_r,temp_m2_25_18_i,temp_m2_25_20_r,temp_m2_25_20_i,temp_m2_27_18_r,temp_m2_27_18_i,temp_m2_27_20_r,temp_m2_27_20_i,temp_b2_25_18_r,temp_b2_25_18_i,temp_b2_25_20_r,temp_b2_25_20_i,temp_b2_27_18_r,temp_b2_27_18_i,temp_b2_27_20_r,temp_b2_27_20_i);
MULT MULT467 (clk,temp_b1_26_17_r,temp_b1_26_17_i,temp_b1_26_19_r,temp_b1_26_19_i,temp_b1_28_17_r,temp_b1_28_17_i,temp_b1_28_19_r,temp_b1_28_19_i,temp_m2_26_17_r,temp_m2_26_17_i,temp_m2_26_19_r,temp_m2_26_19_i,temp_m2_28_17_r,temp_m2_28_17_i,temp_m2_28_19_r,temp_m2_28_19_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly467 (clk,temp_m2_26_17_r,temp_m2_26_17_i,temp_m2_26_19_r,temp_m2_26_19_i,temp_m2_28_17_r,temp_m2_28_17_i,temp_m2_28_19_r,temp_m2_28_19_i,temp_b2_26_17_r,temp_b2_26_17_i,temp_b2_26_19_r,temp_b2_26_19_i,temp_b2_28_17_r,temp_b2_28_17_i,temp_b2_28_19_r,temp_b2_28_19_i);
MULT MULT468 (clk,temp_b1_26_18_r,temp_b1_26_18_i,temp_b1_26_20_r,temp_b1_26_20_i,temp_b1_28_18_r,temp_b1_28_18_i,temp_b1_28_20_r,temp_b1_28_20_i,temp_m2_26_18_r,temp_m2_26_18_i,temp_m2_26_20_r,temp_m2_26_20_i,temp_m2_28_18_r,temp_m2_28_18_i,temp_m2_28_20_r,temp_m2_28_20_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly468 (clk,temp_m2_26_18_r,temp_m2_26_18_i,temp_m2_26_20_r,temp_m2_26_20_i,temp_m2_28_18_r,temp_m2_28_18_i,temp_m2_28_20_r,temp_m2_28_20_i,temp_b2_26_18_r,temp_b2_26_18_i,temp_b2_26_20_r,temp_b2_26_20_i,temp_b2_28_18_r,temp_b2_28_18_i,temp_b2_28_20_r,temp_b2_28_20_i);
MULT MULT469 (clk,temp_b1_25_21_r,temp_b1_25_21_i,temp_b1_25_23_r,temp_b1_25_23_i,temp_b1_27_21_r,temp_b1_27_21_i,temp_b1_27_23_r,temp_b1_27_23_i,temp_m2_25_21_r,temp_m2_25_21_i,temp_m2_25_23_r,temp_m2_25_23_i,temp_m2_27_21_r,temp_m2_27_21_i,temp_m2_27_23_r,temp_m2_27_23_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly469 (clk,temp_m2_25_21_r,temp_m2_25_21_i,temp_m2_25_23_r,temp_m2_25_23_i,temp_m2_27_21_r,temp_m2_27_21_i,temp_m2_27_23_r,temp_m2_27_23_i,temp_b2_25_21_r,temp_b2_25_21_i,temp_b2_25_23_r,temp_b2_25_23_i,temp_b2_27_21_r,temp_b2_27_21_i,temp_b2_27_23_r,temp_b2_27_23_i);
MULT MULT470 (clk,temp_b1_25_22_r,temp_b1_25_22_i,temp_b1_25_24_r,temp_b1_25_24_i,temp_b1_27_22_r,temp_b1_27_22_i,temp_b1_27_24_r,temp_b1_27_24_i,temp_m2_25_22_r,temp_m2_25_22_i,temp_m2_25_24_r,temp_m2_25_24_i,temp_m2_27_22_r,temp_m2_27_22_i,temp_m2_27_24_r,temp_m2_27_24_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly470 (clk,temp_m2_25_22_r,temp_m2_25_22_i,temp_m2_25_24_r,temp_m2_25_24_i,temp_m2_27_22_r,temp_m2_27_22_i,temp_m2_27_24_r,temp_m2_27_24_i,temp_b2_25_22_r,temp_b2_25_22_i,temp_b2_25_24_r,temp_b2_25_24_i,temp_b2_27_22_r,temp_b2_27_22_i,temp_b2_27_24_r,temp_b2_27_24_i);
MULT MULT471 (clk,temp_b1_26_21_r,temp_b1_26_21_i,temp_b1_26_23_r,temp_b1_26_23_i,temp_b1_28_21_r,temp_b1_28_21_i,temp_b1_28_23_r,temp_b1_28_23_i,temp_m2_26_21_r,temp_m2_26_21_i,temp_m2_26_23_r,temp_m2_26_23_i,temp_m2_28_21_r,temp_m2_28_21_i,temp_m2_28_23_r,temp_m2_28_23_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly471 (clk,temp_m2_26_21_r,temp_m2_26_21_i,temp_m2_26_23_r,temp_m2_26_23_i,temp_m2_28_21_r,temp_m2_28_21_i,temp_m2_28_23_r,temp_m2_28_23_i,temp_b2_26_21_r,temp_b2_26_21_i,temp_b2_26_23_r,temp_b2_26_23_i,temp_b2_28_21_r,temp_b2_28_21_i,temp_b2_28_23_r,temp_b2_28_23_i);
MULT MULT472 (clk,temp_b1_26_22_r,temp_b1_26_22_i,temp_b1_26_24_r,temp_b1_26_24_i,temp_b1_28_22_r,temp_b1_28_22_i,temp_b1_28_24_r,temp_b1_28_24_i,temp_m2_26_22_r,temp_m2_26_22_i,temp_m2_26_24_r,temp_m2_26_24_i,temp_m2_28_22_r,temp_m2_28_22_i,temp_m2_28_24_r,temp_m2_28_24_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly472 (clk,temp_m2_26_22_r,temp_m2_26_22_i,temp_m2_26_24_r,temp_m2_26_24_i,temp_m2_28_22_r,temp_m2_28_22_i,temp_m2_28_24_r,temp_m2_28_24_i,temp_b2_26_22_r,temp_b2_26_22_i,temp_b2_26_24_r,temp_b2_26_24_i,temp_b2_28_22_r,temp_b2_28_22_i,temp_b2_28_24_r,temp_b2_28_24_i);
MULT MULT473 (clk,temp_b1_25_25_r,temp_b1_25_25_i,temp_b1_25_27_r,temp_b1_25_27_i,temp_b1_27_25_r,temp_b1_27_25_i,temp_b1_27_27_r,temp_b1_27_27_i,temp_m2_25_25_r,temp_m2_25_25_i,temp_m2_25_27_r,temp_m2_25_27_i,temp_m2_27_25_r,temp_m2_27_25_i,temp_m2_27_27_r,temp_m2_27_27_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly473 (clk,temp_m2_25_25_r,temp_m2_25_25_i,temp_m2_25_27_r,temp_m2_25_27_i,temp_m2_27_25_r,temp_m2_27_25_i,temp_m2_27_27_r,temp_m2_27_27_i,temp_b2_25_25_r,temp_b2_25_25_i,temp_b2_25_27_r,temp_b2_25_27_i,temp_b2_27_25_r,temp_b2_27_25_i,temp_b2_27_27_r,temp_b2_27_27_i);
MULT MULT474 (clk,temp_b1_25_26_r,temp_b1_25_26_i,temp_b1_25_28_r,temp_b1_25_28_i,temp_b1_27_26_r,temp_b1_27_26_i,temp_b1_27_28_r,temp_b1_27_28_i,temp_m2_25_26_r,temp_m2_25_26_i,temp_m2_25_28_r,temp_m2_25_28_i,temp_m2_27_26_r,temp_m2_27_26_i,temp_m2_27_28_r,temp_m2_27_28_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly474 (clk,temp_m2_25_26_r,temp_m2_25_26_i,temp_m2_25_28_r,temp_m2_25_28_i,temp_m2_27_26_r,temp_m2_27_26_i,temp_m2_27_28_r,temp_m2_27_28_i,temp_b2_25_26_r,temp_b2_25_26_i,temp_b2_25_28_r,temp_b2_25_28_i,temp_b2_27_26_r,temp_b2_27_26_i,temp_b2_27_28_r,temp_b2_27_28_i);
MULT MULT475 (clk,temp_b1_26_25_r,temp_b1_26_25_i,temp_b1_26_27_r,temp_b1_26_27_i,temp_b1_28_25_r,temp_b1_28_25_i,temp_b1_28_27_r,temp_b1_28_27_i,temp_m2_26_25_r,temp_m2_26_25_i,temp_m2_26_27_r,temp_m2_26_27_i,temp_m2_28_25_r,temp_m2_28_25_i,temp_m2_28_27_r,temp_m2_28_27_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly475 (clk,temp_m2_26_25_r,temp_m2_26_25_i,temp_m2_26_27_r,temp_m2_26_27_i,temp_m2_28_25_r,temp_m2_28_25_i,temp_m2_28_27_r,temp_m2_28_27_i,temp_b2_26_25_r,temp_b2_26_25_i,temp_b2_26_27_r,temp_b2_26_27_i,temp_b2_28_25_r,temp_b2_28_25_i,temp_b2_28_27_r,temp_b2_28_27_i);
MULT MULT476 (clk,temp_b1_26_26_r,temp_b1_26_26_i,temp_b1_26_28_r,temp_b1_26_28_i,temp_b1_28_26_r,temp_b1_28_26_i,temp_b1_28_28_r,temp_b1_28_28_i,temp_m2_26_26_r,temp_m2_26_26_i,temp_m2_26_28_r,temp_m2_26_28_i,temp_m2_28_26_r,temp_m2_28_26_i,temp_m2_28_28_r,temp_m2_28_28_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly476 (clk,temp_m2_26_26_r,temp_m2_26_26_i,temp_m2_26_28_r,temp_m2_26_28_i,temp_m2_28_26_r,temp_m2_28_26_i,temp_m2_28_28_r,temp_m2_28_28_i,temp_b2_26_26_r,temp_b2_26_26_i,temp_b2_26_28_r,temp_b2_26_28_i,temp_b2_28_26_r,temp_b2_28_26_i,temp_b2_28_28_r,temp_b2_28_28_i);
MULT MULT477 (clk,temp_b1_25_29_r,temp_b1_25_29_i,temp_b1_25_31_r,temp_b1_25_31_i,temp_b1_27_29_r,temp_b1_27_29_i,temp_b1_27_31_r,temp_b1_27_31_i,temp_m2_25_29_r,temp_m2_25_29_i,temp_m2_25_31_r,temp_m2_25_31_i,temp_m2_27_29_r,temp_m2_27_29_i,temp_m2_27_31_r,temp_m2_27_31_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly477 (clk,temp_m2_25_29_r,temp_m2_25_29_i,temp_m2_25_31_r,temp_m2_25_31_i,temp_m2_27_29_r,temp_m2_27_29_i,temp_m2_27_31_r,temp_m2_27_31_i,temp_b2_25_29_r,temp_b2_25_29_i,temp_b2_25_31_r,temp_b2_25_31_i,temp_b2_27_29_r,temp_b2_27_29_i,temp_b2_27_31_r,temp_b2_27_31_i);
MULT MULT478 (clk,temp_b1_25_30_r,temp_b1_25_30_i,temp_b1_25_32_r,temp_b1_25_32_i,temp_b1_27_30_r,temp_b1_27_30_i,temp_b1_27_32_r,temp_b1_27_32_i,temp_m2_25_30_r,temp_m2_25_30_i,temp_m2_25_32_r,temp_m2_25_32_i,temp_m2_27_30_r,temp_m2_27_30_i,temp_m2_27_32_r,temp_m2_27_32_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly478 (clk,temp_m2_25_30_r,temp_m2_25_30_i,temp_m2_25_32_r,temp_m2_25_32_i,temp_m2_27_30_r,temp_m2_27_30_i,temp_m2_27_32_r,temp_m2_27_32_i,temp_b2_25_30_r,temp_b2_25_30_i,temp_b2_25_32_r,temp_b2_25_32_i,temp_b2_27_30_r,temp_b2_27_30_i,temp_b2_27_32_r,temp_b2_27_32_i);
MULT MULT479 (clk,temp_b1_26_29_r,temp_b1_26_29_i,temp_b1_26_31_r,temp_b1_26_31_i,temp_b1_28_29_r,temp_b1_28_29_i,temp_b1_28_31_r,temp_b1_28_31_i,temp_m2_26_29_r,temp_m2_26_29_i,temp_m2_26_31_r,temp_m2_26_31_i,temp_m2_28_29_r,temp_m2_28_29_i,temp_m2_28_31_r,temp_m2_28_31_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly479 (clk,temp_m2_26_29_r,temp_m2_26_29_i,temp_m2_26_31_r,temp_m2_26_31_i,temp_m2_28_29_r,temp_m2_28_29_i,temp_m2_28_31_r,temp_m2_28_31_i,temp_b2_26_29_r,temp_b2_26_29_i,temp_b2_26_31_r,temp_b2_26_31_i,temp_b2_28_29_r,temp_b2_28_29_i,temp_b2_28_31_r,temp_b2_28_31_i);
MULT MULT480 (clk,temp_b1_26_30_r,temp_b1_26_30_i,temp_b1_26_32_r,temp_b1_26_32_i,temp_b1_28_30_r,temp_b1_28_30_i,temp_b1_28_32_r,temp_b1_28_32_i,temp_m2_26_30_r,temp_m2_26_30_i,temp_m2_26_32_r,temp_m2_26_32_i,temp_m2_28_30_r,temp_m2_28_30_i,temp_m2_28_32_r,temp_m2_28_32_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly480 (clk,temp_m2_26_30_r,temp_m2_26_30_i,temp_m2_26_32_r,temp_m2_26_32_i,temp_m2_28_30_r,temp_m2_28_30_i,temp_m2_28_32_r,temp_m2_28_32_i,temp_b2_26_30_r,temp_b2_26_30_i,temp_b2_26_32_r,temp_b2_26_32_i,temp_b2_28_30_r,temp_b2_28_30_i,temp_b2_28_32_r,temp_b2_28_32_i);
MULT MULT481 (clk,temp_b1_29_1_r,temp_b1_29_1_i,temp_b1_29_3_r,temp_b1_29_3_i,temp_b1_31_1_r,temp_b1_31_1_i,temp_b1_31_3_r,temp_b1_31_3_i,temp_m2_29_1_r,temp_m2_29_1_i,temp_m2_29_3_r,temp_m2_29_3_i,temp_m2_31_1_r,temp_m2_31_1_i,temp_m2_31_3_r,temp_m2_31_3_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly481 (clk,temp_m2_29_1_r,temp_m2_29_1_i,temp_m2_29_3_r,temp_m2_29_3_i,temp_m2_31_1_r,temp_m2_31_1_i,temp_m2_31_3_r,temp_m2_31_3_i,temp_b2_29_1_r,temp_b2_29_1_i,temp_b2_29_3_r,temp_b2_29_3_i,temp_b2_31_1_r,temp_b2_31_1_i,temp_b2_31_3_r,temp_b2_31_3_i);
MULT MULT482 (clk,temp_b1_29_2_r,temp_b1_29_2_i,temp_b1_29_4_r,temp_b1_29_4_i,temp_b1_31_2_r,temp_b1_31_2_i,temp_b1_31_4_r,temp_b1_31_4_i,temp_m2_29_2_r,temp_m2_29_2_i,temp_m2_29_4_r,temp_m2_29_4_i,temp_m2_31_2_r,temp_m2_31_2_i,temp_m2_31_4_r,temp_m2_31_4_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly482 (clk,temp_m2_29_2_r,temp_m2_29_2_i,temp_m2_29_4_r,temp_m2_29_4_i,temp_m2_31_2_r,temp_m2_31_2_i,temp_m2_31_4_r,temp_m2_31_4_i,temp_b2_29_2_r,temp_b2_29_2_i,temp_b2_29_4_r,temp_b2_29_4_i,temp_b2_31_2_r,temp_b2_31_2_i,temp_b2_31_4_r,temp_b2_31_4_i);
MULT MULT483 (clk,temp_b1_30_1_r,temp_b1_30_1_i,temp_b1_30_3_r,temp_b1_30_3_i,temp_b1_32_1_r,temp_b1_32_1_i,temp_b1_32_3_r,temp_b1_32_3_i,temp_m2_30_1_r,temp_m2_30_1_i,temp_m2_30_3_r,temp_m2_30_3_i,temp_m2_32_1_r,temp_m2_32_1_i,temp_m2_32_3_r,temp_m2_32_3_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly483 (clk,temp_m2_30_1_r,temp_m2_30_1_i,temp_m2_30_3_r,temp_m2_30_3_i,temp_m2_32_1_r,temp_m2_32_1_i,temp_m2_32_3_r,temp_m2_32_3_i,temp_b2_30_1_r,temp_b2_30_1_i,temp_b2_30_3_r,temp_b2_30_3_i,temp_b2_32_1_r,temp_b2_32_1_i,temp_b2_32_3_r,temp_b2_32_3_i);
MULT MULT484 (clk,temp_b1_30_2_r,temp_b1_30_2_i,temp_b1_30_4_r,temp_b1_30_4_i,temp_b1_32_2_r,temp_b1_32_2_i,temp_b1_32_4_r,temp_b1_32_4_i,temp_m2_30_2_r,temp_m2_30_2_i,temp_m2_30_4_r,temp_m2_30_4_i,temp_m2_32_2_r,temp_m2_32_2_i,temp_m2_32_4_r,temp_m2_32_4_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly484 (clk,temp_m2_30_2_r,temp_m2_30_2_i,temp_m2_30_4_r,temp_m2_30_4_i,temp_m2_32_2_r,temp_m2_32_2_i,temp_m2_32_4_r,temp_m2_32_4_i,temp_b2_30_2_r,temp_b2_30_2_i,temp_b2_30_4_r,temp_b2_30_4_i,temp_b2_32_2_r,temp_b2_32_2_i,temp_b2_32_4_r,temp_b2_32_4_i);
MULT MULT485 (clk,temp_b1_29_5_r,temp_b1_29_5_i,temp_b1_29_7_r,temp_b1_29_7_i,temp_b1_31_5_r,temp_b1_31_5_i,temp_b1_31_7_r,temp_b1_31_7_i,temp_m2_29_5_r,temp_m2_29_5_i,temp_m2_29_7_r,temp_m2_29_7_i,temp_m2_31_5_r,temp_m2_31_5_i,temp_m2_31_7_r,temp_m2_31_7_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly485 (clk,temp_m2_29_5_r,temp_m2_29_5_i,temp_m2_29_7_r,temp_m2_29_7_i,temp_m2_31_5_r,temp_m2_31_5_i,temp_m2_31_7_r,temp_m2_31_7_i,temp_b2_29_5_r,temp_b2_29_5_i,temp_b2_29_7_r,temp_b2_29_7_i,temp_b2_31_5_r,temp_b2_31_5_i,temp_b2_31_7_r,temp_b2_31_7_i);
MULT MULT486 (clk,temp_b1_29_6_r,temp_b1_29_6_i,temp_b1_29_8_r,temp_b1_29_8_i,temp_b1_31_6_r,temp_b1_31_6_i,temp_b1_31_8_r,temp_b1_31_8_i,temp_m2_29_6_r,temp_m2_29_6_i,temp_m2_29_8_r,temp_m2_29_8_i,temp_m2_31_6_r,temp_m2_31_6_i,temp_m2_31_8_r,temp_m2_31_8_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly486 (clk,temp_m2_29_6_r,temp_m2_29_6_i,temp_m2_29_8_r,temp_m2_29_8_i,temp_m2_31_6_r,temp_m2_31_6_i,temp_m2_31_8_r,temp_m2_31_8_i,temp_b2_29_6_r,temp_b2_29_6_i,temp_b2_29_8_r,temp_b2_29_8_i,temp_b2_31_6_r,temp_b2_31_6_i,temp_b2_31_8_r,temp_b2_31_8_i);
MULT MULT487 (clk,temp_b1_30_5_r,temp_b1_30_5_i,temp_b1_30_7_r,temp_b1_30_7_i,temp_b1_32_5_r,temp_b1_32_5_i,temp_b1_32_7_r,temp_b1_32_7_i,temp_m2_30_5_r,temp_m2_30_5_i,temp_m2_30_7_r,temp_m2_30_7_i,temp_m2_32_5_r,temp_m2_32_5_i,temp_m2_32_7_r,temp_m2_32_7_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly487 (clk,temp_m2_30_5_r,temp_m2_30_5_i,temp_m2_30_7_r,temp_m2_30_7_i,temp_m2_32_5_r,temp_m2_32_5_i,temp_m2_32_7_r,temp_m2_32_7_i,temp_b2_30_5_r,temp_b2_30_5_i,temp_b2_30_7_r,temp_b2_30_7_i,temp_b2_32_5_r,temp_b2_32_5_i,temp_b2_32_7_r,temp_b2_32_7_i);
MULT MULT488 (clk,temp_b1_30_6_r,temp_b1_30_6_i,temp_b1_30_8_r,temp_b1_30_8_i,temp_b1_32_6_r,temp_b1_32_6_i,temp_b1_32_8_r,temp_b1_32_8_i,temp_m2_30_6_r,temp_m2_30_6_i,temp_m2_30_8_r,temp_m2_30_8_i,temp_m2_32_6_r,temp_m2_32_6_i,temp_m2_32_8_r,temp_m2_32_8_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly488 (clk,temp_m2_30_6_r,temp_m2_30_6_i,temp_m2_30_8_r,temp_m2_30_8_i,temp_m2_32_6_r,temp_m2_32_6_i,temp_m2_32_8_r,temp_m2_32_8_i,temp_b2_30_6_r,temp_b2_30_6_i,temp_b2_30_8_r,temp_b2_30_8_i,temp_b2_32_6_r,temp_b2_32_6_i,temp_b2_32_8_r,temp_b2_32_8_i);
MULT MULT489 (clk,temp_b1_29_9_r,temp_b1_29_9_i,temp_b1_29_11_r,temp_b1_29_11_i,temp_b1_31_9_r,temp_b1_31_9_i,temp_b1_31_11_r,temp_b1_31_11_i,temp_m2_29_9_r,temp_m2_29_9_i,temp_m2_29_11_r,temp_m2_29_11_i,temp_m2_31_9_r,temp_m2_31_9_i,temp_m2_31_11_r,temp_m2_31_11_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly489 (clk,temp_m2_29_9_r,temp_m2_29_9_i,temp_m2_29_11_r,temp_m2_29_11_i,temp_m2_31_9_r,temp_m2_31_9_i,temp_m2_31_11_r,temp_m2_31_11_i,temp_b2_29_9_r,temp_b2_29_9_i,temp_b2_29_11_r,temp_b2_29_11_i,temp_b2_31_9_r,temp_b2_31_9_i,temp_b2_31_11_r,temp_b2_31_11_i);
MULT MULT490 (clk,temp_b1_29_10_r,temp_b1_29_10_i,temp_b1_29_12_r,temp_b1_29_12_i,temp_b1_31_10_r,temp_b1_31_10_i,temp_b1_31_12_r,temp_b1_31_12_i,temp_m2_29_10_r,temp_m2_29_10_i,temp_m2_29_12_r,temp_m2_29_12_i,temp_m2_31_10_r,temp_m2_31_10_i,temp_m2_31_12_r,temp_m2_31_12_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly490 (clk,temp_m2_29_10_r,temp_m2_29_10_i,temp_m2_29_12_r,temp_m2_29_12_i,temp_m2_31_10_r,temp_m2_31_10_i,temp_m2_31_12_r,temp_m2_31_12_i,temp_b2_29_10_r,temp_b2_29_10_i,temp_b2_29_12_r,temp_b2_29_12_i,temp_b2_31_10_r,temp_b2_31_10_i,temp_b2_31_12_r,temp_b2_31_12_i);
MULT MULT491 (clk,temp_b1_30_9_r,temp_b1_30_9_i,temp_b1_30_11_r,temp_b1_30_11_i,temp_b1_32_9_r,temp_b1_32_9_i,temp_b1_32_11_r,temp_b1_32_11_i,temp_m2_30_9_r,temp_m2_30_9_i,temp_m2_30_11_r,temp_m2_30_11_i,temp_m2_32_9_r,temp_m2_32_9_i,temp_m2_32_11_r,temp_m2_32_11_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly491 (clk,temp_m2_30_9_r,temp_m2_30_9_i,temp_m2_30_11_r,temp_m2_30_11_i,temp_m2_32_9_r,temp_m2_32_9_i,temp_m2_32_11_r,temp_m2_32_11_i,temp_b2_30_9_r,temp_b2_30_9_i,temp_b2_30_11_r,temp_b2_30_11_i,temp_b2_32_9_r,temp_b2_32_9_i,temp_b2_32_11_r,temp_b2_32_11_i);
MULT MULT492 (clk,temp_b1_30_10_r,temp_b1_30_10_i,temp_b1_30_12_r,temp_b1_30_12_i,temp_b1_32_10_r,temp_b1_32_10_i,temp_b1_32_12_r,temp_b1_32_12_i,temp_m2_30_10_r,temp_m2_30_10_i,temp_m2_30_12_r,temp_m2_30_12_i,temp_m2_32_10_r,temp_m2_32_10_i,temp_m2_32_12_r,temp_m2_32_12_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly492 (clk,temp_m2_30_10_r,temp_m2_30_10_i,temp_m2_30_12_r,temp_m2_30_12_i,temp_m2_32_10_r,temp_m2_32_10_i,temp_m2_32_12_r,temp_m2_32_12_i,temp_b2_30_10_r,temp_b2_30_10_i,temp_b2_30_12_r,temp_b2_30_12_i,temp_b2_32_10_r,temp_b2_32_10_i,temp_b2_32_12_r,temp_b2_32_12_i);
MULT MULT493 (clk,temp_b1_29_13_r,temp_b1_29_13_i,temp_b1_29_15_r,temp_b1_29_15_i,temp_b1_31_13_r,temp_b1_31_13_i,temp_b1_31_15_r,temp_b1_31_15_i,temp_m2_29_13_r,temp_m2_29_13_i,temp_m2_29_15_r,temp_m2_29_15_i,temp_m2_31_13_r,temp_m2_31_13_i,temp_m2_31_15_r,temp_m2_31_15_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly493 (clk,temp_m2_29_13_r,temp_m2_29_13_i,temp_m2_29_15_r,temp_m2_29_15_i,temp_m2_31_13_r,temp_m2_31_13_i,temp_m2_31_15_r,temp_m2_31_15_i,temp_b2_29_13_r,temp_b2_29_13_i,temp_b2_29_15_r,temp_b2_29_15_i,temp_b2_31_13_r,temp_b2_31_13_i,temp_b2_31_15_r,temp_b2_31_15_i);
MULT MULT494 (clk,temp_b1_29_14_r,temp_b1_29_14_i,temp_b1_29_16_r,temp_b1_29_16_i,temp_b1_31_14_r,temp_b1_31_14_i,temp_b1_31_16_r,temp_b1_31_16_i,temp_m2_29_14_r,temp_m2_29_14_i,temp_m2_29_16_r,temp_m2_29_16_i,temp_m2_31_14_r,temp_m2_31_14_i,temp_m2_31_16_r,temp_m2_31_16_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly494 (clk,temp_m2_29_14_r,temp_m2_29_14_i,temp_m2_29_16_r,temp_m2_29_16_i,temp_m2_31_14_r,temp_m2_31_14_i,temp_m2_31_16_r,temp_m2_31_16_i,temp_b2_29_14_r,temp_b2_29_14_i,temp_b2_29_16_r,temp_b2_29_16_i,temp_b2_31_14_r,temp_b2_31_14_i,temp_b2_31_16_r,temp_b2_31_16_i);
MULT MULT495 (clk,temp_b1_30_13_r,temp_b1_30_13_i,temp_b1_30_15_r,temp_b1_30_15_i,temp_b1_32_13_r,temp_b1_32_13_i,temp_b1_32_15_r,temp_b1_32_15_i,temp_m2_30_13_r,temp_m2_30_13_i,temp_m2_30_15_r,temp_m2_30_15_i,temp_m2_32_13_r,temp_m2_32_13_i,temp_m2_32_15_r,temp_m2_32_15_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly495 (clk,temp_m2_30_13_r,temp_m2_30_13_i,temp_m2_30_15_r,temp_m2_30_15_i,temp_m2_32_13_r,temp_m2_32_13_i,temp_m2_32_15_r,temp_m2_32_15_i,temp_b2_30_13_r,temp_b2_30_13_i,temp_b2_30_15_r,temp_b2_30_15_i,temp_b2_32_13_r,temp_b2_32_13_i,temp_b2_32_15_r,temp_b2_32_15_i);
MULT MULT496 (clk,temp_b1_30_14_r,temp_b1_30_14_i,temp_b1_30_16_r,temp_b1_30_16_i,temp_b1_32_14_r,temp_b1_32_14_i,temp_b1_32_16_r,temp_b1_32_16_i,temp_m2_30_14_r,temp_m2_30_14_i,temp_m2_30_16_r,temp_m2_30_16_i,temp_m2_32_14_r,temp_m2_32_14_i,temp_m2_32_16_r,temp_m2_32_16_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly496 (clk,temp_m2_30_14_r,temp_m2_30_14_i,temp_m2_30_16_r,temp_m2_30_16_i,temp_m2_32_14_r,temp_m2_32_14_i,temp_m2_32_16_r,temp_m2_32_16_i,temp_b2_30_14_r,temp_b2_30_14_i,temp_b2_30_16_r,temp_b2_30_16_i,temp_b2_32_14_r,temp_b2_32_14_i,temp_b2_32_16_r,temp_b2_32_16_i);
MULT MULT497 (clk,temp_b1_29_17_r,temp_b1_29_17_i,temp_b1_29_19_r,temp_b1_29_19_i,temp_b1_31_17_r,temp_b1_31_17_i,temp_b1_31_19_r,temp_b1_31_19_i,temp_m2_29_17_r,temp_m2_29_17_i,temp_m2_29_19_r,temp_m2_29_19_i,temp_m2_31_17_r,temp_m2_31_17_i,temp_m2_31_19_r,temp_m2_31_19_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly497 (clk,temp_m2_29_17_r,temp_m2_29_17_i,temp_m2_29_19_r,temp_m2_29_19_i,temp_m2_31_17_r,temp_m2_31_17_i,temp_m2_31_19_r,temp_m2_31_19_i,temp_b2_29_17_r,temp_b2_29_17_i,temp_b2_29_19_r,temp_b2_29_19_i,temp_b2_31_17_r,temp_b2_31_17_i,temp_b2_31_19_r,temp_b2_31_19_i);
MULT MULT498 (clk,temp_b1_29_18_r,temp_b1_29_18_i,temp_b1_29_20_r,temp_b1_29_20_i,temp_b1_31_18_r,temp_b1_31_18_i,temp_b1_31_20_r,temp_b1_31_20_i,temp_m2_29_18_r,temp_m2_29_18_i,temp_m2_29_20_r,temp_m2_29_20_i,temp_m2_31_18_r,temp_m2_31_18_i,temp_m2_31_20_r,temp_m2_31_20_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly498 (clk,temp_m2_29_18_r,temp_m2_29_18_i,temp_m2_29_20_r,temp_m2_29_20_i,temp_m2_31_18_r,temp_m2_31_18_i,temp_m2_31_20_r,temp_m2_31_20_i,temp_b2_29_18_r,temp_b2_29_18_i,temp_b2_29_20_r,temp_b2_29_20_i,temp_b2_31_18_r,temp_b2_31_18_i,temp_b2_31_20_r,temp_b2_31_20_i);
MULT MULT499 (clk,temp_b1_30_17_r,temp_b1_30_17_i,temp_b1_30_19_r,temp_b1_30_19_i,temp_b1_32_17_r,temp_b1_32_17_i,temp_b1_32_19_r,temp_b1_32_19_i,temp_m2_30_17_r,temp_m2_30_17_i,temp_m2_30_19_r,temp_m2_30_19_i,temp_m2_32_17_r,temp_m2_32_17_i,temp_m2_32_19_r,temp_m2_32_19_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly499 (clk,temp_m2_30_17_r,temp_m2_30_17_i,temp_m2_30_19_r,temp_m2_30_19_i,temp_m2_32_17_r,temp_m2_32_17_i,temp_m2_32_19_r,temp_m2_32_19_i,temp_b2_30_17_r,temp_b2_30_17_i,temp_b2_30_19_r,temp_b2_30_19_i,temp_b2_32_17_r,temp_b2_32_17_i,temp_b2_32_19_r,temp_b2_32_19_i);
MULT MULT500 (clk,temp_b1_30_18_r,temp_b1_30_18_i,temp_b1_30_20_r,temp_b1_30_20_i,temp_b1_32_18_r,temp_b1_32_18_i,temp_b1_32_20_r,temp_b1_32_20_i,temp_m2_30_18_r,temp_m2_30_18_i,temp_m2_30_20_r,temp_m2_30_20_i,temp_m2_32_18_r,temp_m2_32_18_i,temp_m2_32_20_r,temp_m2_32_20_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly500 (clk,temp_m2_30_18_r,temp_m2_30_18_i,temp_m2_30_20_r,temp_m2_30_20_i,temp_m2_32_18_r,temp_m2_32_18_i,temp_m2_32_20_r,temp_m2_32_20_i,temp_b2_30_18_r,temp_b2_30_18_i,temp_b2_30_20_r,temp_b2_30_20_i,temp_b2_32_18_r,temp_b2_32_18_i,temp_b2_32_20_r,temp_b2_32_20_i);
MULT MULT501 (clk,temp_b1_29_21_r,temp_b1_29_21_i,temp_b1_29_23_r,temp_b1_29_23_i,temp_b1_31_21_r,temp_b1_31_21_i,temp_b1_31_23_r,temp_b1_31_23_i,temp_m2_29_21_r,temp_m2_29_21_i,temp_m2_29_23_r,temp_m2_29_23_i,temp_m2_31_21_r,temp_m2_31_21_i,temp_m2_31_23_r,temp_m2_31_23_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly501 (clk,temp_m2_29_21_r,temp_m2_29_21_i,temp_m2_29_23_r,temp_m2_29_23_i,temp_m2_31_21_r,temp_m2_31_21_i,temp_m2_31_23_r,temp_m2_31_23_i,temp_b2_29_21_r,temp_b2_29_21_i,temp_b2_29_23_r,temp_b2_29_23_i,temp_b2_31_21_r,temp_b2_31_21_i,temp_b2_31_23_r,temp_b2_31_23_i);
MULT MULT502 (clk,temp_b1_29_22_r,temp_b1_29_22_i,temp_b1_29_24_r,temp_b1_29_24_i,temp_b1_31_22_r,temp_b1_31_22_i,temp_b1_31_24_r,temp_b1_31_24_i,temp_m2_29_22_r,temp_m2_29_22_i,temp_m2_29_24_r,temp_m2_29_24_i,temp_m2_31_22_r,temp_m2_31_22_i,temp_m2_31_24_r,temp_m2_31_24_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly502 (clk,temp_m2_29_22_r,temp_m2_29_22_i,temp_m2_29_24_r,temp_m2_29_24_i,temp_m2_31_22_r,temp_m2_31_22_i,temp_m2_31_24_r,temp_m2_31_24_i,temp_b2_29_22_r,temp_b2_29_22_i,temp_b2_29_24_r,temp_b2_29_24_i,temp_b2_31_22_r,temp_b2_31_22_i,temp_b2_31_24_r,temp_b2_31_24_i);
MULT MULT503 (clk,temp_b1_30_21_r,temp_b1_30_21_i,temp_b1_30_23_r,temp_b1_30_23_i,temp_b1_32_21_r,temp_b1_32_21_i,temp_b1_32_23_r,temp_b1_32_23_i,temp_m2_30_21_r,temp_m2_30_21_i,temp_m2_30_23_r,temp_m2_30_23_i,temp_m2_32_21_r,temp_m2_32_21_i,temp_m2_32_23_r,temp_m2_32_23_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly503 (clk,temp_m2_30_21_r,temp_m2_30_21_i,temp_m2_30_23_r,temp_m2_30_23_i,temp_m2_32_21_r,temp_m2_32_21_i,temp_m2_32_23_r,temp_m2_32_23_i,temp_b2_30_21_r,temp_b2_30_21_i,temp_b2_30_23_r,temp_b2_30_23_i,temp_b2_32_21_r,temp_b2_32_21_i,temp_b2_32_23_r,temp_b2_32_23_i);
MULT MULT504 (clk,temp_b1_30_22_r,temp_b1_30_22_i,temp_b1_30_24_r,temp_b1_30_24_i,temp_b1_32_22_r,temp_b1_32_22_i,temp_b1_32_24_r,temp_b1_32_24_i,temp_m2_30_22_r,temp_m2_30_22_i,temp_m2_30_24_r,temp_m2_30_24_i,temp_m2_32_22_r,temp_m2_32_22_i,temp_m2_32_24_r,temp_m2_32_24_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly504 (clk,temp_m2_30_22_r,temp_m2_30_22_i,temp_m2_30_24_r,temp_m2_30_24_i,temp_m2_32_22_r,temp_m2_32_22_i,temp_m2_32_24_r,temp_m2_32_24_i,temp_b2_30_22_r,temp_b2_30_22_i,temp_b2_30_24_r,temp_b2_30_24_i,temp_b2_32_22_r,temp_b2_32_22_i,temp_b2_32_24_r,temp_b2_32_24_i);
MULT MULT505 (clk,temp_b1_29_25_r,temp_b1_29_25_i,temp_b1_29_27_r,temp_b1_29_27_i,temp_b1_31_25_r,temp_b1_31_25_i,temp_b1_31_27_r,temp_b1_31_27_i,temp_m2_29_25_r,temp_m2_29_25_i,temp_m2_29_27_r,temp_m2_29_27_i,temp_m2_31_25_r,temp_m2_31_25_i,temp_m2_31_27_r,temp_m2_31_27_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly505 (clk,temp_m2_29_25_r,temp_m2_29_25_i,temp_m2_29_27_r,temp_m2_29_27_i,temp_m2_31_25_r,temp_m2_31_25_i,temp_m2_31_27_r,temp_m2_31_27_i,temp_b2_29_25_r,temp_b2_29_25_i,temp_b2_29_27_r,temp_b2_29_27_i,temp_b2_31_25_r,temp_b2_31_25_i,temp_b2_31_27_r,temp_b2_31_27_i);
MULT MULT506 (clk,temp_b1_29_26_r,temp_b1_29_26_i,temp_b1_29_28_r,temp_b1_29_28_i,temp_b1_31_26_r,temp_b1_31_26_i,temp_b1_31_28_r,temp_b1_31_28_i,temp_m2_29_26_r,temp_m2_29_26_i,temp_m2_29_28_r,temp_m2_29_28_i,temp_m2_31_26_r,temp_m2_31_26_i,temp_m2_31_28_r,temp_m2_31_28_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly506 (clk,temp_m2_29_26_r,temp_m2_29_26_i,temp_m2_29_28_r,temp_m2_29_28_i,temp_m2_31_26_r,temp_m2_31_26_i,temp_m2_31_28_r,temp_m2_31_28_i,temp_b2_29_26_r,temp_b2_29_26_i,temp_b2_29_28_r,temp_b2_29_28_i,temp_b2_31_26_r,temp_b2_31_26_i,temp_b2_31_28_r,temp_b2_31_28_i);
MULT MULT507 (clk,temp_b1_30_25_r,temp_b1_30_25_i,temp_b1_30_27_r,temp_b1_30_27_i,temp_b1_32_25_r,temp_b1_32_25_i,temp_b1_32_27_r,temp_b1_32_27_i,temp_m2_30_25_r,temp_m2_30_25_i,temp_m2_30_27_r,temp_m2_30_27_i,temp_m2_32_25_r,temp_m2_32_25_i,temp_m2_32_27_r,temp_m2_32_27_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly507 (clk,temp_m2_30_25_r,temp_m2_30_25_i,temp_m2_30_27_r,temp_m2_30_27_i,temp_m2_32_25_r,temp_m2_32_25_i,temp_m2_32_27_r,temp_m2_32_27_i,temp_b2_30_25_r,temp_b2_30_25_i,temp_b2_30_27_r,temp_b2_30_27_i,temp_b2_32_25_r,temp_b2_32_25_i,temp_b2_32_27_r,temp_b2_32_27_i);
MULT MULT508 (clk,temp_b1_30_26_r,temp_b1_30_26_i,temp_b1_30_28_r,temp_b1_30_28_i,temp_b1_32_26_r,temp_b1_32_26_i,temp_b1_32_28_r,temp_b1_32_28_i,temp_m2_30_26_r,temp_m2_30_26_i,temp_m2_30_28_r,temp_m2_30_28_i,temp_m2_32_26_r,temp_m2_32_26_i,temp_m2_32_28_r,temp_m2_32_28_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly508 (clk,temp_m2_30_26_r,temp_m2_30_26_i,temp_m2_30_28_r,temp_m2_30_28_i,temp_m2_32_26_r,temp_m2_32_26_i,temp_m2_32_28_r,temp_m2_32_28_i,temp_b2_30_26_r,temp_b2_30_26_i,temp_b2_30_28_r,temp_b2_30_28_i,temp_b2_32_26_r,temp_b2_32_26_i,temp_b2_32_28_r,temp_b2_32_28_i);
MULT MULT509 (clk,temp_b1_29_29_r,temp_b1_29_29_i,temp_b1_29_31_r,temp_b1_29_31_i,temp_b1_31_29_r,temp_b1_31_29_i,temp_b1_31_31_r,temp_b1_31_31_i,temp_m2_29_29_r,temp_m2_29_29_i,temp_m2_29_31_r,temp_m2_29_31_i,temp_m2_31_29_r,temp_m2_31_29_i,temp_m2_31_31_r,temp_m2_31_31_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly509 (clk,temp_m2_29_29_r,temp_m2_29_29_i,temp_m2_29_31_r,temp_m2_29_31_i,temp_m2_31_29_r,temp_m2_31_29_i,temp_m2_31_31_r,temp_m2_31_31_i,temp_b2_29_29_r,temp_b2_29_29_i,temp_b2_29_31_r,temp_b2_29_31_i,temp_b2_31_29_r,temp_b2_31_29_i,temp_b2_31_31_r,temp_b2_31_31_i);
MULT MULT510 (clk,temp_b1_29_30_r,temp_b1_29_30_i,temp_b1_29_32_r,temp_b1_29_32_i,temp_b1_31_30_r,temp_b1_31_30_i,temp_b1_31_32_r,temp_b1_31_32_i,temp_m2_29_30_r,temp_m2_29_30_i,temp_m2_29_32_r,temp_m2_29_32_i,temp_m2_31_30_r,temp_m2_31_30_i,temp_m2_31_32_r,temp_m2_31_32_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly510 (clk,temp_m2_29_30_r,temp_m2_29_30_i,temp_m2_29_32_r,temp_m2_29_32_i,temp_m2_31_30_r,temp_m2_31_30_i,temp_m2_31_32_r,temp_m2_31_32_i,temp_b2_29_30_r,temp_b2_29_30_i,temp_b2_29_32_r,temp_b2_29_32_i,temp_b2_31_30_r,temp_b2_31_30_i,temp_b2_31_32_r,temp_b2_31_32_i);
MULT MULT511 (clk,temp_b1_30_29_r,temp_b1_30_29_i,temp_b1_30_31_r,temp_b1_30_31_i,temp_b1_32_29_r,temp_b1_32_29_i,temp_b1_32_31_r,temp_b1_32_31_i,temp_m2_30_29_r,temp_m2_30_29_i,temp_m2_30_31_r,temp_m2_30_31_i,temp_m2_32_29_r,temp_m2_32_29_i,temp_m2_32_31_r,temp_m2_32_31_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly511 (clk,temp_m2_30_29_r,temp_m2_30_29_i,temp_m2_30_31_r,temp_m2_30_31_i,temp_m2_32_29_r,temp_m2_32_29_i,temp_m2_32_31_r,temp_m2_32_31_i,temp_b2_30_29_r,temp_b2_30_29_i,temp_b2_30_31_r,temp_b2_30_31_i,temp_b2_32_29_r,temp_b2_32_29_i,temp_b2_32_31_r,temp_b2_32_31_i);
MULT MULT512 (clk,temp_b1_30_30_r,temp_b1_30_30_i,temp_b1_30_32_r,temp_b1_30_32_i,temp_b1_32_30_r,temp_b1_32_30_i,temp_b1_32_32_r,temp_b1_32_32_i,temp_m2_30_30_r,temp_m2_30_30_i,temp_m2_30_32_r,temp_m2_30_32_i,temp_m2_32_30_r,temp_m2_32_30_i,temp_m2_32_32_r,temp_m2_32_32_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly512 (clk,temp_m2_30_30_r,temp_m2_30_30_i,temp_m2_30_32_r,temp_m2_30_32_i,temp_m2_32_30_r,temp_m2_32_30_i,temp_m2_32_32_r,temp_m2_32_32_i,temp_b2_30_30_r,temp_b2_30_30_i,temp_b2_30_32_r,temp_b2_30_32_i,temp_b2_32_30_r,temp_b2_32_30_i,temp_b2_32_32_r,temp_b2_32_32_i);
MULT MULT513 (clk,temp_b2_1_1_r,temp_b2_1_1_i,temp_b2_1_5_r,temp_b2_1_5_i,temp_b2_5_1_r,temp_b2_5_1_i,temp_b2_5_5_r,temp_b2_5_5_i,temp_m3_1_1_r,temp_m3_1_1_i,temp_m3_1_5_r,temp_m3_1_5_i,temp_m3_5_1_r,temp_m3_5_1_i,temp_m3_5_5_r,temp_m3_5_5_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly513 (clk,temp_m3_1_1_r,temp_m3_1_1_i,temp_m3_1_5_r,temp_m3_1_5_i,temp_m3_5_1_r,temp_m3_5_1_i,temp_m3_5_5_r,temp_m3_5_5_i,temp_b3_1_1_r,temp_b3_1_1_i,temp_b3_1_5_r,temp_b3_1_5_i,temp_b3_5_1_r,temp_b3_5_1_i,temp_b3_5_5_r,temp_b3_5_5_i);
MULT MULT514 (clk,temp_b2_1_2_r,temp_b2_1_2_i,temp_b2_1_6_r,temp_b2_1_6_i,temp_b2_5_2_r,temp_b2_5_2_i,temp_b2_5_6_r,temp_b2_5_6_i,temp_m3_1_2_r,temp_m3_1_2_i,temp_m3_1_6_r,temp_m3_1_6_i,temp_m3_5_2_r,temp_m3_5_2_i,temp_m3_5_6_r,temp_m3_5_6_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly514 (clk,temp_m3_1_2_r,temp_m3_1_2_i,temp_m3_1_6_r,temp_m3_1_6_i,temp_m3_5_2_r,temp_m3_5_2_i,temp_m3_5_6_r,temp_m3_5_6_i,temp_b3_1_2_r,temp_b3_1_2_i,temp_b3_1_6_r,temp_b3_1_6_i,temp_b3_5_2_r,temp_b3_5_2_i,temp_b3_5_6_r,temp_b3_5_6_i);
MULT MULT515 (clk,temp_b2_1_3_r,temp_b2_1_3_i,temp_b2_1_7_r,temp_b2_1_7_i,temp_b2_5_3_r,temp_b2_5_3_i,temp_b2_5_7_r,temp_b2_5_7_i,temp_m3_1_3_r,temp_m3_1_3_i,temp_m3_1_7_r,temp_m3_1_7_i,temp_m3_5_3_r,temp_m3_5_3_i,temp_m3_5_7_r,temp_m3_5_7_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly515 (clk,temp_m3_1_3_r,temp_m3_1_3_i,temp_m3_1_7_r,temp_m3_1_7_i,temp_m3_5_3_r,temp_m3_5_3_i,temp_m3_5_7_r,temp_m3_5_7_i,temp_b3_1_3_r,temp_b3_1_3_i,temp_b3_1_7_r,temp_b3_1_7_i,temp_b3_5_3_r,temp_b3_5_3_i,temp_b3_5_7_r,temp_b3_5_7_i);
MULT MULT516 (clk,temp_b2_1_4_r,temp_b2_1_4_i,temp_b2_1_8_r,temp_b2_1_8_i,temp_b2_5_4_r,temp_b2_5_4_i,temp_b2_5_8_r,temp_b2_5_8_i,temp_m3_1_4_r,temp_m3_1_4_i,temp_m3_1_8_r,temp_m3_1_8_i,temp_m3_5_4_r,temp_m3_5_4_i,temp_m3_5_8_r,temp_m3_5_8_i,`W12_real,`W12_imag,`W0_real,`W0_imag,`W12_real,`W12_imag);
butterfly butterfly516 (clk,temp_m3_1_4_r,temp_m3_1_4_i,temp_m3_1_8_r,temp_m3_1_8_i,temp_m3_5_4_r,temp_m3_5_4_i,temp_m3_5_8_r,temp_m3_5_8_i,temp_b3_1_4_r,temp_b3_1_4_i,temp_b3_1_8_r,temp_b3_1_8_i,temp_b3_5_4_r,temp_b3_5_4_i,temp_b3_5_8_r,temp_b3_5_8_i);
MULT MULT517 (clk,temp_b2_2_1_r,temp_b2_2_1_i,temp_b2_2_5_r,temp_b2_2_5_i,temp_b2_6_1_r,temp_b2_6_1_i,temp_b2_6_5_r,temp_b2_6_5_i,temp_m3_2_1_r,temp_m3_2_1_i,temp_m3_2_5_r,temp_m3_2_5_i,temp_m3_6_1_r,temp_m3_6_1_i,temp_m3_6_5_r,temp_m3_6_5_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly517 (clk,temp_m3_2_1_r,temp_m3_2_1_i,temp_m3_2_5_r,temp_m3_2_5_i,temp_m3_6_1_r,temp_m3_6_1_i,temp_m3_6_5_r,temp_m3_6_5_i,temp_b3_2_1_r,temp_b3_2_1_i,temp_b3_2_5_r,temp_b3_2_5_i,temp_b3_6_1_r,temp_b3_6_1_i,temp_b3_6_5_r,temp_b3_6_5_i);
MULT MULT518 (clk,temp_b2_2_2_r,temp_b2_2_2_i,temp_b2_2_6_r,temp_b2_2_6_i,temp_b2_6_2_r,temp_b2_6_2_i,temp_b2_6_6_r,temp_b2_6_6_i,temp_m3_2_2_r,temp_m3_2_2_i,temp_m3_2_6_r,temp_m3_2_6_i,temp_m3_6_2_r,temp_m3_6_2_i,temp_m3_6_6_r,temp_m3_6_6_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly518 (clk,temp_m3_2_2_r,temp_m3_2_2_i,temp_m3_2_6_r,temp_m3_2_6_i,temp_m3_6_2_r,temp_m3_6_2_i,temp_m3_6_6_r,temp_m3_6_6_i,temp_b3_2_2_r,temp_b3_2_2_i,temp_b3_2_6_r,temp_b3_2_6_i,temp_b3_6_2_r,temp_b3_6_2_i,temp_b3_6_6_r,temp_b3_6_6_i);
MULT MULT519 (clk,temp_b2_2_3_r,temp_b2_2_3_i,temp_b2_2_7_r,temp_b2_2_7_i,temp_b2_6_3_r,temp_b2_6_3_i,temp_b2_6_7_r,temp_b2_6_7_i,temp_m3_2_3_r,temp_m3_2_3_i,temp_m3_2_7_r,temp_m3_2_7_i,temp_m3_6_3_r,temp_m3_6_3_i,temp_m3_6_7_r,temp_m3_6_7_i,`W8_real,`W8_imag,`W4_real,`W4_imag,`W12_real,`W12_imag);
butterfly butterfly519 (clk,temp_m3_2_3_r,temp_m3_2_3_i,temp_m3_2_7_r,temp_m3_2_7_i,temp_m3_6_3_r,temp_m3_6_3_i,temp_m3_6_7_r,temp_m3_6_7_i,temp_b3_2_3_r,temp_b3_2_3_i,temp_b3_2_7_r,temp_b3_2_7_i,temp_b3_6_3_r,temp_b3_6_3_i,temp_b3_6_7_r,temp_b3_6_7_i);
MULT MULT520 (clk,temp_b2_2_4_r,temp_b2_2_4_i,temp_b2_2_8_r,temp_b2_2_8_i,temp_b2_6_4_r,temp_b2_6_4_i,temp_b2_6_8_r,temp_b2_6_8_i,temp_m3_2_4_r,temp_m3_2_4_i,temp_m3_2_8_r,temp_m3_2_8_i,temp_m3_6_4_r,temp_m3_6_4_i,temp_m3_6_8_r,temp_m3_6_8_i,`W12_real,`W12_imag,`W4_real,`W4_imag,`W16_real,`W16_imag);
butterfly butterfly520 (clk,temp_m3_2_4_r,temp_m3_2_4_i,temp_m3_2_8_r,temp_m3_2_8_i,temp_m3_6_4_r,temp_m3_6_4_i,temp_m3_6_8_r,temp_m3_6_8_i,temp_b3_2_4_r,temp_b3_2_4_i,temp_b3_2_8_r,temp_b3_2_8_i,temp_b3_6_4_r,temp_b3_6_4_i,temp_b3_6_8_r,temp_b3_6_8_i);
MULT MULT521 (clk,temp_b2_3_1_r,temp_b2_3_1_i,temp_b2_3_5_r,temp_b2_3_5_i,temp_b2_7_1_r,temp_b2_7_1_i,temp_b2_7_5_r,temp_b2_7_5_i,temp_m3_3_1_r,temp_m3_3_1_i,temp_m3_3_5_r,temp_m3_3_5_i,temp_m3_7_1_r,temp_m3_7_1_i,temp_m3_7_5_r,temp_m3_7_5_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly521 (clk,temp_m3_3_1_r,temp_m3_3_1_i,temp_m3_3_5_r,temp_m3_3_5_i,temp_m3_7_1_r,temp_m3_7_1_i,temp_m3_7_5_r,temp_m3_7_5_i,temp_b3_3_1_r,temp_b3_3_1_i,temp_b3_3_5_r,temp_b3_3_5_i,temp_b3_7_1_r,temp_b3_7_1_i,temp_b3_7_5_r,temp_b3_7_5_i);
MULT MULT522 (clk,temp_b2_3_2_r,temp_b2_3_2_i,temp_b2_3_6_r,temp_b2_3_6_i,temp_b2_7_2_r,temp_b2_7_2_i,temp_b2_7_6_r,temp_b2_7_6_i,temp_m3_3_2_r,temp_m3_3_2_i,temp_m3_3_6_r,temp_m3_3_6_i,temp_m3_7_2_r,temp_m3_7_2_i,temp_m3_7_6_r,temp_m3_7_6_i,`W4_real,`W4_imag,`W8_real,`W8_imag,`W12_real,`W12_imag);
butterfly butterfly522 (clk,temp_m3_3_2_r,temp_m3_3_2_i,temp_m3_3_6_r,temp_m3_3_6_i,temp_m3_7_2_r,temp_m3_7_2_i,temp_m3_7_6_r,temp_m3_7_6_i,temp_b3_3_2_r,temp_b3_3_2_i,temp_b3_3_6_r,temp_b3_3_6_i,temp_b3_7_2_r,temp_b3_7_2_i,temp_b3_7_6_r,temp_b3_7_6_i);
MULT MULT523 (clk,temp_b2_3_3_r,temp_b2_3_3_i,temp_b2_3_7_r,temp_b2_3_7_i,temp_b2_7_3_r,temp_b2_7_3_i,temp_b2_7_7_r,temp_b2_7_7_i,temp_m3_3_3_r,temp_m3_3_3_i,temp_m3_3_7_r,temp_m3_3_7_i,temp_m3_7_3_r,temp_m3_7_3_i,temp_m3_7_7_r,temp_m3_7_7_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly523 (clk,temp_m3_3_3_r,temp_m3_3_3_i,temp_m3_3_7_r,temp_m3_3_7_i,temp_m3_7_3_r,temp_m3_7_3_i,temp_m3_7_7_r,temp_m3_7_7_i,temp_b3_3_3_r,temp_b3_3_3_i,temp_b3_3_7_r,temp_b3_3_7_i,temp_b3_7_3_r,temp_b3_7_3_i,temp_b3_7_7_r,temp_b3_7_7_i);
MULT MULT524 (clk,temp_b2_3_4_r,temp_b2_3_4_i,temp_b2_3_8_r,temp_b2_3_8_i,temp_b2_7_4_r,temp_b2_7_4_i,temp_b2_7_8_r,temp_b2_7_8_i,temp_m3_3_4_r,temp_m3_3_4_i,temp_m3_3_8_r,temp_m3_3_8_i,temp_m3_7_4_r,temp_m3_7_4_i,temp_m3_7_8_r,temp_m3_7_8_i,`W12_real,`W12_imag,`W8_real,`W8_imag,`W20_real,`W20_imag);
butterfly butterfly524 (clk,temp_m3_3_4_r,temp_m3_3_4_i,temp_m3_3_8_r,temp_m3_3_8_i,temp_m3_7_4_r,temp_m3_7_4_i,temp_m3_7_8_r,temp_m3_7_8_i,temp_b3_3_4_r,temp_b3_3_4_i,temp_b3_3_8_r,temp_b3_3_8_i,temp_b3_7_4_r,temp_b3_7_4_i,temp_b3_7_8_r,temp_b3_7_8_i);
MULT MULT525 (clk,temp_b2_4_1_r,temp_b2_4_1_i,temp_b2_4_5_r,temp_b2_4_5_i,temp_b2_8_1_r,temp_b2_8_1_i,temp_b2_8_5_r,temp_b2_8_5_i,temp_m3_4_1_r,temp_m3_4_1_i,temp_m3_4_5_r,temp_m3_4_5_i,temp_m3_8_1_r,temp_m3_8_1_i,temp_m3_8_5_r,temp_m3_8_5_i,`W0_real,`W0_imag,`W12_real,`W12_imag,`W12_real,`W12_imag);
butterfly butterfly525 (clk,temp_m3_4_1_r,temp_m3_4_1_i,temp_m3_4_5_r,temp_m3_4_5_i,temp_m3_8_1_r,temp_m3_8_1_i,temp_m3_8_5_r,temp_m3_8_5_i,temp_b3_4_1_r,temp_b3_4_1_i,temp_b3_4_5_r,temp_b3_4_5_i,temp_b3_8_1_r,temp_b3_8_1_i,temp_b3_8_5_r,temp_b3_8_5_i);
MULT MULT526 (clk,temp_b2_4_2_r,temp_b2_4_2_i,temp_b2_4_6_r,temp_b2_4_6_i,temp_b2_8_2_r,temp_b2_8_2_i,temp_b2_8_6_r,temp_b2_8_6_i,temp_m3_4_2_r,temp_m3_4_2_i,temp_m3_4_6_r,temp_m3_4_6_i,temp_m3_8_2_r,temp_m3_8_2_i,temp_m3_8_6_r,temp_m3_8_6_i,`W4_real,`W4_imag,`W12_real,`W12_imag,`W16_real,`W16_imag);
butterfly butterfly526 (clk,temp_m3_4_2_r,temp_m3_4_2_i,temp_m3_4_6_r,temp_m3_4_6_i,temp_m3_8_2_r,temp_m3_8_2_i,temp_m3_8_6_r,temp_m3_8_6_i,temp_b3_4_2_r,temp_b3_4_2_i,temp_b3_4_6_r,temp_b3_4_6_i,temp_b3_8_2_r,temp_b3_8_2_i,temp_b3_8_6_r,temp_b3_8_6_i);
MULT MULT527 (clk,temp_b2_4_3_r,temp_b2_4_3_i,temp_b2_4_7_r,temp_b2_4_7_i,temp_b2_8_3_r,temp_b2_8_3_i,temp_b2_8_7_r,temp_b2_8_7_i,temp_m3_4_3_r,temp_m3_4_3_i,temp_m3_4_7_r,temp_m3_4_7_i,temp_m3_8_3_r,temp_m3_8_3_i,temp_m3_8_7_r,temp_m3_8_7_i,`W8_real,`W8_imag,`W12_real,`W12_imag,`W20_real,`W20_imag);
butterfly butterfly527 (clk,temp_m3_4_3_r,temp_m3_4_3_i,temp_m3_4_7_r,temp_m3_4_7_i,temp_m3_8_3_r,temp_m3_8_3_i,temp_m3_8_7_r,temp_m3_8_7_i,temp_b3_4_3_r,temp_b3_4_3_i,temp_b3_4_7_r,temp_b3_4_7_i,temp_b3_8_3_r,temp_b3_8_3_i,temp_b3_8_7_r,temp_b3_8_7_i);
MULT MULT528 (clk,temp_b2_4_4_r,temp_b2_4_4_i,temp_b2_4_8_r,temp_b2_4_8_i,temp_b2_8_4_r,temp_b2_8_4_i,temp_b2_8_8_r,temp_b2_8_8_i,temp_m3_4_4_r,temp_m3_4_4_i,temp_m3_4_8_r,temp_m3_4_8_i,temp_m3_8_4_r,temp_m3_8_4_i,temp_m3_8_8_r,temp_m3_8_8_i,`W12_real,`W12_imag,`W12_real,`W12_imag,`W24_real,`W24_imag);
butterfly butterfly528 (clk,temp_m3_4_4_r,temp_m3_4_4_i,temp_m3_4_8_r,temp_m3_4_8_i,temp_m3_8_4_r,temp_m3_8_4_i,temp_m3_8_8_r,temp_m3_8_8_i,temp_b3_4_4_r,temp_b3_4_4_i,temp_b3_4_8_r,temp_b3_4_8_i,temp_b3_8_4_r,temp_b3_8_4_i,temp_b3_8_8_r,temp_b3_8_8_i);
MULT MULT529 (clk,temp_b2_1_9_r,temp_b2_1_9_i,temp_b2_1_13_r,temp_b2_1_13_i,temp_b2_5_9_r,temp_b2_5_9_i,temp_b2_5_13_r,temp_b2_5_13_i,temp_m3_1_9_r,temp_m3_1_9_i,temp_m3_1_13_r,temp_m3_1_13_i,temp_m3_5_9_r,temp_m3_5_9_i,temp_m3_5_13_r,temp_m3_5_13_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly529 (clk,temp_m3_1_9_r,temp_m3_1_9_i,temp_m3_1_13_r,temp_m3_1_13_i,temp_m3_5_9_r,temp_m3_5_9_i,temp_m3_5_13_r,temp_m3_5_13_i,temp_b3_1_9_r,temp_b3_1_9_i,temp_b3_1_13_r,temp_b3_1_13_i,temp_b3_5_9_r,temp_b3_5_9_i,temp_b3_5_13_r,temp_b3_5_13_i);
MULT MULT530 (clk,temp_b2_1_10_r,temp_b2_1_10_i,temp_b2_1_14_r,temp_b2_1_14_i,temp_b2_5_10_r,temp_b2_5_10_i,temp_b2_5_14_r,temp_b2_5_14_i,temp_m3_1_10_r,temp_m3_1_10_i,temp_m3_1_14_r,temp_m3_1_14_i,temp_m3_5_10_r,temp_m3_5_10_i,temp_m3_5_14_r,temp_m3_5_14_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly530 (clk,temp_m3_1_10_r,temp_m3_1_10_i,temp_m3_1_14_r,temp_m3_1_14_i,temp_m3_5_10_r,temp_m3_5_10_i,temp_m3_5_14_r,temp_m3_5_14_i,temp_b3_1_10_r,temp_b3_1_10_i,temp_b3_1_14_r,temp_b3_1_14_i,temp_b3_5_10_r,temp_b3_5_10_i,temp_b3_5_14_r,temp_b3_5_14_i);
MULT MULT531 (clk,temp_b2_1_11_r,temp_b2_1_11_i,temp_b2_1_15_r,temp_b2_1_15_i,temp_b2_5_11_r,temp_b2_5_11_i,temp_b2_5_15_r,temp_b2_5_15_i,temp_m3_1_11_r,temp_m3_1_11_i,temp_m3_1_15_r,temp_m3_1_15_i,temp_m3_5_11_r,temp_m3_5_11_i,temp_m3_5_15_r,temp_m3_5_15_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly531 (clk,temp_m3_1_11_r,temp_m3_1_11_i,temp_m3_1_15_r,temp_m3_1_15_i,temp_m3_5_11_r,temp_m3_5_11_i,temp_m3_5_15_r,temp_m3_5_15_i,temp_b3_1_11_r,temp_b3_1_11_i,temp_b3_1_15_r,temp_b3_1_15_i,temp_b3_5_11_r,temp_b3_5_11_i,temp_b3_5_15_r,temp_b3_5_15_i);
MULT MULT532 (clk,temp_b2_1_12_r,temp_b2_1_12_i,temp_b2_1_16_r,temp_b2_1_16_i,temp_b2_5_12_r,temp_b2_5_12_i,temp_b2_5_16_r,temp_b2_5_16_i,temp_m3_1_12_r,temp_m3_1_12_i,temp_m3_1_16_r,temp_m3_1_16_i,temp_m3_5_12_r,temp_m3_5_12_i,temp_m3_5_16_r,temp_m3_5_16_i,`W12_real,`W12_imag,`W0_real,`W0_imag,`W12_real,`W12_imag);
butterfly butterfly532 (clk,temp_m3_1_12_r,temp_m3_1_12_i,temp_m3_1_16_r,temp_m3_1_16_i,temp_m3_5_12_r,temp_m3_5_12_i,temp_m3_5_16_r,temp_m3_5_16_i,temp_b3_1_12_r,temp_b3_1_12_i,temp_b3_1_16_r,temp_b3_1_16_i,temp_b3_5_12_r,temp_b3_5_12_i,temp_b3_5_16_r,temp_b3_5_16_i);
MULT MULT533 (clk,temp_b2_2_9_r,temp_b2_2_9_i,temp_b2_2_13_r,temp_b2_2_13_i,temp_b2_6_9_r,temp_b2_6_9_i,temp_b2_6_13_r,temp_b2_6_13_i,temp_m3_2_9_r,temp_m3_2_9_i,temp_m3_2_13_r,temp_m3_2_13_i,temp_m3_6_9_r,temp_m3_6_9_i,temp_m3_6_13_r,temp_m3_6_13_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly533 (clk,temp_m3_2_9_r,temp_m3_2_9_i,temp_m3_2_13_r,temp_m3_2_13_i,temp_m3_6_9_r,temp_m3_6_9_i,temp_m3_6_13_r,temp_m3_6_13_i,temp_b3_2_9_r,temp_b3_2_9_i,temp_b3_2_13_r,temp_b3_2_13_i,temp_b3_6_9_r,temp_b3_6_9_i,temp_b3_6_13_r,temp_b3_6_13_i);
MULT MULT534 (clk,temp_b2_2_10_r,temp_b2_2_10_i,temp_b2_2_14_r,temp_b2_2_14_i,temp_b2_6_10_r,temp_b2_6_10_i,temp_b2_6_14_r,temp_b2_6_14_i,temp_m3_2_10_r,temp_m3_2_10_i,temp_m3_2_14_r,temp_m3_2_14_i,temp_m3_6_10_r,temp_m3_6_10_i,temp_m3_6_14_r,temp_m3_6_14_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly534 (clk,temp_m3_2_10_r,temp_m3_2_10_i,temp_m3_2_14_r,temp_m3_2_14_i,temp_m3_6_10_r,temp_m3_6_10_i,temp_m3_6_14_r,temp_m3_6_14_i,temp_b3_2_10_r,temp_b3_2_10_i,temp_b3_2_14_r,temp_b3_2_14_i,temp_b3_6_10_r,temp_b3_6_10_i,temp_b3_6_14_r,temp_b3_6_14_i);
MULT MULT535 (clk,temp_b2_2_11_r,temp_b2_2_11_i,temp_b2_2_15_r,temp_b2_2_15_i,temp_b2_6_11_r,temp_b2_6_11_i,temp_b2_6_15_r,temp_b2_6_15_i,temp_m3_2_11_r,temp_m3_2_11_i,temp_m3_2_15_r,temp_m3_2_15_i,temp_m3_6_11_r,temp_m3_6_11_i,temp_m3_6_15_r,temp_m3_6_15_i,`W8_real,`W8_imag,`W4_real,`W4_imag,`W12_real,`W12_imag);
butterfly butterfly535 (clk,temp_m3_2_11_r,temp_m3_2_11_i,temp_m3_2_15_r,temp_m3_2_15_i,temp_m3_6_11_r,temp_m3_6_11_i,temp_m3_6_15_r,temp_m3_6_15_i,temp_b3_2_11_r,temp_b3_2_11_i,temp_b3_2_15_r,temp_b3_2_15_i,temp_b3_6_11_r,temp_b3_6_11_i,temp_b3_6_15_r,temp_b3_6_15_i);
MULT MULT536 (clk,temp_b2_2_12_r,temp_b2_2_12_i,temp_b2_2_16_r,temp_b2_2_16_i,temp_b2_6_12_r,temp_b2_6_12_i,temp_b2_6_16_r,temp_b2_6_16_i,temp_m3_2_12_r,temp_m3_2_12_i,temp_m3_2_16_r,temp_m3_2_16_i,temp_m3_6_12_r,temp_m3_6_12_i,temp_m3_6_16_r,temp_m3_6_16_i,`W12_real,`W12_imag,`W4_real,`W4_imag,`W16_real,`W16_imag);
butterfly butterfly536 (clk,temp_m3_2_12_r,temp_m3_2_12_i,temp_m3_2_16_r,temp_m3_2_16_i,temp_m3_6_12_r,temp_m3_6_12_i,temp_m3_6_16_r,temp_m3_6_16_i,temp_b3_2_12_r,temp_b3_2_12_i,temp_b3_2_16_r,temp_b3_2_16_i,temp_b3_6_12_r,temp_b3_6_12_i,temp_b3_6_16_r,temp_b3_6_16_i);
MULT MULT537 (clk,temp_b2_3_9_r,temp_b2_3_9_i,temp_b2_3_13_r,temp_b2_3_13_i,temp_b2_7_9_r,temp_b2_7_9_i,temp_b2_7_13_r,temp_b2_7_13_i,temp_m3_3_9_r,temp_m3_3_9_i,temp_m3_3_13_r,temp_m3_3_13_i,temp_m3_7_9_r,temp_m3_7_9_i,temp_m3_7_13_r,temp_m3_7_13_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly537 (clk,temp_m3_3_9_r,temp_m3_3_9_i,temp_m3_3_13_r,temp_m3_3_13_i,temp_m3_7_9_r,temp_m3_7_9_i,temp_m3_7_13_r,temp_m3_7_13_i,temp_b3_3_9_r,temp_b3_3_9_i,temp_b3_3_13_r,temp_b3_3_13_i,temp_b3_7_9_r,temp_b3_7_9_i,temp_b3_7_13_r,temp_b3_7_13_i);
MULT MULT538 (clk,temp_b2_3_10_r,temp_b2_3_10_i,temp_b2_3_14_r,temp_b2_3_14_i,temp_b2_7_10_r,temp_b2_7_10_i,temp_b2_7_14_r,temp_b2_7_14_i,temp_m3_3_10_r,temp_m3_3_10_i,temp_m3_3_14_r,temp_m3_3_14_i,temp_m3_7_10_r,temp_m3_7_10_i,temp_m3_7_14_r,temp_m3_7_14_i,`W4_real,`W4_imag,`W8_real,`W8_imag,`W12_real,`W12_imag);
butterfly butterfly538 (clk,temp_m3_3_10_r,temp_m3_3_10_i,temp_m3_3_14_r,temp_m3_3_14_i,temp_m3_7_10_r,temp_m3_7_10_i,temp_m3_7_14_r,temp_m3_7_14_i,temp_b3_3_10_r,temp_b3_3_10_i,temp_b3_3_14_r,temp_b3_3_14_i,temp_b3_7_10_r,temp_b3_7_10_i,temp_b3_7_14_r,temp_b3_7_14_i);
MULT MULT539 (clk,temp_b2_3_11_r,temp_b2_3_11_i,temp_b2_3_15_r,temp_b2_3_15_i,temp_b2_7_11_r,temp_b2_7_11_i,temp_b2_7_15_r,temp_b2_7_15_i,temp_m3_3_11_r,temp_m3_3_11_i,temp_m3_3_15_r,temp_m3_3_15_i,temp_m3_7_11_r,temp_m3_7_11_i,temp_m3_7_15_r,temp_m3_7_15_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly539 (clk,temp_m3_3_11_r,temp_m3_3_11_i,temp_m3_3_15_r,temp_m3_3_15_i,temp_m3_7_11_r,temp_m3_7_11_i,temp_m3_7_15_r,temp_m3_7_15_i,temp_b3_3_11_r,temp_b3_3_11_i,temp_b3_3_15_r,temp_b3_3_15_i,temp_b3_7_11_r,temp_b3_7_11_i,temp_b3_7_15_r,temp_b3_7_15_i);
MULT MULT540 (clk,temp_b2_3_12_r,temp_b2_3_12_i,temp_b2_3_16_r,temp_b2_3_16_i,temp_b2_7_12_r,temp_b2_7_12_i,temp_b2_7_16_r,temp_b2_7_16_i,temp_m3_3_12_r,temp_m3_3_12_i,temp_m3_3_16_r,temp_m3_3_16_i,temp_m3_7_12_r,temp_m3_7_12_i,temp_m3_7_16_r,temp_m3_7_16_i,`W12_real,`W12_imag,`W8_real,`W8_imag,`W20_real,`W20_imag);
butterfly butterfly540 (clk,temp_m3_3_12_r,temp_m3_3_12_i,temp_m3_3_16_r,temp_m3_3_16_i,temp_m3_7_12_r,temp_m3_7_12_i,temp_m3_7_16_r,temp_m3_7_16_i,temp_b3_3_12_r,temp_b3_3_12_i,temp_b3_3_16_r,temp_b3_3_16_i,temp_b3_7_12_r,temp_b3_7_12_i,temp_b3_7_16_r,temp_b3_7_16_i);
MULT MULT541 (clk,temp_b2_4_9_r,temp_b2_4_9_i,temp_b2_4_13_r,temp_b2_4_13_i,temp_b2_8_9_r,temp_b2_8_9_i,temp_b2_8_13_r,temp_b2_8_13_i,temp_m3_4_9_r,temp_m3_4_9_i,temp_m3_4_13_r,temp_m3_4_13_i,temp_m3_8_9_r,temp_m3_8_9_i,temp_m3_8_13_r,temp_m3_8_13_i,`W0_real,`W0_imag,`W12_real,`W12_imag,`W12_real,`W12_imag);
butterfly butterfly541 (clk,temp_m3_4_9_r,temp_m3_4_9_i,temp_m3_4_13_r,temp_m3_4_13_i,temp_m3_8_9_r,temp_m3_8_9_i,temp_m3_8_13_r,temp_m3_8_13_i,temp_b3_4_9_r,temp_b3_4_9_i,temp_b3_4_13_r,temp_b3_4_13_i,temp_b3_8_9_r,temp_b3_8_9_i,temp_b3_8_13_r,temp_b3_8_13_i);
MULT MULT542 (clk,temp_b2_4_10_r,temp_b2_4_10_i,temp_b2_4_14_r,temp_b2_4_14_i,temp_b2_8_10_r,temp_b2_8_10_i,temp_b2_8_14_r,temp_b2_8_14_i,temp_m3_4_10_r,temp_m3_4_10_i,temp_m3_4_14_r,temp_m3_4_14_i,temp_m3_8_10_r,temp_m3_8_10_i,temp_m3_8_14_r,temp_m3_8_14_i,`W4_real,`W4_imag,`W12_real,`W12_imag,`W16_real,`W16_imag);
butterfly butterfly542 (clk,temp_m3_4_10_r,temp_m3_4_10_i,temp_m3_4_14_r,temp_m3_4_14_i,temp_m3_8_10_r,temp_m3_8_10_i,temp_m3_8_14_r,temp_m3_8_14_i,temp_b3_4_10_r,temp_b3_4_10_i,temp_b3_4_14_r,temp_b3_4_14_i,temp_b3_8_10_r,temp_b3_8_10_i,temp_b3_8_14_r,temp_b3_8_14_i);
MULT MULT543 (clk,temp_b2_4_11_r,temp_b2_4_11_i,temp_b2_4_15_r,temp_b2_4_15_i,temp_b2_8_11_r,temp_b2_8_11_i,temp_b2_8_15_r,temp_b2_8_15_i,temp_m3_4_11_r,temp_m3_4_11_i,temp_m3_4_15_r,temp_m3_4_15_i,temp_m3_8_11_r,temp_m3_8_11_i,temp_m3_8_15_r,temp_m3_8_15_i,`W8_real,`W8_imag,`W12_real,`W12_imag,`W20_real,`W20_imag);
butterfly butterfly543 (clk,temp_m3_4_11_r,temp_m3_4_11_i,temp_m3_4_15_r,temp_m3_4_15_i,temp_m3_8_11_r,temp_m3_8_11_i,temp_m3_8_15_r,temp_m3_8_15_i,temp_b3_4_11_r,temp_b3_4_11_i,temp_b3_4_15_r,temp_b3_4_15_i,temp_b3_8_11_r,temp_b3_8_11_i,temp_b3_8_15_r,temp_b3_8_15_i);
MULT MULT544 (clk,temp_b2_4_12_r,temp_b2_4_12_i,temp_b2_4_16_r,temp_b2_4_16_i,temp_b2_8_12_r,temp_b2_8_12_i,temp_b2_8_16_r,temp_b2_8_16_i,temp_m3_4_12_r,temp_m3_4_12_i,temp_m3_4_16_r,temp_m3_4_16_i,temp_m3_8_12_r,temp_m3_8_12_i,temp_m3_8_16_r,temp_m3_8_16_i,`W12_real,`W12_imag,`W12_real,`W12_imag,`W24_real,`W24_imag);
butterfly butterfly544 (clk,temp_m3_4_12_r,temp_m3_4_12_i,temp_m3_4_16_r,temp_m3_4_16_i,temp_m3_8_12_r,temp_m3_8_12_i,temp_m3_8_16_r,temp_m3_8_16_i,temp_b3_4_12_r,temp_b3_4_12_i,temp_b3_4_16_r,temp_b3_4_16_i,temp_b3_8_12_r,temp_b3_8_12_i,temp_b3_8_16_r,temp_b3_8_16_i);
MULT MULT545 (clk,temp_b2_1_17_r,temp_b2_1_17_i,temp_b2_1_21_r,temp_b2_1_21_i,temp_b2_5_17_r,temp_b2_5_17_i,temp_b2_5_21_r,temp_b2_5_21_i,temp_m3_1_17_r,temp_m3_1_17_i,temp_m3_1_21_r,temp_m3_1_21_i,temp_m3_5_17_r,temp_m3_5_17_i,temp_m3_5_21_r,temp_m3_5_21_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly545 (clk,temp_m3_1_17_r,temp_m3_1_17_i,temp_m3_1_21_r,temp_m3_1_21_i,temp_m3_5_17_r,temp_m3_5_17_i,temp_m3_5_21_r,temp_m3_5_21_i,temp_b3_1_17_r,temp_b3_1_17_i,temp_b3_1_21_r,temp_b3_1_21_i,temp_b3_5_17_r,temp_b3_5_17_i,temp_b3_5_21_r,temp_b3_5_21_i);
MULT MULT546 (clk,temp_b2_1_18_r,temp_b2_1_18_i,temp_b2_1_22_r,temp_b2_1_22_i,temp_b2_5_18_r,temp_b2_5_18_i,temp_b2_5_22_r,temp_b2_5_22_i,temp_m3_1_18_r,temp_m3_1_18_i,temp_m3_1_22_r,temp_m3_1_22_i,temp_m3_5_18_r,temp_m3_5_18_i,temp_m3_5_22_r,temp_m3_5_22_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly546 (clk,temp_m3_1_18_r,temp_m3_1_18_i,temp_m3_1_22_r,temp_m3_1_22_i,temp_m3_5_18_r,temp_m3_5_18_i,temp_m3_5_22_r,temp_m3_5_22_i,temp_b3_1_18_r,temp_b3_1_18_i,temp_b3_1_22_r,temp_b3_1_22_i,temp_b3_5_18_r,temp_b3_5_18_i,temp_b3_5_22_r,temp_b3_5_22_i);
MULT MULT547 (clk,temp_b2_1_19_r,temp_b2_1_19_i,temp_b2_1_23_r,temp_b2_1_23_i,temp_b2_5_19_r,temp_b2_5_19_i,temp_b2_5_23_r,temp_b2_5_23_i,temp_m3_1_19_r,temp_m3_1_19_i,temp_m3_1_23_r,temp_m3_1_23_i,temp_m3_5_19_r,temp_m3_5_19_i,temp_m3_5_23_r,temp_m3_5_23_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly547 (clk,temp_m3_1_19_r,temp_m3_1_19_i,temp_m3_1_23_r,temp_m3_1_23_i,temp_m3_5_19_r,temp_m3_5_19_i,temp_m3_5_23_r,temp_m3_5_23_i,temp_b3_1_19_r,temp_b3_1_19_i,temp_b3_1_23_r,temp_b3_1_23_i,temp_b3_5_19_r,temp_b3_5_19_i,temp_b3_5_23_r,temp_b3_5_23_i);
MULT MULT548 (clk,temp_b2_1_20_r,temp_b2_1_20_i,temp_b2_1_24_r,temp_b2_1_24_i,temp_b2_5_20_r,temp_b2_5_20_i,temp_b2_5_24_r,temp_b2_5_24_i,temp_m3_1_20_r,temp_m3_1_20_i,temp_m3_1_24_r,temp_m3_1_24_i,temp_m3_5_20_r,temp_m3_5_20_i,temp_m3_5_24_r,temp_m3_5_24_i,`W12_real,`W12_imag,`W0_real,`W0_imag,`W12_real,`W12_imag);
butterfly butterfly548 (clk,temp_m3_1_20_r,temp_m3_1_20_i,temp_m3_1_24_r,temp_m3_1_24_i,temp_m3_5_20_r,temp_m3_5_20_i,temp_m3_5_24_r,temp_m3_5_24_i,temp_b3_1_20_r,temp_b3_1_20_i,temp_b3_1_24_r,temp_b3_1_24_i,temp_b3_5_20_r,temp_b3_5_20_i,temp_b3_5_24_r,temp_b3_5_24_i);
MULT MULT549 (clk,temp_b2_2_17_r,temp_b2_2_17_i,temp_b2_2_21_r,temp_b2_2_21_i,temp_b2_6_17_r,temp_b2_6_17_i,temp_b2_6_21_r,temp_b2_6_21_i,temp_m3_2_17_r,temp_m3_2_17_i,temp_m3_2_21_r,temp_m3_2_21_i,temp_m3_6_17_r,temp_m3_6_17_i,temp_m3_6_21_r,temp_m3_6_21_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly549 (clk,temp_m3_2_17_r,temp_m3_2_17_i,temp_m3_2_21_r,temp_m3_2_21_i,temp_m3_6_17_r,temp_m3_6_17_i,temp_m3_6_21_r,temp_m3_6_21_i,temp_b3_2_17_r,temp_b3_2_17_i,temp_b3_2_21_r,temp_b3_2_21_i,temp_b3_6_17_r,temp_b3_6_17_i,temp_b3_6_21_r,temp_b3_6_21_i);
MULT MULT550 (clk,temp_b2_2_18_r,temp_b2_2_18_i,temp_b2_2_22_r,temp_b2_2_22_i,temp_b2_6_18_r,temp_b2_6_18_i,temp_b2_6_22_r,temp_b2_6_22_i,temp_m3_2_18_r,temp_m3_2_18_i,temp_m3_2_22_r,temp_m3_2_22_i,temp_m3_6_18_r,temp_m3_6_18_i,temp_m3_6_22_r,temp_m3_6_22_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly550 (clk,temp_m3_2_18_r,temp_m3_2_18_i,temp_m3_2_22_r,temp_m3_2_22_i,temp_m3_6_18_r,temp_m3_6_18_i,temp_m3_6_22_r,temp_m3_6_22_i,temp_b3_2_18_r,temp_b3_2_18_i,temp_b3_2_22_r,temp_b3_2_22_i,temp_b3_6_18_r,temp_b3_6_18_i,temp_b3_6_22_r,temp_b3_6_22_i);
MULT MULT551 (clk,temp_b2_2_19_r,temp_b2_2_19_i,temp_b2_2_23_r,temp_b2_2_23_i,temp_b2_6_19_r,temp_b2_6_19_i,temp_b2_6_23_r,temp_b2_6_23_i,temp_m3_2_19_r,temp_m3_2_19_i,temp_m3_2_23_r,temp_m3_2_23_i,temp_m3_6_19_r,temp_m3_6_19_i,temp_m3_6_23_r,temp_m3_6_23_i,`W8_real,`W8_imag,`W4_real,`W4_imag,`W12_real,`W12_imag);
butterfly butterfly551 (clk,temp_m3_2_19_r,temp_m3_2_19_i,temp_m3_2_23_r,temp_m3_2_23_i,temp_m3_6_19_r,temp_m3_6_19_i,temp_m3_6_23_r,temp_m3_6_23_i,temp_b3_2_19_r,temp_b3_2_19_i,temp_b3_2_23_r,temp_b3_2_23_i,temp_b3_6_19_r,temp_b3_6_19_i,temp_b3_6_23_r,temp_b3_6_23_i);
MULT MULT552 (clk,temp_b2_2_20_r,temp_b2_2_20_i,temp_b2_2_24_r,temp_b2_2_24_i,temp_b2_6_20_r,temp_b2_6_20_i,temp_b2_6_24_r,temp_b2_6_24_i,temp_m3_2_20_r,temp_m3_2_20_i,temp_m3_2_24_r,temp_m3_2_24_i,temp_m3_6_20_r,temp_m3_6_20_i,temp_m3_6_24_r,temp_m3_6_24_i,`W12_real,`W12_imag,`W4_real,`W4_imag,`W16_real,`W16_imag);
butterfly butterfly552 (clk,temp_m3_2_20_r,temp_m3_2_20_i,temp_m3_2_24_r,temp_m3_2_24_i,temp_m3_6_20_r,temp_m3_6_20_i,temp_m3_6_24_r,temp_m3_6_24_i,temp_b3_2_20_r,temp_b3_2_20_i,temp_b3_2_24_r,temp_b3_2_24_i,temp_b3_6_20_r,temp_b3_6_20_i,temp_b3_6_24_r,temp_b3_6_24_i);
MULT MULT553 (clk,temp_b2_3_17_r,temp_b2_3_17_i,temp_b2_3_21_r,temp_b2_3_21_i,temp_b2_7_17_r,temp_b2_7_17_i,temp_b2_7_21_r,temp_b2_7_21_i,temp_m3_3_17_r,temp_m3_3_17_i,temp_m3_3_21_r,temp_m3_3_21_i,temp_m3_7_17_r,temp_m3_7_17_i,temp_m3_7_21_r,temp_m3_7_21_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly553 (clk,temp_m3_3_17_r,temp_m3_3_17_i,temp_m3_3_21_r,temp_m3_3_21_i,temp_m3_7_17_r,temp_m3_7_17_i,temp_m3_7_21_r,temp_m3_7_21_i,temp_b3_3_17_r,temp_b3_3_17_i,temp_b3_3_21_r,temp_b3_3_21_i,temp_b3_7_17_r,temp_b3_7_17_i,temp_b3_7_21_r,temp_b3_7_21_i);
MULT MULT554 (clk,temp_b2_3_18_r,temp_b2_3_18_i,temp_b2_3_22_r,temp_b2_3_22_i,temp_b2_7_18_r,temp_b2_7_18_i,temp_b2_7_22_r,temp_b2_7_22_i,temp_m3_3_18_r,temp_m3_3_18_i,temp_m3_3_22_r,temp_m3_3_22_i,temp_m3_7_18_r,temp_m3_7_18_i,temp_m3_7_22_r,temp_m3_7_22_i,`W4_real,`W4_imag,`W8_real,`W8_imag,`W12_real,`W12_imag);
butterfly butterfly554 (clk,temp_m3_3_18_r,temp_m3_3_18_i,temp_m3_3_22_r,temp_m3_3_22_i,temp_m3_7_18_r,temp_m3_7_18_i,temp_m3_7_22_r,temp_m3_7_22_i,temp_b3_3_18_r,temp_b3_3_18_i,temp_b3_3_22_r,temp_b3_3_22_i,temp_b3_7_18_r,temp_b3_7_18_i,temp_b3_7_22_r,temp_b3_7_22_i);
MULT MULT555 (clk,temp_b2_3_19_r,temp_b2_3_19_i,temp_b2_3_23_r,temp_b2_3_23_i,temp_b2_7_19_r,temp_b2_7_19_i,temp_b2_7_23_r,temp_b2_7_23_i,temp_m3_3_19_r,temp_m3_3_19_i,temp_m3_3_23_r,temp_m3_3_23_i,temp_m3_7_19_r,temp_m3_7_19_i,temp_m3_7_23_r,temp_m3_7_23_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly555 (clk,temp_m3_3_19_r,temp_m3_3_19_i,temp_m3_3_23_r,temp_m3_3_23_i,temp_m3_7_19_r,temp_m3_7_19_i,temp_m3_7_23_r,temp_m3_7_23_i,temp_b3_3_19_r,temp_b3_3_19_i,temp_b3_3_23_r,temp_b3_3_23_i,temp_b3_7_19_r,temp_b3_7_19_i,temp_b3_7_23_r,temp_b3_7_23_i);
MULT MULT556 (clk,temp_b2_3_20_r,temp_b2_3_20_i,temp_b2_3_24_r,temp_b2_3_24_i,temp_b2_7_20_r,temp_b2_7_20_i,temp_b2_7_24_r,temp_b2_7_24_i,temp_m3_3_20_r,temp_m3_3_20_i,temp_m3_3_24_r,temp_m3_3_24_i,temp_m3_7_20_r,temp_m3_7_20_i,temp_m3_7_24_r,temp_m3_7_24_i,`W12_real,`W12_imag,`W8_real,`W8_imag,`W20_real,`W20_imag);
butterfly butterfly556 (clk,temp_m3_3_20_r,temp_m3_3_20_i,temp_m3_3_24_r,temp_m3_3_24_i,temp_m3_7_20_r,temp_m3_7_20_i,temp_m3_7_24_r,temp_m3_7_24_i,temp_b3_3_20_r,temp_b3_3_20_i,temp_b3_3_24_r,temp_b3_3_24_i,temp_b3_7_20_r,temp_b3_7_20_i,temp_b3_7_24_r,temp_b3_7_24_i);
MULT MULT557 (clk,temp_b2_4_17_r,temp_b2_4_17_i,temp_b2_4_21_r,temp_b2_4_21_i,temp_b2_8_17_r,temp_b2_8_17_i,temp_b2_8_21_r,temp_b2_8_21_i,temp_m3_4_17_r,temp_m3_4_17_i,temp_m3_4_21_r,temp_m3_4_21_i,temp_m3_8_17_r,temp_m3_8_17_i,temp_m3_8_21_r,temp_m3_8_21_i,`W0_real,`W0_imag,`W12_real,`W12_imag,`W12_real,`W12_imag);
butterfly butterfly557 (clk,temp_m3_4_17_r,temp_m3_4_17_i,temp_m3_4_21_r,temp_m3_4_21_i,temp_m3_8_17_r,temp_m3_8_17_i,temp_m3_8_21_r,temp_m3_8_21_i,temp_b3_4_17_r,temp_b3_4_17_i,temp_b3_4_21_r,temp_b3_4_21_i,temp_b3_8_17_r,temp_b3_8_17_i,temp_b3_8_21_r,temp_b3_8_21_i);
MULT MULT558 (clk,temp_b2_4_18_r,temp_b2_4_18_i,temp_b2_4_22_r,temp_b2_4_22_i,temp_b2_8_18_r,temp_b2_8_18_i,temp_b2_8_22_r,temp_b2_8_22_i,temp_m3_4_18_r,temp_m3_4_18_i,temp_m3_4_22_r,temp_m3_4_22_i,temp_m3_8_18_r,temp_m3_8_18_i,temp_m3_8_22_r,temp_m3_8_22_i,`W4_real,`W4_imag,`W12_real,`W12_imag,`W16_real,`W16_imag);
butterfly butterfly558 (clk,temp_m3_4_18_r,temp_m3_4_18_i,temp_m3_4_22_r,temp_m3_4_22_i,temp_m3_8_18_r,temp_m3_8_18_i,temp_m3_8_22_r,temp_m3_8_22_i,temp_b3_4_18_r,temp_b3_4_18_i,temp_b3_4_22_r,temp_b3_4_22_i,temp_b3_8_18_r,temp_b3_8_18_i,temp_b3_8_22_r,temp_b3_8_22_i);
MULT MULT559 (clk,temp_b2_4_19_r,temp_b2_4_19_i,temp_b2_4_23_r,temp_b2_4_23_i,temp_b2_8_19_r,temp_b2_8_19_i,temp_b2_8_23_r,temp_b2_8_23_i,temp_m3_4_19_r,temp_m3_4_19_i,temp_m3_4_23_r,temp_m3_4_23_i,temp_m3_8_19_r,temp_m3_8_19_i,temp_m3_8_23_r,temp_m3_8_23_i,`W8_real,`W8_imag,`W12_real,`W12_imag,`W20_real,`W20_imag);
butterfly butterfly559 (clk,temp_m3_4_19_r,temp_m3_4_19_i,temp_m3_4_23_r,temp_m3_4_23_i,temp_m3_8_19_r,temp_m3_8_19_i,temp_m3_8_23_r,temp_m3_8_23_i,temp_b3_4_19_r,temp_b3_4_19_i,temp_b3_4_23_r,temp_b3_4_23_i,temp_b3_8_19_r,temp_b3_8_19_i,temp_b3_8_23_r,temp_b3_8_23_i);
MULT MULT560 (clk,temp_b2_4_20_r,temp_b2_4_20_i,temp_b2_4_24_r,temp_b2_4_24_i,temp_b2_8_20_r,temp_b2_8_20_i,temp_b2_8_24_r,temp_b2_8_24_i,temp_m3_4_20_r,temp_m3_4_20_i,temp_m3_4_24_r,temp_m3_4_24_i,temp_m3_8_20_r,temp_m3_8_20_i,temp_m3_8_24_r,temp_m3_8_24_i,`W12_real,`W12_imag,`W12_real,`W12_imag,`W24_real,`W24_imag);
butterfly butterfly560 (clk,temp_m3_4_20_r,temp_m3_4_20_i,temp_m3_4_24_r,temp_m3_4_24_i,temp_m3_8_20_r,temp_m3_8_20_i,temp_m3_8_24_r,temp_m3_8_24_i,temp_b3_4_20_r,temp_b3_4_20_i,temp_b3_4_24_r,temp_b3_4_24_i,temp_b3_8_20_r,temp_b3_8_20_i,temp_b3_8_24_r,temp_b3_8_24_i);
MULT MULT561 (clk,temp_b2_1_25_r,temp_b2_1_25_i,temp_b2_1_29_r,temp_b2_1_29_i,temp_b2_5_25_r,temp_b2_5_25_i,temp_b2_5_29_r,temp_b2_5_29_i,temp_m3_1_25_r,temp_m3_1_25_i,temp_m3_1_29_r,temp_m3_1_29_i,temp_m3_5_25_r,temp_m3_5_25_i,temp_m3_5_29_r,temp_m3_5_29_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly561 (clk,temp_m3_1_25_r,temp_m3_1_25_i,temp_m3_1_29_r,temp_m3_1_29_i,temp_m3_5_25_r,temp_m3_5_25_i,temp_m3_5_29_r,temp_m3_5_29_i,temp_b3_1_25_r,temp_b3_1_25_i,temp_b3_1_29_r,temp_b3_1_29_i,temp_b3_5_25_r,temp_b3_5_25_i,temp_b3_5_29_r,temp_b3_5_29_i);
MULT MULT562 (clk,temp_b2_1_26_r,temp_b2_1_26_i,temp_b2_1_30_r,temp_b2_1_30_i,temp_b2_5_26_r,temp_b2_5_26_i,temp_b2_5_30_r,temp_b2_5_30_i,temp_m3_1_26_r,temp_m3_1_26_i,temp_m3_1_30_r,temp_m3_1_30_i,temp_m3_5_26_r,temp_m3_5_26_i,temp_m3_5_30_r,temp_m3_5_30_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly562 (clk,temp_m3_1_26_r,temp_m3_1_26_i,temp_m3_1_30_r,temp_m3_1_30_i,temp_m3_5_26_r,temp_m3_5_26_i,temp_m3_5_30_r,temp_m3_5_30_i,temp_b3_1_26_r,temp_b3_1_26_i,temp_b3_1_30_r,temp_b3_1_30_i,temp_b3_5_26_r,temp_b3_5_26_i,temp_b3_5_30_r,temp_b3_5_30_i);
MULT MULT563 (clk,temp_b2_1_27_r,temp_b2_1_27_i,temp_b2_1_31_r,temp_b2_1_31_i,temp_b2_5_27_r,temp_b2_5_27_i,temp_b2_5_31_r,temp_b2_5_31_i,temp_m3_1_27_r,temp_m3_1_27_i,temp_m3_1_31_r,temp_m3_1_31_i,temp_m3_5_27_r,temp_m3_5_27_i,temp_m3_5_31_r,temp_m3_5_31_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly563 (clk,temp_m3_1_27_r,temp_m3_1_27_i,temp_m3_1_31_r,temp_m3_1_31_i,temp_m3_5_27_r,temp_m3_5_27_i,temp_m3_5_31_r,temp_m3_5_31_i,temp_b3_1_27_r,temp_b3_1_27_i,temp_b3_1_31_r,temp_b3_1_31_i,temp_b3_5_27_r,temp_b3_5_27_i,temp_b3_5_31_r,temp_b3_5_31_i);
MULT MULT564 (clk,temp_b2_1_28_r,temp_b2_1_28_i,temp_b2_1_32_r,temp_b2_1_32_i,temp_b2_5_28_r,temp_b2_5_28_i,temp_b2_5_32_r,temp_b2_5_32_i,temp_m3_1_28_r,temp_m3_1_28_i,temp_m3_1_32_r,temp_m3_1_32_i,temp_m3_5_28_r,temp_m3_5_28_i,temp_m3_5_32_r,temp_m3_5_32_i,`W12_real,`W12_imag,`W0_real,`W0_imag,`W12_real,`W12_imag);
butterfly butterfly564 (clk,temp_m3_1_28_r,temp_m3_1_28_i,temp_m3_1_32_r,temp_m3_1_32_i,temp_m3_5_28_r,temp_m3_5_28_i,temp_m3_5_32_r,temp_m3_5_32_i,temp_b3_1_28_r,temp_b3_1_28_i,temp_b3_1_32_r,temp_b3_1_32_i,temp_b3_5_28_r,temp_b3_5_28_i,temp_b3_5_32_r,temp_b3_5_32_i);
MULT MULT565 (clk,temp_b2_2_25_r,temp_b2_2_25_i,temp_b2_2_29_r,temp_b2_2_29_i,temp_b2_6_25_r,temp_b2_6_25_i,temp_b2_6_29_r,temp_b2_6_29_i,temp_m3_2_25_r,temp_m3_2_25_i,temp_m3_2_29_r,temp_m3_2_29_i,temp_m3_6_25_r,temp_m3_6_25_i,temp_m3_6_29_r,temp_m3_6_29_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly565 (clk,temp_m3_2_25_r,temp_m3_2_25_i,temp_m3_2_29_r,temp_m3_2_29_i,temp_m3_6_25_r,temp_m3_6_25_i,temp_m3_6_29_r,temp_m3_6_29_i,temp_b3_2_25_r,temp_b3_2_25_i,temp_b3_2_29_r,temp_b3_2_29_i,temp_b3_6_25_r,temp_b3_6_25_i,temp_b3_6_29_r,temp_b3_6_29_i);
MULT MULT566 (clk,temp_b2_2_26_r,temp_b2_2_26_i,temp_b2_2_30_r,temp_b2_2_30_i,temp_b2_6_26_r,temp_b2_6_26_i,temp_b2_6_30_r,temp_b2_6_30_i,temp_m3_2_26_r,temp_m3_2_26_i,temp_m3_2_30_r,temp_m3_2_30_i,temp_m3_6_26_r,temp_m3_6_26_i,temp_m3_6_30_r,temp_m3_6_30_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly566 (clk,temp_m3_2_26_r,temp_m3_2_26_i,temp_m3_2_30_r,temp_m3_2_30_i,temp_m3_6_26_r,temp_m3_6_26_i,temp_m3_6_30_r,temp_m3_6_30_i,temp_b3_2_26_r,temp_b3_2_26_i,temp_b3_2_30_r,temp_b3_2_30_i,temp_b3_6_26_r,temp_b3_6_26_i,temp_b3_6_30_r,temp_b3_6_30_i);
MULT MULT567 (clk,temp_b2_2_27_r,temp_b2_2_27_i,temp_b2_2_31_r,temp_b2_2_31_i,temp_b2_6_27_r,temp_b2_6_27_i,temp_b2_6_31_r,temp_b2_6_31_i,temp_m3_2_27_r,temp_m3_2_27_i,temp_m3_2_31_r,temp_m3_2_31_i,temp_m3_6_27_r,temp_m3_6_27_i,temp_m3_6_31_r,temp_m3_6_31_i,`W8_real,`W8_imag,`W4_real,`W4_imag,`W12_real,`W12_imag);
butterfly butterfly567 (clk,temp_m3_2_27_r,temp_m3_2_27_i,temp_m3_2_31_r,temp_m3_2_31_i,temp_m3_6_27_r,temp_m3_6_27_i,temp_m3_6_31_r,temp_m3_6_31_i,temp_b3_2_27_r,temp_b3_2_27_i,temp_b3_2_31_r,temp_b3_2_31_i,temp_b3_6_27_r,temp_b3_6_27_i,temp_b3_6_31_r,temp_b3_6_31_i);
MULT MULT568 (clk,temp_b2_2_28_r,temp_b2_2_28_i,temp_b2_2_32_r,temp_b2_2_32_i,temp_b2_6_28_r,temp_b2_6_28_i,temp_b2_6_32_r,temp_b2_6_32_i,temp_m3_2_28_r,temp_m3_2_28_i,temp_m3_2_32_r,temp_m3_2_32_i,temp_m3_6_28_r,temp_m3_6_28_i,temp_m3_6_32_r,temp_m3_6_32_i,`W12_real,`W12_imag,`W4_real,`W4_imag,`W16_real,`W16_imag);
butterfly butterfly568 (clk,temp_m3_2_28_r,temp_m3_2_28_i,temp_m3_2_32_r,temp_m3_2_32_i,temp_m3_6_28_r,temp_m3_6_28_i,temp_m3_6_32_r,temp_m3_6_32_i,temp_b3_2_28_r,temp_b3_2_28_i,temp_b3_2_32_r,temp_b3_2_32_i,temp_b3_6_28_r,temp_b3_6_28_i,temp_b3_6_32_r,temp_b3_6_32_i);
MULT MULT569 (clk,temp_b2_3_25_r,temp_b2_3_25_i,temp_b2_3_29_r,temp_b2_3_29_i,temp_b2_7_25_r,temp_b2_7_25_i,temp_b2_7_29_r,temp_b2_7_29_i,temp_m3_3_25_r,temp_m3_3_25_i,temp_m3_3_29_r,temp_m3_3_29_i,temp_m3_7_25_r,temp_m3_7_25_i,temp_m3_7_29_r,temp_m3_7_29_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly569 (clk,temp_m3_3_25_r,temp_m3_3_25_i,temp_m3_3_29_r,temp_m3_3_29_i,temp_m3_7_25_r,temp_m3_7_25_i,temp_m3_7_29_r,temp_m3_7_29_i,temp_b3_3_25_r,temp_b3_3_25_i,temp_b3_3_29_r,temp_b3_3_29_i,temp_b3_7_25_r,temp_b3_7_25_i,temp_b3_7_29_r,temp_b3_7_29_i);
MULT MULT570 (clk,temp_b2_3_26_r,temp_b2_3_26_i,temp_b2_3_30_r,temp_b2_3_30_i,temp_b2_7_26_r,temp_b2_7_26_i,temp_b2_7_30_r,temp_b2_7_30_i,temp_m3_3_26_r,temp_m3_3_26_i,temp_m3_3_30_r,temp_m3_3_30_i,temp_m3_7_26_r,temp_m3_7_26_i,temp_m3_7_30_r,temp_m3_7_30_i,`W4_real,`W4_imag,`W8_real,`W8_imag,`W12_real,`W12_imag);
butterfly butterfly570 (clk,temp_m3_3_26_r,temp_m3_3_26_i,temp_m3_3_30_r,temp_m3_3_30_i,temp_m3_7_26_r,temp_m3_7_26_i,temp_m3_7_30_r,temp_m3_7_30_i,temp_b3_3_26_r,temp_b3_3_26_i,temp_b3_3_30_r,temp_b3_3_30_i,temp_b3_7_26_r,temp_b3_7_26_i,temp_b3_7_30_r,temp_b3_7_30_i);
MULT MULT571 (clk,temp_b2_3_27_r,temp_b2_3_27_i,temp_b2_3_31_r,temp_b2_3_31_i,temp_b2_7_27_r,temp_b2_7_27_i,temp_b2_7_31_r,temp_b2_7_31_i,temp_m3_3_27_r,temp_m3_3_27_i,temp_m3_3_31_r,temp_m3_3_31_i,temp_m3_7_27_r,temp_m3_7_27_i,temp_m3_7_31_r,temp_m3_7_31_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly571 (clk,temp_m3_3_27_r,temp_m3_3_27_i,temp_m3_3_31_r,temp_m3_3_31_i,temp_m3_7_27_r,temp_m3_7_27_i,temp_m3_7_31_r,temp_m3_7_31_i,temp_b3_3_27_r,temp_b3_3_27_i,temp_b3_3_31_r,temp_b3_3_31_i,temp_b3_7_27_r,temp_b3_7_27_i,temp_b3_7_31_r,temp_b3_7_31_i);
MULT MULT572 (clk,temp_b2_3_28_r,temp_b2_3_28_i,temp_b2_3_32_r,temp_b2_3_32_i,temp_b2_7_28_r,temp_b2_7_28_i,temp_b2_7_32_r,temp_b2_7_32_i,temp_m3_3_28_r,temp_m3_3_28_i,temp_m3_3_32_r,temp_m3_3_32_i,temp_m3_7_28_r,temp_m3_7_28_i,temp_m3_7_32_r,temp_m3_7_32_i,`W12_real,`W12_imag,`W8_real,`W8_imag,`W20_real,`W20_imag);
butterfly butterfly572 (clk,temp_m3_3_28_r,temp_m3_3_28_i,temp_m3_3_32_r,temp_m3_3_32_i,temp_m3_7_28_r,temp_m3_7_28_i,temp_m3_7_32_r,temp_m3_7_32_i,temp_b3_3_28_r,temp_b3_3_28_i,temp_b3_3_32_r,temp_b3_3_32_i,temp_b3_7_28_r,temp_b3_7_28_i,temp_b3_7_32_r,temp_b3_7_32_i);
MULT MULT573 (clk,temp_b2_4_25_r,temp_b2_4_25_i,temp_b2_4_29_r,temp_b2_4_29_i,temp_b2_8_25_r,temp_b2_8_25_i,temp_b2_8_29_r,temp_b2_8_29_i,temp_m3_4_25_r,temp_m3_4_25_i,temp_m3_4_29_r,temp_m3_4_29_i,temp_m3_8_25_r,temp_m3_8_25_i,temp_m3_8_29_r,temp_m3_8_29_i,`W0_real,`W0_imag,`W12_real,`W12_imag,`W12_real,`W12_imag);
butterfly butterfly573 (clk,temp_m3_4_25_r,temp_m3_4_25_i,temp_m3_4_29_r,temp_m3_4_29_i,temp_m3_8_25_r,temp_m3_8_25_i,temp_m3_8_29_r,temp_m3_8_29_i,temp_b3_4_25_r,temp_b3_4_25_i,temp_b3_4_29_r,temp_b3_4_29_i,temp_b3_8_25_r,temp_b3_8_25_i,temp_b3_8_29_r,temp_b3_8_29_i);
MULT MULT574 (clk,temp_b2_4_26_r,temp_b2_4_26_i,temp_b2_4_30_r,temp_b2_4_30_i,temp_b2_8_26_r,temp_b2_8_26_i,temp_b2_8_30_r,temp_b2_8_30_i,temp_m3_4_26_r,temp_m3_4_26_i,temp_m3_4_30_r,temp_m3_4_30_i,temp_m3_8_26_r,temp_m3_8_26_i,temp_m3_8_30_r,temp_m3_8_30_i,`W4_real,`W4_imag,`W12_real,`W12_imag,`W16_real,`W16_imag);
butterfly butterfly574 (clk,temp_m3_4_26_r,temp_m3_4_26_i,temp_m3_4_30_r,temp_m3_4_30_i,temp_m3_8_26_r,temp_m3_8_26_i,temp_m3_8_30_r,temp_m3_8_30_i,temp_b3_4_26_r,temp_b3_4_26_i,temp_b3_4_30_r,temp_b3_4_30_i,temp_b3_8_26_r,temp_b3_8_26_i,temp_b3_8_30_r,temp_b3_8_30_i);
MULT MULT575 (clk,temp_b2_4_27_r,temp_b2_4_27_i,temp_b2_4_31_r,temp_b2_4_31_i,temp_b2_8_27_r,temp_b2_8_27_i,temp_b2_8_31_r,temp_b2_8_31_i,temp_m3_4_27_r,temp_m3_4_27_i,temp_m3_4_31_r,temp_m3_4_31_i,temp_m3_8_27_r,temp_m3_8_27_i,temp_m3_8_31_r,temp_m3_8_31_i,`W8_real,`W8_imag,`W12_real,`W12_imag,`W20_real,`W20_imag);
butterfly butterfly575 (clk,temp_m3_4_27_r,temp_m3_4_27_i,temp_m3_4_31_r,temp_m3_4_31_i,temp_m3_8_27_r,temp_m3_8_27_i,temp_m3_8_31_r,temp_m3_8_31_i,temp_b3_4_27_r,temp_b3_4_27_i,temp_b3_4_31_r,temp_b3_4_31_i,temp_b3_8_27_r,temp_b3_8_27_i,temp_b3_8_31_r,temp_b3_8_31_i);
MULT MULT576 (clk,temp_b2_4_28_r,temp_b2_4_28_i,temp_b2_4_32_r,temp_b2_4_32_i,temp_b2_8_28_r,temp_b2_8_28_i,temp_b2_8_32_r,temp_b2_8_32_i,temp_m3_4_28_r,temp_m3_4_28_i,temp_m3_4_32_r,temp_m3_4_32_i,temp_m3_8_28_r,temp_m3_8_28_i,temp_m3_8_32_r,temp_m3_8_32_i,`W12_real,`W12_imag,`W12_real,`W12_imag,`W24_real,`W24_imag);
butterfly butterfly576 (clk,temp_m3_4_28_r,temp_m3_4_28_i,temp_m3_4_32_r,temp_m3_4_32_i,temp_m3_8_28_r,temp_m3_8_28_i,temp_m3_8_32_r,temp_m3_8_32_i,temp_b3_4_28_r,temp_b3_4_28_i,temp_b3_4_32_r,temp_b3_4_32_i,temp_b3_8_28_r,temp_b3_8_28_i,temp_b3_8_32_r,temp_b3_8_32_i);
MULT MULT577 (clk,temp_b2_9_1_r,temp_b2_9_1_i,temp_b2_9_5_r,temp_b2_9_5_i,temp_b2_13_1_r,temp_b2_13_1_i,temp_b2_13_5_r,temp_b2_13_5_i,temp_m3_9_1_r,temp_m3_9_1_i,temp_m3_9_5_r,temp_m3_9_5_i,temp_m3_13_1_r,temp_m3_13_1_i,temp_m3_13_5_r,temp_m3_13_5_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly577 (clk,temp_m3_9_1_r,temp_m3_9_1_i,temp_m3_9_5_r,temp_m3_9_5_i,temp_m3_13_1_r,temp_m3_13_1_i,temp_m3_13_5_r,temp_m3_13_5_i,temp_b3_9_1_r,temp_b3_9_1_i,temp_b3_9_5_r,temp_b3_9_5_i,temp_b3_13_1_r,temp_b3_13_1_i,temp_b3_13_5_r,temp_b3_13_5_i);
MULT MULT578 (clk,temp_b2_9_2_r,temp_b2_9_2_i,temp_b2_9_6_r,temp_b2_9_6_i,temp_b2_13_2_r,temp_b2_13_2_i,temp_b2_13_6_r,temp_b2_13_6_i,temp_m3_9_2_r,temp_m3_9_2_i,temp_m3_9_6_r,temp_m3_9_6_i,temp_m3_13_2_r,temp_m3_13_2_i,temp_m3_13_6_r,temp_m3_13_6_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly578 (clk,temp_m3_9_2_r,temp_m3_9_2_i,temp_m3_9_6_r,temp_m3_9_6_i,temp_m3_13_2_r,temp_m3_13_2_i,temp_m3_13_6_r,temp_m3_13_6_i,temp_b3_9_2_r,temp_b3_9_2_i,temp_b3_9_6_r,temp_b3_9_6_i,temp_b3_13_2_r,temp_b3_13_2_i,temp_b3_13_6_r,temp_b3_13_6_i);
MULT MULT579 (clk,temp_b2_9_3_r,temp_b2_9_3_i,temp_b2_9_7_r,temp_b2_9_7_i,temp_b2_13_3_r,temp_b2_13_3_i,temp_b2_13_7_r,temp_b2_13_7_i,temp_m3_9_3_r,temp_m3_9_3_i,temp_m3_9_7_r,temp_m3_9_7_i,temp_m3_13_3_r,temp_m3_13_3_i,temp_m3_13_7_r,temp_m3_13_7_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly579 (clk,temp_m3_9_3_r,temp_m3_9_3_i,temp_m3_9_7_r,temp_m3_9_7_i,temp_m3_13_3_r,temp_m3_13_3_i,temp_m3_13_7_r,temp_m3_13_7_i,temp_b3_9_3_r,temp_b3_9_3_i,temp_b3_9_7_r,temp_b3_9_7_i,temp_b3_13_3_r,temp_b3_13_3_i,temp_b3_13_7_r,temp_b3_13_7_i);
MULT MULT580 (clk,temp_b2_9_4_r,temp_b2_9_4_i,temp_b2_9_8_r,temp_b2_9_8_i,temp_b2_13_4_r,temp_b2_13_4_i,temp_b2_13_8_r,temp_b2_13_8_i,temp_m3_9_4_r,temp_m3_9_4_i,temp_m3_9_8_r,temp_m3_9_8_i,temp_m3_13_4_r,temp_m3_13_4_i,temp_m3_13_8_r,temp_m3_13_8_i,`W12_real,`W12_imag,`W0_real,`W0_imag,`W12_real,`W12_imag);
butterfly butterfly580 (clk,temp_m3_9_4_r,temp_m3_9_4_i,temp_m3_9_8_r,temp_m3_9_8_i,temp_m3_13_4_r,temp_m3_13_4_i,temp_m3_13_8_r,temp_m3_13_8_i,temp_b3_9_4_r,temp_b3_9_4_i,temp_b3_9_8_r,temp_b3_9_8_i,temp_b3_13_4_r,temp_b3_13_4_i,temp_b3_13_8_r,temp_b3_13_8_i);
MULT MULT581 (clk,temp_b2_10_1_r,temp_b2_10_1_i,temp_b2_10_5_r,temp_b2_10_5_i,temp_b2_14_1_r,temp_b2_14_1_i,temp_b2_14_5_r,temp_b2_14_5_i,temp_m3_10_1_r,temp_m3_10_1_i,temp_m3_10_5_r,temp_m3_10_5_i,temp_m3_14_1_r,temp_m3_14_1_i,temp_m3_14_5_r,temp_m3_14_5_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly581 (clk,temp_m3_10_1_r,temp_m3_10_1_i,temp_m3_10_5_r,temp_m3_10_5_i,temp_m3_14_1_r,temp_m3_14_1_i,temp_m3_14_5_r,temp_m3_14_5_i,temp_b3_10_1_r,temp_b3_10_1_i,temp_b3_10_5_r,temp_b3_10_5_i,temp_b3_14_1_r,temp_b3_14_1_i,temp_b3_14_5_r,temp_b3_14_5_i);
MULT MULT582 (clk,temp_b2_10_2_r,temp_b2_10_2_i,temp_b2_10_6_r,temp_b2_10_6_i,temp_b2_14_2_r,temp_b2_14_2_i,temp_b2_14_6_r,temp_b2_14_6_i,temp_m3_10_2_r,temp_m3_10_2_i,temp_m3_10_6_r,temp_m3_10_6_i,temp_m3_14_2_r,temp_m3_14_2_i,temp_m3_14_6_r,temp_m3_14_6_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly582 (clk,temp_m3_10_2_r,temp_m3_10_2_i,temp_m3_10_6_r,temp_m3_10_6_i,temp_m3_14_2_r,temp_m3_14_2_i,temp_m3_14_6_r,temp_m3_14_6_i,temp_b3_10_2_r,temp_b3_10_2_i,temp_b3_10_6_r,temp_b3_10_6_i,temp_b3_14_2_r,temp_b3_14_2_i,temp_b3_14_6_r,temp_b3_14_6_i);
MULT MULT583 (clk,temp_b2_10_3_r,temp_b2_10_3_i,temp_b2_10_7_r,temp_b2_10_7_i,temp_b2_14_3_r,temp_b2_14_3_i,temp_b2_14_7_r,temp_b2_14_7_i,temp_m3_10_3_r,temp_m3_10_3_i,temp_m3_10_7_r,temp_m3_10_7_i,temp_m3_14_3_r,temp_m3_14_3_i,temp_m3_14_7_r,temp_m3_14_7_i,`W8_real,`W8_imag,`W4_real,`W4_imag,`W12_real,`W12_imag);
butterfly butterfly583 (clk,temp_m3_10_3_r,temp_m3_10_3_i,temp_m3_10_7_r,temp_m3_10_7_i,temp_m3_14_3_r,temp_m3_14_3_i,temp_m3_14_7_r,temp_m3_14_7_i,temp_b3_10_3_r,temp_b3_10_3_i,temp_b3_10_7_r,temp_b3_10_7_i,temp_b3_14_3_r,temp_b3_14_3_i,temp_b3_14_7_r,temp_b3_14_7_i);
MULT MULT584 (clk,temp_b2_10_4_r,temp_b2_10_4_i,temp_b2_10_8_r,temp_b2_10_8_i,temp_b2_14_4_r,temp_b2_14_4_i,temp_b2_14_8_r,temp_b2_14_8_i,temp_m3_10_4_r,temp_m3_10_4_i,temp_m3_10_8_r,temp_m3_10_8_i,temp_m3_14_4_r,temp_m3_14_4_i,temp_m3_14_8_r,temp_m3_14_8_i,`W12_real,`W12_imag,`W4_real,`W4_imag,`W16_real,`W16_imag);
butterfly butterfly584 (clk,temp_m3_10_4_r,temp_m3_10_4_i,temp_m3_10_8_r,temp_m3_10_8_i,temp_m3_14_4_r,temp_m3_14_4_i,temp_m3_14_8_r,temp_m3_14_8_i,temp_b3_10_4_r,temp_b3_10_4_i,temp_b3_10_8_r,temp_b3_10_8_i,temp_b3_14_4_r,temp_b3_14_4_i,temp_b3_14_8_r,temp_b3_14_8_i);
MULT MULT585 (clk,temp_b2_11_1_r,temp_b2_11_1_i,temp_b2_11_5_r,temp_b2_11_5_i,temp_b2_15_1_r,temp_b2_15_1_i,temp_b2_15_5_r,temp_b2_15_5_i,temp_m3_11_1_r,temp_m3_11_1_i,temp_m3_11_5_r,temp_m3_11_5_i,temp_m3_15_1_r,temp_m3_15_1_i,temp_m3_15_5_r,temp_m3_15_5_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly585 (clk,temp_m3_11_1_r,temp_m3_11_1_i,temp_m3_11_5_r,temp_m3_11_5_i,temp_m3_15_1_r,temp_m3_15_1_i,temp_m3_15_5_r,temp_m3_15_5_i,temp_b3_11_1_r,temp_b3_11_1_i,temp_b3_11_5_r,temp_b3_11_5_i,temp_b3_15_1_r,temp_b3_15_1_i,temp_b3_15_5_r,temp_b3_15_5_i);
MULT MULT586 (clk,temp_b2_11_2_r,temp_b2_11_2_i,temp_b2_11_6_r,temp_b2_11_6_i,temp_b2_15_2_r,temp_b2_15_2_i,temp_b2_15_6_r,temp_b2_15_6_i,temp_m3_11_2_r,temp_m3_11_2_i,temp_m3_11_6_r,temp_m3_11_6_i,temp_m3_15_2_r,temp_m3_15_2_i,temp_m3_15_6_r,temp_m3_15_6_i,`W4_real,`W4_imag,`W8_real,`W8_imag,`W12_real,`W12_imag);
butterfly butterfly586 (clk,temp_m3_11_2_r,temp_m3_11_2_i,temp_m3_11_6_r,temp_m3_11_6_i,temp_m3_15_2_r,temp_m3_15_2_i,temp_m3_15_6_r,temp_m3_15_6_i,temp_b3_11_2_r,temp_b3_11_2_i,temp_b3_11_6_r,temp_b3_11_6_i,temp_b3_15_2_r,temp_b3_15_2_i,temp_b3_15_6_r,temp_b3_15_6_i);
MULT MULT587 (clk,temp_b2_11_3_r,temp_b2_11_3_i,temp_b2_11_7_r,temp_b2_11_7_i,temp_b2_15_3_r,temp_b2_15_3_i,temp_b2_15_7_r,temp_b2_15_7_i,temp_m3_11_3_r,temp_m3_11_3_i,temp_m3_11_7_r,temp_m3_11_7_i,temp_m3_15_3_r,temp_m3_15_3_i,temp_m3_15_7_r,temp_m3_15_7_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly587 (clk,temp_m3_11_3_r,temp_m3_11_3_i,temp_m3_11_7_r,temp_m3_11_7_i,temp_m3_15_3_r,temp_m3_15_3_i,temp_m3_15_7_r,temp_m3_15_7_i,temp_b3_11_3_r,temp_b3_11_3_i,temp_b3_11_7_r,temp_b3_11_7_i,temp_b3_15_3_r,temp_b3_15_3_i,temp_b3_15_7_r,temp_b3_15_7_i);
MULT MULT588 (clk,temp_b2_11_4_r,temp_b2_11_4_i,temp_b2_11_8_r,temp_b2_11_8_i,temp_b2_15_4_r,temp_b2_15_4_i,temp_b2_15_8_r,temp_b2_15_8_i,temp_m3_11_4_r,temp_m3_11_4_i,temp_m3_11_8_r,temp_m3_11_8_i,temp_m3_15_4_r,temp_m3_15_4_i,temp_m3_15_8_r,temp_m3_15_8_i,`W12_real,`W12_imag,`W8_real,`W8_imag,`W20_real,`W20_imag);
butterfly butterfly588 (clk,temp_m3_11_4_r,temp_m3_11_4_i,temp_m3_11_8_r,temp_m3_11_8_i,temp_m3_15_4_r,temp_m3_15_4_i,temp_m3_15_8_r,temp_m3_15_8_i,temp_b3_11_4_r,temp_b3_11_4_i,temp_b3_11_8_r,temp_b3_11_8_i,temp_b3_15_4_r,temp_b3_15_4_i,temp_b3_15_8_r,temp_b3_15_8_i);
MULT MULT589 (clk,temp_b2_12_1_r,temp_b2_12_1_i,temp_b2_12_5_r,temp_b2_12_5_i,temp_b2_16_1_r,temp_b2_16_1_i,temp_b2_16_5_r,temp_b2_16_5_i,temp_m3_12_1_r,temp_m3_12_1_i,temp_m3_12_5_r,temp_m3_12_5_i,temp_m3_16_1_r,temp_m3_16_1_i,temp_m3_16_5_r,temp_m3_16_5_i,`W0_real,`W0_imag,`W12_real,`W12_imag,`W12_real,`W12_imag);
butterfly butterfly589 (clk,temp_m3_12_1_r,temp_m3_12_1_i,temp_m3_12_5_r,temp_m3_12_5_i,temp_m3_16_1_r,temp_m3_16_1_i,temp_m3_16_5_r,temp_m3_16_5_i,temp_b3_12_1_r,temp_b3_12_1_i,temp_b3_12_5_r,temp_b3_12_5_i,temp_b3_16_1_r,temp_b3_16_1_i,temp_b3_16_5_r,temp_b3_16_5_i);
MULT MULT590 (clk,temp_b2_12_2_r,temp_b2_12_2_i,temp_b2_12_6_r,temp_b2_12_6_i,temp_b2_16_2_r,temp_b2_16_2_i,temp_b2_16_6_r,temp_b2_16_6_i,temp_m3_12_2_r,temp_m3_12_2_i,temp_m3_12_6_r,temp_m3_12_6_i,temp_m3_16_2_r,temp_m3_16_2_i,temp_m3_16_6_r,temp_m3_16_6_i,`W4_real,`W4_imag,`W12_real,`W12_imag,`W16_real,`W16_imag);
butterfly butterfly590 (clk,temp_m3_12_2_r,temp_m3_12_2_i,temp_m3_12_6_r,temp_m3_12_6_i,temp_m3_16_2_r,temp_m3_16_2_i,temp_m3_16_6_r,temp_m3_16_6_i,temp_b3_12_2_r,temp_b3_12_2_i,temp_b3_12_6_r,temp_b3_12_6_i,temp_b3_16_2_r,temp_b3_16_2_i,temp_b3_16_6_r,temp_b3_16_6_i);
MULT MULT591 (clk,temp_b2_12_3_r,temp_b2_12_3_i,temp_b2_12_7_r,temp_b2_12_7_i,temp_b2_16_3_r,temp_b2_16_3_i,temp_b2_16_7_r,temp_b2_16_7_i,temp_m3_12_3_r,temp_m3_12_3_i,temp_m3_12_7_r,temp_m3_12_7_i,temp_m3_16_3_r,temp_m3_16_3_i,temp_m3_16_7_r,temp_m3_16_7_i,`W8_real,`W8_imag,`W12_real,`W12_imag,`W20_real,`W20_imag);
butterfly butterfly591 (clk,temp_m3_12_3_r,temp_m3_12_3_i,temp_m3_12_7_r,temp_m3_12_7_i,temp_m3_16_3_r,temp_m3_16_3_i,temp_m3_16_7_r,temp_m3_16_7_i,temp_b3_12_3_r,temp_b3_12_3_i,temp_b3_12_7_r,temp_b3_12_7_i,temp_b3_16_3_r,temp_b3_16_3_i,temp_b3_16_7_r,temp_b3_16_7_i);
MULT MULT592 (clk,temp_b2_12_4_r,temp_b2_12_4_i,temp_b2_12_8_r,temp_b2_12_8_i,temp_b2_16_4_r,temp_b2_16_4_i,temp_b2_16_8_r,temp_b2_16_8_i,temp_m3_12_4_r,temp_m3_12_4_i,temp_m3_12_8_r,temp_m3_12_8_i,temp_m3_16_4_r,temp_m3_16_4_i,temp_m3_16_8_r,temp_m3_16_8_i,`W12_real,`W12_imag,`W12_real,`W12_imag,`W24_real,`W24_imag);
butterfly butterfly592 (clk,temp_m3_12_4_r,temp_m3_12_4_i,temp_m3_12_8_r,temp_m3_12_8_i,temp_m3_16_4_r,temp_m3_16_4_i,temp_m3_16_8_r,temp_m3_16_8_i,temp_b3_12_4_r,temp_b3_12_4_i,temp_b3_12_8_r,temp_b3_12_8_i,temp_b3_16_4_r,temp_b3_16_4_i,temp_b3_16_8_r,temp_b3_16_8_i);
MULT MULT593 (clk,temp_b2_9_9_r,temp_b2_9_9_i,temp_b2_9_13_r,temp_b2_9_13_i,temp_b2_13_9_r,temp_b2_13_9_i,temp_b2_13_13_r,temp_b2_13_13_i,temp_m3_9_9_r,temp_m3_9_9_i,temp_m3_9_13_r,temp_m3_9_13_i,temp_m3_13_9_r,temp_m3_13_9_i,temp_m3_13_13_r,temp_m3_13_13_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly593 (clk,temp_m3_9_9_r,temp_m3_9_9_i,temp_m3_9_13_r,temp_m3_9_13_i,temp_m3_13_9_r,temp_m3_13_9_i,temp_m3_13_13_r,temp_m3_13_13_i,temp_b3_9_9_r,temp_b3_9_9_i,temp_b3_9_13_r,temp_b3_9_13_i,temp_b3_13_9_r,temp_b3_13_9_i,temp_b3_13_13_r,temp_b3_13_13_i);
MULT MULT594 (clk,temp_b2_9_10_r,temp_b2_9_10_i,temp_b2_9_14_r,temp_b2_9_14_i,temp_b2_13_10_r,temp_b2_13_10_i,temp_b2_13_14_r,temp_b2_13_14_i,temp_m3_9_10_r,temp_m3_9_10_i,temp_m3_9_14_r,temp_m3_9_14_i,temp_m3_13_10_r,temp_m3_13_10_i,temp_m3_13_14_r,temp_m3_13_14_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly594 (clk,temp_m3_9_10_r,temp_m3_9_10_i,temp_m3_9_14_r,temp_m3_9_14_i,temp_m3_13_10_r,temp_m3_13_10_i,temp_m3_13_14_r,temp_m3_13_14_i,temp_b3_9_10_r,temp_b3_9_10_i,temp_b3_9_14_r,temp_b3_9_14_i,temp_b3_13_10_r,temp_b3_13_10_i,temp_b3_13_14_r,temp_b3_13_14_i);
MULT MULT595 (clk,temp_b2_9_11_r,temp_b2_9_11_i,temp_b2_9_15_r,temp_b2_9_15_i,temp_b2_13_11_r,temp_b2_13_11_i,temp_b2_13_15_r,temp_b2_13_15_i,temp_m3_9_11_r,temp_m3_9_11_i,temp_m3_9_15_r,temp_m3_9_15_i,temp_m3_13_11_r,temp_m3_13_11_i,temp_m3_13_15_r,temp_m3_13_15_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly595 (clk,temp_m3_9_11_r,temp_m3_9_11_i,temp_m3_9_15_r,temp_m3_9_15_i,temp_m3_13_11_r,temp_m3_13_11_i,temp_m3_13_15_r,temp_m3_13_15_i,temp_b3_9_11_r,temp_b3_9_11_i,temp_b3_9_15_r,temp_b3_9_15_i,temp_b3_13_11_r,temp_b3_13_11_i,temp_b3_13_15_r,temp_b3_13_15_i);
MULT MULT596 (clk,temp_b2_9_12_r,temp_b2_9_12_i,temp_b2_9_16_r,temp_b2_9_16_i,temp_b2_13_12_r,temp_b2_13_12_i,temp_b2_13_16_r,temp_b2_13_16_i,temp_m3_9_12_r,temp_m3_9_12_i,temp_m3_9_16_r,temp_m3_9_16_i,temp_m3_13_12_r,temp_m3_13_12_i,temp_m3_13_16_r,temp_m3_13_16_i,`W12_real,`W12_imag,`W0_real,`W0_imag,`W12_real,`W12_imag);
butterfly butterfly596 (clk,temp_m3_9_12_r,temp_m3_9_12_i,temp_m3_9_16_r,temp_m3_9_16_i,temp_m3_13_12_r,temp_m3_13_12_i,temp_m3_13_16_r,temp_m3_13_16_i,temp_b3_9_12_r,temp_b3_9_12_i,temp_b3_9_16_r,temp_b3_9_16_i,temp_b3_13_12_r,temp_b3_13_12_i,temp_b3_13_16_r,temp_b3_13_16_i);
MULT MULT597 (clk,temp_b2_10_9_r,temp_b2_10_9_i,temp_b2_10_13_r,temp_b2_10_13_i,temp_b2_14_9_r,temp_b2_14_9_i,temp_b2_14_13_r,temp_b2_14_13_i,temp_m3_10_9_r,temp_m3_10_9_i,temp_m3_10_13_r,temp_m3_10_13_i,temp_m3_14_9_r,temp_m3_14_9_i,temp_m3_14_13_r,temp_m3_14_13_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly597 (clk,temp_m3_10_9_r,temp_m3_10_9_i,temp_m3_10_13_r,temp_m3_10_13_i,temp_m3_14_9_r,temp_m3_14_9_i,temp_m3_14_13_r,temp_m3_14_13_i,temp_b3_10_9_r,temp_b3_10_9_i,temp_b3_10_13_r,temp_b3_10_13_i,temp_b3_14_9_r,temp_b3_14_9_i,temp_b3_14_13_r,temp_b3_14_13_i);
MULT MULT598 (clk,temp_b2_10_10_r,temp_b2_10_10_i,temp_b2_10_14_r,temp_b2_10_14_i,temp_b2_14_10_r,temp_b2_14_10_i,temp_b2_14_14_r,temp_b2_14_14_i,temp_m3_10_10_r,temp_m3_10_10_i,temp_m3_10_14_r,temp_m3_10_14_i,temp_m3_14_10_r,temp_m3_14_10_i,temp_m3_14_14_r,temp_m3_14_14_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly598 (clk,temp_m3_10_10_r,temp_m3_10_10_i,temp_m3_10_14_r,temp_m3_10_14_i,temp_m3_14_10_r,temp_m3_14_10_i,temp_m3_14_14_r,temp_m3_14_14_i,temp_b3_10_10_r,temp_b3_10_10_i,temp_b3_10_14_r,temp_b3_10_14_i,temp_b3_14_10_r,temp_b3_14_10_i,temp_b3_14_14_r,temp_b3_14_14_i);
MULT MULT599 (clk,temp_b2_10_11_r,temp_b2_10_11_i,temp_b2_10_15_r,temp_b2_10_15_i,temp_b2_14_11_r,temp_b2_14_11_i,temp_b2_14_15_r,temp_b2_14_15_i,temp_m3_10_11_r,temp_m3_10_11_i,temp_m3_10_15_r,temp_m3_10_15_i,temp_m3_14_11_r,temp_m3_14_11_i,temp_m3_14_15_r,temp_m3_14_15_i,`W8_real,`W8_imag,`W4_real,`W4_imag,`W12_real,`W12_imag);
butterfly butterfly599 (clk,temp_m3_10_11_r,temp_m3_10_11_i,temp_m3_10_15_r,temp_m3_10_15_i,temp_m3_14_11_r,temp_m3_14_11_i,temp_m3_14_15_r,temp_m3_14_15_i,temp_b3_10_11_r,temp_b3_10_11_i,temp_b3_10_15_r,temp_b3_10_15_i,temp_b3_14_11_r,temp_b3_14_11_i,temp_b3_14_15_r,temp_b3_14_15_i);
MULT MULT600 (clk,temp_b2_10_12_r,temp_b2_10_12_i,temp_b2_10_16_r,temp_b2_10_16_i,temp_b2_14_12_r,temp_b2_14_12_i,temp_b2_14_16_r,temp_b2_14_16_i,temp_m3_10_12_r,temp_m3_10_12_i,temp_m3_10_16_r,temp_m3_10_16_i,temp_m3_14_12_r,temp_m3_14_12_i,temp_m3_14_16_r,temp_m3_14_16_i,`W12_real,`W12_imag,`W4_real,`W4_imag,`W16_real,`W16_imag);
butterfly butterfly600 (clk,temp_m3_10_12_r,temp_m3_10_12_i,temp_m3_10_16_r,temp_m3_10_16_i,temp_m3_14_12_r,temp_m3_14_12_i,temp_m3_14_16_r,temp_m3_14_16_i,temp_b3_10_12_r,temp_b3_10_12_i,temp_b3_10_16_r,temp_b3_10_16_i,temp_b3_14_12_r,temp_b3_14_12_i,temp_b3_14_16_r,temp_b3_14_16_i);
MULT MULT601 (clk,temp_b2_11_9_r,temp_b2_11_9_i,temp_b2_11_13_r,temp_b2_11_13_i,temp_b2_15_9_r,temp_b2_15_9_i,temp_b2_15_13_r,temp_b2_15_13_i,temp_m3_11_9_r,temp_m3_11_9_i,temp_m3_11_13_r,temp_m3_11_13_i,temp_m3_15_9_r,temp_m3_15_9_i,temp_m3_15_13_r,temp_m3_15_13_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly601 (clk,temp_m3_11_9_r,temp_m3_11_9_i,temp_m3_11_13_r,temp_m3_11_13_i,temp_m3_15_9_r,temp_m3_15_9_i,temp_m3_15_13_r,temp_m3_15_13_i,temp_b3_11_9_r,temp_b3_11_9_i,temp_b3_11_13_r,temp_b3_11_13_i,temp_b3_15_9_r,temp_b3_15_9_i,temp_b3_15_13_r,temp_b3_15_13_i);
MULT MULT602 (clk,temp_b2_11_10_r,temp_b2_11_10_i,temp_b2_11_14_r,temp_b2_11_14_i,temp_b2_15_10_r,temp_b2_15_10_i,temp_b2_15_14_r,temp_b2_15_14_i,temp_m3_11_10_r,temp_m3_11_10_i,temp_m3_11_14_r,temp_m3_11_14_i,temp_m3_15_10_r,temp_m3_15_10_i,temp_m3_15_14_r,temp_m3_15_14_i,`W4_real,`W4_imag,`W8_real,`W8_imag,`W12_real,`W12_imag);
butterfly butterfly602 (clk,temp_m3_11_10_r,temp_m3_11_10_i,temp_m3_11_14_r,temp_m3_11_14_i,temp_m3_15_10_r,temp_m3_15_10_i,temp_m3_15_14_r,temp_m3_15_14_i,temp_b3_11_10_r,temp_b3_11_10_i,temp_b3_11_14_r,temp_b3_11_14_i,temp_b3_15_10_r,temp_b3_15_10_i,temp_b3_15_14_r,temp_b3_15_14_i);
MULT MULT603 (clk,temp_b2_11_11_r,temp_b2_11_11_i,temp_b2_11_15_r,temp_b2_11_15_i,temp_b2_15_11_r,temp_b2_15_11_i,temp_b2_15_15_r,temp_b2_15_15_i,temp_m3_11_11_r,temp_m3_11_11_i,temp_m3_11_15_r,temp_m3_11_15_i,temp_m3_15_11_r,temp_m3_15_11_i,temp_m3_15_15_r,temp_m3_15_15_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly603 (clk,temp_m3_11_11_r,temp_m3_11_11_i,temp_m3_11_15_r,temp_m3_11_15_i,temp_m3_15_11_r,temp_m3_15_11_i,temp_m3_15_15_r,temp_m3_15_15_i,temp_b3_11_11_r,temp_b3_11_11_i,temp_b3_11_15_r,temp_b3_11_15_i,temp_b3_15_11_r,temp_b3_15_11_i,temp_b3_15_15_r,temp_b3_15_15_i);
MULT MULT604 (clk,temp_b2_11_12_r,temp_b2_11_12_i,temp_b2_11_16_r,temp_b2_11_16_i,temp_b2_15_12_r,temp_b2_15_12_i,temp_b2_15_16_r,temp_b2_15_16_i,temp_m3_11_12_r,temp_m3_11_12_i,temp_m3_11_16_r,temp_m3_11_16_i,temp_m3_15_12_r,temp_m3_15_12_i,temp_m3_15_16_r,temp_m3_15_16_i,`W12_real,`W12_imag,`W8_real,`W8_imag,`W20_real,`W20_imag);
butterfly butterfly604 (clk,temp_m3_11_12_r,temp_m3_11_12_i,temp_m3_11_16_r,temp_m3_11_16_i,temp_m3_15_12_r,temp_m3_15_12_i,temp_m3_15_16_r,temp_m3_15_16_i,temp_b3_11_12_r,temp_b3_11_12_i,temp_b3_11_16_r,temp_b3_11_16_i,temp_b3_15_12_r,temp_b3_15_12_i,temp_b3_15_16_r,temp_b3_15_16_i);
MULT MULT605 (clk,temp_b2_12_9_r,temp_b2_12_9_i,temp_b2_12_13_r,temp_b2_12_13_i,temp_b2_16_9_r,temp_b2_16_9_i,temp_b2_16_13_r,temp_b2_16_13_i,temp_m3_12_9_r,temp_m3_12_9_i,temp_m3_12_13_r,temp_m3_12_13_i,temp_m3_16_9_r,temp_m3_16_9_i,temp_m3_16_13_r,temp_m3_16_13_i,`W0_real,`W0_imag,`W12_real,`W12_imag,`W12_real,`W12_imag);
butterfly butterfly605 (clk,temp_m3_12_9_r,temp_m3_12_9_i,temp_m3_12_13_r,temp_m3_12_13_i,temp_m3_16_9_r,temp_m3_16_9_i,temp_m3_16_13_r,temp_m3_16_13_i,temp_b3_12_9_r,temp_b3_12_9_i,temp_b3_12_13_r,temp_b3_12_13_i,temp_b3_16_9_r,temp_b3_16_9_i,temp_b3_16_13_r,temp_b3_16_13_i);
MULT MULT606 (clk,temp_b2_12_10_r,temp_b2_12_10_i,temp_b2_12_14_r,temp_b2_12_14_i,temp_b2_16_10_r,temp_b2_16_10_i,temp_b2_16_14_r,temp_b2_16_14_i,temp_m3_12_10_r,temp_m3_12_10_i,temp_m3_12_14_r,temp_m3_12_14_i,temp_m3_16_10_r,temp_m3_16_10_i,temp_m3_16_14_r,temp_m3_16_14_i,`W4_real,`W4_imag,`W12_real,`W12_imag,`W16_real,`W16_imag);
butterfly butterfly606 (clk,temp_m3_12_10_r,temp_m3_12_10_i,temp_m3_12_14_r,temp_m3_12_14_i,temp_m3_16_10_r,temp_m3_16_10_i,temp_m3_16_14_r,temp_m3_16_14_i,temp_b3_12_10_r,temp_b3_12_10_i,temp_b3_12_14_r,temp_b3_12_14_i,temp_b3_16_10_r,temp_b3_16_10_i,temp_b3_16_14_r,temp_b3_16_14_i);
MULT MULT607 (clk,temp_b2_12_11_r,temp_b2_12_11_i,temp_b2_12_15_r,temp_b2_12_15_i,temp_b2_16_11_r,temp_b2_16_11_i,temp_b2_16_15_r,temp_b2_16_15_i,temp_m3_12_11_r,temp_m3_12_11_i,temp_m3_12_15_r,temp_m3_12_15_i,temp_m3_16_11_r,temp_m3_16_11_i,temp_m3_16_15_r,temp_m3_16_15_i,`W8_real,`W8_imag,`W12_real,`W12_imag,`W20_real,`W20_imag);
butterfly butterfly607 (clk,temp_m3_12_11_r,temp_m3_12_11_i,temp_m3_12_15_r,temp_m3_12_15_i,temp_m3_16_11_r,temp_m3_16_11_i,temp_m3_16_15_r,temp_m3_16_15_i,temp_b3_12_11_r,temp_b3_12_11_i,temp_b3_12_15_r,temp_b3_12_15_i,temp_b3_16_11_r,temp_b3_16_11_i,temp_b3_16_15_r,temp_b3_16_15_i);
MULT MULT608 (clk,temp_b2_12_12_r,temp_b2_12_12_i,temp_b2_12_16_r,temp_b2_12_16_i,temp_b2_16_12_r,temp_b2_16_12_i,temp_b2_16_16_r,temp_b2_16_16_i,temp_m3_12_12_r,temp_m3_12_12_i,temp_m3_12_16_r,temp_m3_12_16_i,temp_m3_16_12_r,temp_m3_16_12_i,temp_m3_16_16_r,temp_m3_16_16_i,`W12_real,`W12_imag,`W12_real,`W12_imag,`W24_real,`W24_imag);
butterfly butterfly608 (clk,temp_m3_12_12_r,temp_m3_12_12_i,temp_m3_12_16_r,temp_m3_12_16_i,temp_m3_16_12_r,temp_m3_16_12_i,temp_m3_16_16_r,temp_m3_16_16_i,temp_b3_12_12_r,temp_b3_12_12_i,temp_b3_12_16_r,temp_b3_12_16_i,temp_b3_16_12_r,temp_b3_16_12_i,temp_b3_16_16_r,temp_b3_16_16_i);
MULT MULT609 (clk,temp_b2_9_17_r,temp_b2_9_17_i,temp_b2_9_21_r,temp_b2_9_21_i,temp_b2_13_17_r,temp_b2_13_17_i,temp_b2_13_21_r,temp_b2_13_21_i,temp_m3_9_17_r,temp_m3_9_17_i,temp_m3_9_21_r,temp_m3_9_21_i,temp_m3_13_17_r,temp_m3_13_17_i,temp_m3_13_21_r,temp_m3_13_21_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly609 (clk,temp_m3_9_17_r,temp_m3_9_17_i,temp_m3_9_21_r,temp_m3_9_21_i,temp_m3_13_17_r,temp_m3_13_17_i,temp_m3_13_21_r,temp_m3_13_21_i,temp_b3_9_17_r,temp_b3_9_17_i,temp_b3_9_21_r,temp_b3_9_21_i,temp_b3_13_17_r,temp_b3_13_17_i,temp_b3_13_21_r,temp_b3_13_21_i);
MULT MULT610 (clk,temp_b2_9_18_r,temp_b2_9_18_i,temp_b2_9_22_r,temp_b2_9_22_i,temp_b2_13_18_r,temp_b2_13_18_i,temp_b2_13_22_r,temp_b2_13_22_i,temp_m3_9_18_r,temp_m3_9_18_i,temp_m3_9_22_r,temp_m3_9_22_i,temp_m3_13_18_r,temp_m3_13_18_i,temp_m3_13_22_r,temp_m3_13_22_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly610 (clk,temp_m3_9_18_r,temp_m3_9_18_i,temp_m3_9_22_r,temp_m3_9_22_i,temp_m3_13_18_r,temp_m3_13_18_i,temp_m3_13_22_r,temp_m3_13_22_i,temp_b3_9_18_r,temp_b3_9_18_i,temp_b3_9_22_r,temp_b3_9_22_i,temp_b3_13_18_r,temp_b3_13_18_i,temp_b3_13_22_r,temp_b3_13_22_i);
MULT MULT611 (clk,temp_b2_9_19_r,temp_b2_9_19_i,temp_b2_9_23_r,temp_b2_9_23_i,temp_b2_13_19_r,temp_b2_13_19_i,temp_b2_13_23_r,temp_b2_13_23_i,temp_m3_9_19_r,temp_m3_9_19_i,temp_m3_9_23_r,temp_m3_9_23_i,temp_m3_13_19_r,temp_m3_13_19_i,temp_m3_13_23_r,temp_m3_13_23_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly611 (clk,temp_m3_9_19_r,temp_m3_9_19_i,temp_m3_9_23_r,temp_m3_9_23_i,temp_m3_13_19_r,temp_m3_13_19_i,temp_m3_13_23_r,temp_m3_13_23_i,temp_b3_9_19_r,temp_b3_9_19_i,temp_b3_9_23_r,temp_b3_9_23_i,temp_b3_13_19_r,temp_b3_13_19_i,temp_b3_13_23_r,temp_b3_13_23_i);
MULT MULT612 (clk,temp_b2_9_20_r,temp_b2_9_20_i,temp_b2_9_24_r,temp_b2_9_24_i,temp_b2_13_20_r,temp_b2_13_20_i,temp_b2_13_24_r,temp_b2_13_24_i,temp_m3_9_20_r,temp_m3_9_20_i,temp_m3_9_24_r,temp_m3_9_24_i,temp_m3_13_20_r,temp_m3_13_20_i,temp_m3_13_24_r,temp_m3_13_24_i,`W12_real,`W12_imag,`W0_real,`W0_imag,`W12_real,`W12_imag);
butterfly butterfly612 (clk,temp_m3_9_20_r,temp_m3_9_20_i,temp_m3_9_24_r,temp_m3_9_24_i,temp_m3_13_20_r,temp_m3_13_20_i,temp_m3_13_24_r,temp_m3_13_24_i,temp_b3_9_20_r,temp_b3_9_20_i,temp_b3_9_24_r,temp_b3_9_24_i,temp_b3_13_20_r,temp_b3_13_20_i,temp_b3_13_24_r,temp_b3_13_24_i);
MULT MULT613 (clk,temp_b2_10_17_r,temp_b2_10_17_i,temp_b2_10_21_r,temp_b2_10_21_i,temp_b2_14_17_r,temp_b2_14_17_i,temp_b2_14_21_r,temp_b2_14_21_i,temp_m3_10_17_r,temp_m3_10_17_i,temp_m3_10_21_r,temp_m3_10_21_i,temp_m3_14_17_r,temp_m3_14_17_i,temp_m3_14_21_r,temp_m3_14_21_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly613 (clk,temp_m3_10_17_r,temp_m3_10_17_i,temp_m3_10_21_r,temp_m3_10_21_i,temp_m3_14_17_r,temp_m3_14_17_i,temp_m3_14_21_r,temp_m3_14_21_i,temp_b3_10_17_r,temp_b3_10_17_i,temp_b3_10_21_r,temp_b3_10_21_i,temp_b3_14_17_r,temp_b3_14_17_i,temp_b3_14_21_r,temp_b3_14_21_i);
MULT MULT614 (clk,temp_b2_10_18_r,temp_b2_10_18_i,temp_b2_10_22_r,temp_b2_10_22_i,temp_b2_14_18_r,temp_b2_14_18_i,temp_b2_14_22_r,temp_b2_14_22_i,temp_m3_10_18_r,temp_m3_10_18_i,temp_m3_10_22_r,temp_m3_10_22_i,temp_m3_14_18_r,temp_m3_14_18_i,temp_m3_14_22_r,temp_m3_14_22_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly614 (clk,temp_m3_10_18_r,temp_m3_10_18_i,temp_m3_10_22_r,temp_m3_10_22_i,temp_m3_14_18_r,temp_m3_14_18_i,temp_m3_14_22_r,temp_m3_14_22_i,temp_b3_10_18_r,temp_b3_10_18_i,temp_b3_10_22_r,temp_b3_10_22_i,temp_b3_14_18_r,temp_b3_14_18_i,temp_b3_14_22_r,temp_b3_14_22_i);
MULT MULT615 (clk,temp_b2_10_19_r,temp_b2_10_19_i,temp_b2_10_23_r,temp_b2_10_23_i,temp_b2_14_19_r,temp_b2_14_19_i,temp_b2_14_23_r,temp_b2_14_23_i,temp_m3_10_19_r,temp_m3_10_19_i,temp_m3_10_23_r,temp_m3_10_23_i,temp_m3_14_19_r,temp_m3_14_19_i,temp_m3_14_23_r,temp_m3_14_23_i,`W8_real,`W8_imag,`W4_real,`W4_imag,`W12_real,`W12_imag);
butterfly butterfly615 (clk,temp_m3_10_19_r,temp_m3_10_19_i,temp_m3_10_23_r,temp_m3_10_23_i,temp_m3_14_19_r,temp_m3_14_19_i,temp_m3_14_23_r,temp_m3_14_23_i,temp_b3_10_19_r,temp_b3_10_19_i,temp_b3_10_23_r,temp_b3_10_23_i,temp_b3_14_19_r,temp_b3_14_19_i,temp_b3_14_23_r,temp_b3_14_23_i);
MULT MULT616 (clk,temp_b2_10_20_r,temp_b2_10_20_i,temp_b2_10_24_r,temp_b2_10_24_i,temp_b2_14_20_r,temp_b2_14_20_i,temp_b2_14_24_r,temp_b2_14_24_i,temp_m3_10_20_r,temp_m3_10_20_i,temp_m3_10_24_r,temp_m3_10_24_i,temp_m3_14_20_r,temp_m3_14_20_i,temp_m3_14_24_r,temp_m3_14_24_i,`W12_real,`W12_imag,`W4_real,`W4_imag,`W16_real,`W16_imag);
butterfly butterfly616 (clk,temp_m3_10_20_r,temp_m3_10_20_i,temp_m3_10_24_r,temp_m3_10_24_i,temp_m3_14_20_r,temp_m3_14_20_i,temp_m3_14_24_r,temp_m3_14_24_i,temp_b3_10_20_r,temp_b3_10_20_i,temp_b3_10_24_r,temp_b3_10_24_i,temp_b3_14_20_r,temp_b3_14_20_i,temp_b3_14_24_r,temp_b3_14_24_i);
MULT MULT617 (clk,temp_b2_11_17_r,temp_b2_11_17_i,temp_b2_11_21_r,temp_b2_11_21_i,temp_b2_15_17_r,temp_b2_15_17_i,temp_b2_15_21_r,temp_b2_15_21_i,temp_m3_11_17_r,temp_m3_11_17_i,temp_m3_11_21_r,temp_m3_11_21_i,temp_m3_15_17_r,temp_m3_15_17_i,temp_m3_15_21_r,temp_m3_15_21_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly617 (clk,temp_m3_11_17_r,temp_m3_11_17_i,temp_m3_11_21_r,temp_m3_11_21_i,temp_m3_15_17_r,temp_m3_15_17_i,temp_m3_15_21_r,temp_m3_15_21_i,temp_b3_11_17_r,temp_b3_11_17_i,temp_b3_11_21_r,temp_b3_11_21_i,temp_b3_15_17_r,temp_b3_15_17_i,temp_b3_15_21_r,temp_b3_15_21_i);
MULT MULT618 (clk,temp_b2_11_18_r,temp_b2_11_18_i,temp_b2_11_22_r,temp_b2_11_22_i,temp_b2_15_18_r,temp_b2_15_18_i,temp_b2_15_22_r,temp_b2_15_22_i,temp_m3_11_18_r,temp_m3_11_18_i,temp_m3_11_22_r,temp_m3_11_22_i,temp_m3_15_18_r,temp_m3_15_18_i,temp_m3_15_22_r,temp_m3_15_22_i,`W4_real,`W4_imag,`W8_real,`W8_imag,`W12_real,`W12_imag);
butterfly butterfly618 (clk,temp_m3_11_18_r,temp_m3_11_18_i,temp_m3_11_22_r,temp_m3_11_22_i,temp_m3_15_18_r,temp_m3_15_18_i,temp_m3_15_22_r,temp_m3_15_22_i,temp_b3_11_18_r,temp_b3_11_18_i,temp_b3_11_22_r,temp_b3_11_22_i,temp_b3_15_18_r,temp_b3_15_18_i,temp_b3_15_22_r,temp_b3_15_22_i);
MULT MULT619 (clk,temp_b2_11_19_r,temp_b2_11_19_i,temp_b2_11_23_r,temp_b2_11_23_i,temp_b2_15_19_r,temp_b2_15_19_i,temp_b2_15_23_r,temp_b2_15_23_i,temp_m3_11_19_r,temp_m3_11_19_i,temp_m3_11_23_r,temp_m3_11_23_i,temp_m3_15_19_r,temp_m3_15_19_i,temp_m3_15_23_r,temp_m3_15_23_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly619 (clk,temp_m3_11_19_r,temp_m3_11_19_i,temp_m3_11_23_r,temp_m3_11_23_i,temp_m3_15_19_r,temp_m3_15_19_i,temp_m3_15_23_r,temp_m3_15_23_i,temp_b3_11_19_r,temp_b3_11_19_i,temp_b3_11_23_r,temp_b3_11_23_i,temp_b3_15_19_r,temp_b3_15_19_i,temp_b3_15_23_r,temp_b3_15_23_i);
MULT MULT620 (clk,temp_b2_11_20_r,temp_b2_11_20_i,temp_b2_11_24_r,temp_b2_11_24_i,temp_b2_15_20_r,temp_b2_15_20_i,temp_b2_15_24_r,temp_b2_15_24_i,temp_m3_11_20_r,temp_m3_11_20_i,temp_m3_11_24_r,temp_m3_11_24_i,temp_m3_15_20_r,temp_m3_15_20_i,temp_m3_15_24_r,temp_m3_15_24_i,`W12_real,`W12_imag,`W8_real,`W8_imag,`W20_real,`W20_imag);
butterfly butterfly620 (clk,temp_m3_11_20_r,temp_m3_11_20_i,temp_m3_11_24_r,temp_m3_11_24_i,temp_m3_15_20_r,temp_m3_15_20_i,temp_m3_15_24_r,temp_m3_15_24_i,temp_b3_11_20_r,temp_b3_11_20_i,temp_b3_11_24_r,temp_b3_11_24_i,temp_b3_15_20_r,temp_b3_15_20_i,temp_b3_15_24_r,temp_b3_15_24_i);
MULT MULT621 (clk,temp_b2_12_17_r,temp_b2_12_17_i,temp_b2_12_21_r,temp_b2_12_21_i,temp_b2_16_17_r,temp_b2_16_17_i,temp_b2_16_21_r,temp_b2_16_21_i,temp_m3_12_17_r,temp_m3_12_17_i,temp_m3_12_21_r,temp_m3_12_21_i,temp_m3_16_17_r,temp_m3_16_17_i,temp_m3_16_21_r,temp_m3_16_21_i,`W0_real,`W0_imag,`W12_real,`W12_imag,`W12_real,`W12_imag);
butterfly butterfly621 (clk,temp_m3_12_17_r,temp_m3_12_17_i,temp_m3_12_21_r,temp_m3_12_21_i,temp_m3_16_17_r,temp_m3_16_17_i,temp_m3_16_21_r,temp_m3_16_21_i,temp_b3_12_17_r,temp_b3_12_17_i,temp_b3_12_21_r,temp_b3_12_21_i,temp_b3_16_17_r,temp_b3_16_17_i,temp_b3_16_21_r,temp_b3_16_21_i);
MULT MULT622 (clk,temp_b2_12_18_r,temp_b2_12_18_i,temp_b2_12_22_r,temp_b2_12_22_i,temp_b2_16_18_r,temp_b2_16_18_i,temp_b2_16_22_r,temp_b2_16_22_i,temp_m3_12_18_r,temp_m3_12_18_i,temp_m3_12_22_r,temp_m3_12_22_i,temp_m3_16_18_r,temp_m3_16_18_i,temp_m3_16_22_r,temp_m3_16_22_i,`W4_real,`W4_imag,`W12_real,`W12_imag,`W16_real,`W16_imag);
butterfly butterfly622 (clk,temp_m3_12_18_r,temp_m3_12_18_i,temp_m3_12_22_r,temp_m3_12_22_i,temp_m3_16_18_r,temp_m3_16_18_i,temp_m3_16_22_r,temp_m3_16_22_i,temp_b3_12_18_r,temp_b3_12_18_i,temp_b3_12_22_r,temp_b3_12_22_i,temp_b3_16_18_r,temp_b3_16_18_i,temp_b3_16_22_r,temp_b3_16_22_i);
MULT MULT623 (clk,temp_b2_12_19_r,temp_b2_12_19_i,temp_b2_12_23_r,temp_b2_12_23_i,temp_b2_16_19_r,temp_b2_16_19_i,temp_b2_16_23_r,temp_b2_16_23_i,temp_m3_12_19_r,temp_m3_12_19_i,temp_m3_12_23_r,temp_m3_12_23_i,temp_m3_16_19_r,temp_m3_16_19_i,temp_m3_16_23_r,temp_m3_16_23_i,`W8_real,`W8_imag,`W12_real,`W12_imag,`W20_real,`W20_imag);
butterfly butterfly623 (clk,temp_m3_12_19_r,temp_m3_12_19_i,temp_m3_12_23_r,temp_m3_12_23_i,temp_m3_16_19_r,temp_m3_16_19_i,temp_m3_16_23_r,temp_m3_16_23_i,temp_b3_12_19_r,temp_b3_12_19_i,temp_b3_12_23_r,temp_b3_12_23_i,temp_b3_16_19_r,temp_b3_16_19_i,temp_b3_16_23_r,temp_b3_16_23_i);
MULT MULT624 (clk,temp_b2_12_20_r,temp_b2_12_20_i,temp_b2_12_24_r,temp_b2_12_24_i,temp_b2_16_20_r,temp_b2_16_20_i,temp_b2_16_24_r,temp_b2_16_24_i,temp_m3_12_20_r,temp_m3_12_20_i,temp_m3_12_24_r,temp_m3_12_24_i,temp_m3_16_20_r,temp_m3_16_20_i,temp_m3_16_24_r,temp_m3_16_24_i,`W12_real,`W12_imag,`W12_real,`W12_imag,`W24_real,`W24_imag);
butterfly butterfly624 (clk,temp_m3_12_20_r,temp_m3_12_20_i,temp_m3_12_24_r,temp_m3_12_24_i,temp_m3_16_20_r,temp_m3_16_20_i,temp_m3_16_24_r,temp_m3_16_24_i,temp_b3_12_20_r,temp_b3_12_20_i,temp_b3_12_24_r,temp_b3_12_24_i,temp_b3_16_20_r,temp_b3_16_20_i,temp_b3_16_24_r,temp_b3_16_24_i);
MULT MULT625 (clk,temp_b2_9_25_r,temp_b2_9_25_i,temp_b2_9_29_r,temp_b2_9_29_i,temp_b2_13_25_r,temp_b2_13_25_i,temp_b2_13_29_r,temp_b2_13_29_i,temp_m3_9_25_r,temp_m3_9_25_i,temp_m3_9_29_r,temp_m3_9_29_i,temp_m3_13_25_r,temp_m3_13_25_i,temp_m3_13_29_r,temp_m3_13_29_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly625 (clk,temp_m3_9_25_r,temp_m3_9_25_i,temp_m3_9_29_r,temp_m3_9_29_i,temp_m3_13_25_r,temp_m3_13_25_i,temp_m3_13_29_r,temp_m3_13_29_i,temp_b3_9_25_r,temp_b3_9_25_i,temp_b3_9_29_r,temp_b3_9_29_i,temp_b3_13_25_r,temp_b3_13_25_i,temp_b3_13_29_r,temp_b3_13_29_i);
MULT MULT626 (clk,temp_b2_9_26_r,temp_b2_9_26_i,temp_b2_9_30_r,temp_b2_9_30_i,temp_b2_13_26_r,temp_b2_13_26_i,temp_b2_13_30_r,temp_b2_13_30_i,temp_m3_9_26_r,temp_m3_9_26_i,temp_m3_9_30_r,temp_m3_9_30_i,temp_m3_13_26_r,temp_m3_13_26_i,temp_m3_13_30_r,temp_m3_13_30_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly626 (clk,temp_m3_9_26_r,temp_m3_9_26_i,temp_m3_9_30_r,temp_m3_9_30_i,temp_m3_13_26_r,temp_m3_13_26_i,temp_m3_13_30_r,temp_m3_13_30_i,temp_b3_9_26_r,temp_b3_9_26_i,temp_b3_9_30_r,temp_b3_9_30_i,temp_b3_13_26_r,temp_b3_13_26_i,temp_b3_13_30_r,temp_b3_13_30_i);
MULT MULT627 (clk,temp_b2_9_27_r,temp_b2_9_27_i,temp_b2_9_31_r,temp_b2_9_31_i,temp_b2_13_27_r,temp_b2_13_27_i,temp_b2_13_31_r,temp_b2_13_31_i,temp_m3_9_27_r,temp_m3_9_27_i,temp_m3_9_31_r,temp_m3_9_31_i,temp_m3_13_27_r,temp_m3_13_27_i,temp_m3_13_31_r,temp_m3_13_31_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly627 (clk,temp_m3_9_27_r,temp_m3_9_27_i,temp_m3_9_31_r,temp_m3_9_31_i,temp_m3_13_27_r,temp_m3_13_27_i,temp_m3_13_31_r,temp_m3_13_31_i,temp_b3_9_27_r,temp_b3_9_27_i,temp_b3_9_31_r,temp_b3_9_31_i,temp_b3_13_27_r,temp_b3_13_27_i,temp_b3_13_31_r,temp_b3_13_31_i);
MULT MULT628 (clk,temp_b2_9_28_r,temp_b2_9_28_i,temp_b2_9_32_r,temp_b2_9_32_i,temp_b2_13_28_r,temp_b2_13_28_i,temp_b2_13_32_r,temp_b2_13_32_i,temp_m3_9_28_r,temp_m3_9_28_i,temp_m3_9_32_r,temp_m3_9_32_i,temp_m3_13_28_r,temp_m3_13_28_i,temp_m3_13_32_r,temp_m3_13_32_i,`W12_real,`W12_imag,`W0_real,`W0_imag,`W12_real,`W12_imag);
butterfly butterfly628 (clk,temp_m3_9_28_r,temp_m3_9_28_i,temp_m3_9_32_r,temp_m3_9_32_i,temp_m3_13_28_r,temp_m3_13_28_i,temp_m3_13_32_r,temp_m3_13_32_i,temp_b3_9_28_r,temp_b3_9_28_i,temp_b3_9_32_r,temp_b3_9_32_i,temp_b3_13_28_r,temp_b3_13_28_i,temp_b3_13_32_r,temp_b3_13_32_i);
MULT MULT629 (clk,temp_b2_10_25_r,temp_b2_10_25_i,temp_b2_10_29_r,temp_b2_10_29_i,temp_b2_14_25_r,temp_b2_14_25_i,temp_b2_14_29_r,temp_b2_14_29_i,temp_m3_10_25_r,temp_m3_10_25_i,temp_m3_10_29_r,temp_m3_10_29_i,temp_m3_14_25_r,temp_m3_14_25_i,temp_m3_14_29_r,temp_m3_14_29_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly629 (clk,temp_m3_10_25_r,temp_m3_10_25_i,temp_m3_10_29_r,temp_m3_10_29_i,temp_m3_14_25_r,temp_m3_14_25_i,temp_m3_14_29_r,temp_m3_14_29_i,temp_b3_10_25_r,temp_b3_10_25_i,temp_b3_10_29_r,temp_b3_10_29_i,temp_b3_14_25_r,temp_b3_14_25_i,temp_b3_14_29_r,temp_b3_14_29_i);
MULT MULT630 (clk,temp_b2_10_26_r,temp_b2_10_26_i,temp_b2_10_30_r,temp_b2_10_30_i,temp_b2_14_26_r,temp_b2_14_26_i,temp_b2_14_30_r,temp_b2_14_30_i,temp_m3_10_26_r,temp_m3_10_26_i,temp_m3_10_30_r,temp_m3_10_30_i,temp_m3_14_26_r,temp_m3_14_26_i,temp_m3_14_30_r,temp_m3_14_30_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly630 (clk,temp_m3_10_26_r,temp_m3_10_26_i,temp_m3_10_30_r,temp_m3_10_30_i,temp_m3_14_26_r,temp_m3_14_26_i,temp_m3_14_30_r,temp_m3_14_30_i,temp_b3_10_26_r,temp_b3_10_26_i,temp_b3_10_30_r,temp_b3_10_30_i,temp_b3_14_26_r,temp_b3_14_26_i,temp_b3_14_30_r,temp_b3_14_30_i);
MULT MULT631 (clk,temp_b2_10_27_r,temp_b2_10_27_i,temp_b2_10_31_r,temp_b2_10_31_i,temp_b2_14_27_r,temp_b2_14_27_i,temp_b2_14_31_r,temp_b2_14_31_i,temp_m3_10_27_r,temp_m3_10_27_i,temp_m3_10_31_r,temp_m3_10_31_i,temp_m3_14_27_r,temp_m3_14_27_i,temp_m3_14_31_r,temp_m3_14_31_i,`W8_real,`W8_imag,`W4_real,`W4_imag,`W12_real,`W12_imag);
butterfly butterfly631 (clk,temp_m3_10_27_r,temp_m3_10_27_i,temp_m3_10_31_r,temp_m3_10_31_i,temp_m3_14_27_r,temp_m3_14_27_i,temp_m3_14_31_r,temp_m3_14_31_i,temp_b3_10_27_r,temp_b3_10_27_i,temp_b3_10_31_r,temp_b3_10_31_i,temp_b3_14_27_r,temp_b3_14_27_i,temp_b3_14_31_r,temp_b3_14_31_i);
MULT MULT632 (clk,temp_b2_10_28_r,temp_b2_10_28_i,temp_b2_10_32_r,temp_b2_10_32_i,temp_b2_14_28_r,temp_b2_14_28_i,temp_b2_14_32_r,temp_b2_14_32_i,temp_m3_10_28_r,temp_m3_10_28_i,temp_m3_10_32_r,temp_m3_10_32_i,temp_m3_14_28_r,temp_m3_14_28_i,temp_m3_14_32_r,temp_m3_14_32_i,`W12_real,`W12_imag,`W4_real,`W4_imag,`W16_real,`W16_imag);
butterfly butterfly632 (clk,temp_m3_10_28_r,temp_m3_10_28_i,temp_m3_10_32_r,temp_m3_10_32_i,temp_m3_14_28_r,temp_m3_14_28_i,temp_m3_14_32_r,temp_m3_14_32_i,temp_b3_10_28_r,temp_b3_10_28_i,temp_b3_10_32_r,temp_b3_10_32_i,temp_b3_14_28_r,temp_b3_14_28_i,temp_b3_14_32_r,temp_b3_14_32_i);
MULT MULT633 (clk,temp_b2_11_25_r,temp_b2_11_25_i,temp_b2_11_29_r,temp_b2_11_29_i,temp_b2_15_25_r,temp_b2_15_25_i,temp_b2_15_29_r,temp_b2_15_29_i,temp_m3_11_25_r,temp_m3_11_25_i,temp_m3_11_29_r,temp_m3_11_29_i,temp_m3_15_25_r,temp_m3_15_25_i,temp_m3_15_29_r,temp_m3_15_29_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly633 (clk,temp_m3_11_25_r,temp_m3_11_25_i,temp_m3_11_29_r,temp_m3_11_29_i,temp_m3_15_25_r,temp_m3_15_25_i,temp_m3_15_29_r,temp_m3_15_29_i,temp_b3_11_25_r,temp_b3_11_25_i,temp_b3_11_29_r,temp_b3_11_29_i,temp_b3_15_25_r,temp_b3_15_25_i,temp_b3_15_29_r,temp_b3_15_29_i);
MULT MULT634 (clk,temp_b2_11_26_r,temp_b2_11_26_i,temp_b2_11_30_r,temp_b2_11_30_i,temp_b2_15_26_r,temp_b2_15_26_i,temp_b2_15_30_r,temp_b2_15_30_i,temp_m3_11_26_r,temp_m3_11_26_i,temp_m3_11_30_r,temp_m3_11_30_i,temp_m3_15_26_r,temp_m3_15_26_i,temp_m3_15_30_r,temp_m3_15_30_i,`W4_real,`W4_imag,`W8_real,`W8_imag,`W12_real,`W12_imag);
butterfly butterfly634 (clk,temp_m3_11_26_r,temp_m3_11_26_i,temp_m3_11_30_r,temp_m3_11_30_i,temp_m3_15_26_r,temp_m3_15_26_i,temp_m3_15_30_r,temp_m3_15_30_i,temp_b3_11_26_r,temp_b3_11_26_i,temp_b3_11_30_r,temp_b3_11_30_i,temp_b3_15_26_r,temp_b3_15_26_i,temp_b3_15_30_r,temp_b3_15_30_i);
MULT MULT635 (clk,temp_b2_11_27_r,temp_b2_11_27_i,temp_b2_11_31_r,temp_b2_11_31_i,temp_b2_15_27_r,temp_b2_15_27_i,temp_b2_15_31_r,temp_b2_15_31_i,temp_m3_11_27_r,temp_m3_11_27_i,temp_m3_11_31_r,temp_m3_11_31_i,temp_m3_15_27_r,temp_m3_15_27_i,temp_m3_15_31_r,temp_m3_15_31_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly635 (clk,temp_m3_11_27_r,temp_m3_11_27_i,temp_m3_11_31_r,temp_m3_11_31_i,temp_m3_15_27_r,temp_m3_15_27_i,temp_m3_15_31_r,temp_m3_15_31_i,temp_b3_11_27_r,temp_b3_11_27_i,temp_b3_11_31_r,temp_b3_11_31_i,temp_b3_15_27_r,temp_b3_15_27_i,temp_b3_15_31_r,temp_b3_15_31_i);
MULT MULT636 (clk,temp_b2_11_28_r,temp_b2_11_28_i,temp_b2_11_32_r,temp_b2_11_32_i,temp_b2_15_28_r,temp_b2_15_28_i,temp_b2_15_32_r,temp_b2_15_32_i,temp_m3_11_28_r,temp_m3_11_28_i,temp_m3_11_32_r,temp_m3_11_32_i,temp_m3_15_28_r,temp_m3_15_28_i,temp_m3_15_32_r,temp_m3_15_32_i,`W12_real,`W12_imag,`W8_real,`W8_imag,`W20_real,`W20_imag);
butterfly butterfly636 (clk,temp_m3_11_28_r,temp_m3_11_28_i,temp_m3_11_32_r,temp_m3_11_32_i,temp_m3_15_28_r,temp_m3_15_28_i,temp_m3_15_32_r,temp_m3_15_32_i,temp_b3_11_28_r,temp_b3_11_28_i,temp_b3_11_32_r,temp_b3_11_32_i,temp_b3_15_28_r,temp_b3_15_28_i,temp_b3_15_32_r,temp_b3_15_32_i);
MULT MULT637 (clk,temp_b2_12_25_r,temp_b2_12_25_i,temp_b2_12_29_r,temp_b2_12_29_i,temp_b2_16_25_r,temp_b2_16_25_i,temp_b2_16_29_r,temp_b2_16_29_i,temp_m3_12_25_r,temp_m3_12_25_i,temp_m3_12_29_r,temp_m3_12_29_i,temp_m3_16_25_r,temp_m3_16_25_i,temp_m3_16_29_r,temp_m3_16_29_i,`W0_real,`W0_imag,`W12_real,`W12_imag,`W12_real,`W12_imag);
butterfly butterfly637 (clk,temp_m3_12_25_r,temp_m3_12_25_i,temp_m3_12_29_r,temp_m3_12_29_i,temp_m3_16_25_r,temp_m3_16_25_i,temp_m3_16_29_r,temp_m3_16_29_i,temp_b3_12_25_r,temp_b3_12_25_i,temp_b3_12_29_r,temp_b3_12_29_i,temp_b3_16_25_r,temp_b3_16_25_i,temp_b3_16_29_r,temp_b3_16_29_i);
MULT MULT638 (clk,temp_b2_12_26_r,temp_b2_12_26_i,temp_b2_12_30_r,temp_b2_12_30_i,temp_b2_16_26_r,temp_b2_16_26_i,temp_b2_16_30_r,temp_b2_16_30_i,temp_m3_12_26_r,temp_m3_12_26_i,temp_m3_12_30_r,temp_m3_12_30_i,temp_m3_16_26_r,temp_m3_16_26_i,temp_m3_16_30_r,temp_m3_16_30_i,`W4_real,`W4_imag,`W12_real,`W12_imag,`W16_real,`W16_imag);
butterfly butterfly638 (clk,temp_m3_12_26_r,temp_m3_12_26_i,temp_m3_12_30_r,temp_m3_12_30_i,temp_m3_16_26_r,temp_m3_16_26_i,temp_m3_16_30_r,temp_m3_16_30_i,temp_b3_12_26_r,temp_b3_12_26_i,temp_b3_12_30_r,temp_b3_12_30_i,temp_b3_16_26_r,temp_b3_16_26_i,temp_b3_16_30_r,temp_b3_16_30_i);
MULT MULT639 (clk,temp_b2_12_27_r,temp_b2_12_27_i,temp_b2_12_31_r,temp_b2_12_31_i,temp_b2_16_27_r,temp_b2_16_27_i,temp_b2_16_31_r,temp_b2_16_31_i,temp_m3_12_27_r,temp_m3_12_27_i,temp_m3_12_31_r,temp_m3_12_31_i,temp_m3_16_27_r,temp_m3_16_27_i,temp_m3_16_31_r,temp_m3_16_31_i,`W8_real,`W8_imag,`W12_real,`W12_imag,`W20_real,`W20_imag);
butterfly butterfly639 (clk,temp_m3_12_27_r,temp_m3_12_27_i,temp_m3_12_31_r,temp_m3_12_31_i,temp_m3_16_27_r,temp_m3_16_27_i,temp_m3_16_31_r,temp_m3_16_31_i,temp_b3_12_27_r,temp_b3_12_27_i,temp_b3_12_31_r,temp_b3_12_31_i,temp_b3_16_27_r,temp_b3_16_27_i,temp_b3_16_31_r,temp_b3_16_31_i);
MULT MULT640 (clk,temp_b2_12_28_r,temp_b2_12_28_i,temp_b2_12_32_r,temp_b2_12_32_i,temp_b2_16_28_r,temp_b2_16_28_i,temp_b2_16_32_r,temp_b2_16_32_i,temp_m3_12_28_r,temp_m3_12_28_i,temp_m3_12_32_r,temp_m3_12_32_i,temp_m3_16_28_r,temp_m3_16_28_i,temp_m3_16_32_r,temp_m3_16_32_i,`W12_real,`W12_imag,`W12_real,`W12_imag,`W24_real,`W24_imag);
butterfly butterfly640 (clk,temp_m3_12_28_r,temp_m3_12_28_i,temp_m3_12_32_r,temp_m3_12_32_i,temp_m3_16_28_r,temp_m3_16_28_i,temp_m3_16_32_r,temp_m3_16_32_i,temp_b3_12_28_r,temp_b3_12_28_i,temp_b3_12_32_r,temp_b3_12_32_i,temp_b3_16_28_r,temp_b3_16_28_i,temp_b3_16_32_r,temp_b3_16_32_i);
MULT MULT641 (clk,temp_b2_17_1_r,temp_b2_17_1_i,temp_b2_17_5_r,temp_b2_17_5_i,temp_b2_21_1_r,temp_b2_21_1_i,temp_b2_21_5_r,temp_b2_21_5_i,temp_m3_17_1_r,temp_m3_17_1_i,temp_m3_17_5_r,temp_m3_17_5_i,temp_m3_21_1_r,temp_m3_21_1_i,temp_m3_21_5_r,temp_m3_21_5_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly641 (clk,temp_m3_17_1_r,temp_m3_17_1_i,temp_m3_17_5_r,temp_m3_17_5_i,temp_m3_21_1_r,temp_m3_21_1_i,temp_m3_21_5_r,temp_m3_21_5_i,temp_b3_17_1_r,temp_b3_17_1_i,temp_b3_17_5_r,temp_b3_17_5_i,temp_b3_21_1_r,temp_b3_21_1_i,temp_b3_21_5_r,temp_b3_21_5_i);
MULT MULT642 (clk,temp_b2_17_2_r,temp_b2_17_2_i,temp_b2_17_6_r,temp_b2_17_6_i,temp_b2_21_2_r,temp_b2_21_2_i,temp_b2_21_6_r,temp_b2_21_6_i,temp_m3_17_2_r,temp_m3_17_2_i,temp_m3_17_6_r,temp_m3_17_6_i,temp_m3_21_2_r,temp_m3_21_2_i,temp_m3_21_6_r,temp_m3_21_6_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly642 (clk,temp_m3_17_2_r,temp_m3_17_2_i,temp_m3_17_6_r,temp_m3_17_6_i,temp_m3_21_2_r,temp_m3_21_2_i,temp_m3_21_6_r,temp_m3_21_6_i,temp_b3_17_2_r,temp_b3_17_2_i,temp_b3_17_6_r,temp_b3_17_6_i,temp_b3_21_2_r,temp_b3_21_2_i,temp_b3_21_6_r,temp_b3_21_6_i);
MULT MULT643 (clk,temp_b2_17_3_r,temp_b2_17_3_i,temp_b2_17_7_r,temp_b2_17_7_i,temp_b2_21_3_r,temp_b2_21_3_i,temp_b2_21_7_r,temp_b2_21_7_i,temp_m3_17_3_r,temp_m3_17_3_i,temp_m3_17_7_r,temp_m3_17_7_i,temp_m3_21_3_r,temp_m3_21_3_i,temp_m3_21_7_r,temp_m3_21_7_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly643 (clk,temp_m3_17_3_r,temp_m3_17_3_i,temp_m3_17_7_r,temp_m3_17_7_i,temp_m3_21_3_r,temp_m3_21_3_i,temp_m3_21_7_r,temp_m3_21_7_i,temp_b3_17_3_r,temp_b3_17_3_i,temp_b3_17_7_r,temp_b3_17_7_i,temp_b3_21_3_r,temp_b3_21_3_i,temp_b3_21_7_r,temp_b3_21_7_i);
MULT MULT644 (clk,temp_b2_17_4_r,temp_b2_17_4_i,temp_b2_17_8_r,temp_b2_17_8_i,temp_b2_21_4_r,temp_b2_21_4_i,temp_b2_21_8_r,temp_b2_21_8_i,temp_m3_17_4_r,temp_m3_17_4_i,temp_m3_17_8_r,temp_m3_17_8_i,temp_m3_21_4_r,temp_m3_21_4_i,temp_m3_21_8_r,temp_m3_21_8_i,`W12_real,`W12_imag,`W0_real,`W0_imag,`W12_real,`W12_imag);
butterfly butterfly644 (clk,temp_m3_17_4_r,temp_m3_17_4_i,temp_m3_17_8_r,temp_m3_17_8_i,temp_m3_21_4_r,temp_m3_21_4_i,temp_m3_21_8_r,temp_m3_21_8_i,temp_b3_17_4_r,temp_b3_17_4_i,temp_b3_17_8_r,temp_b3_17_8_i,temp_b3_21_4_r,temp_b3_21_4_i,temp_b3_21_8_r,temp_b3_21_8_i);
MULT MULT645 (clk,temp_b2_18_1_r,temp_b2_18_1_i,temp_b2_18_5_r,temp_b2_18_5_i,temp_b2_22_1_r,temp_b2_22_1_i,temp_b2_22_5_r,temp_b2_22_5_i,temp_m3_18_1_r,temp_m3_18_1_i,temp_m3_18_5_r,temp_m3_18_5_i,temp_m3_22_1_r,temp_m3_22_1_i,temp_m3_22_5_r,temp_m3_22_5_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly645 (clk,temp_m3_18_1_r,temp_m3_18_1_i,temp_m3_18_5_r,temp_m3_18_5_i,temp_m3_22_1_r,temp_m3_22_1_i,temp_m3_22_5_r,temp_m3_22_5_i,temp_b3_18_1_r,temp_b3_18_1_i,temp_b3_18_5_r,temp_b3_18_5_i,temp_b3_22_1_r,temp_b3_22_1_i,temp_b3_22_5_r,temp_b3_22_5_i);
MULT MULT646 (clk,temp_b2_18_2_r,temp_b2_18_2_i,temp_b2_18_6_r,temp_b2_18_6_i,temp_b2_22_2_r,temp_b2_22_2_i,temp_b2_22_6_r,temp_b2_22_6_i,temp_m3_18_2_r,temp_m3_18_2_i,temp_m3_18_6_r,temp_m3_18_6_i,temp_m3_22_2_r,temp_m3_22_2_i,temp_m3_22_6_r,temp_m3_22_6_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly646 (clk,temp_m3_18_2_r,temp_m3_18_2_i,temp_m3_18_6_r,temp_m3_18_6_i,temp_m3_22_2_r,temp_m3_22_2_i,temp_m3_22_6_r,temp_m3_22_6_i,temp_b3_18_2_r,temp_b3_18_2_i,temp_b3_18_6_r,temp_b3_18_6_i,temp_b3_22_2_r,temp_b3_22_2_i,temp_b3_22_6_r,temp_b3_22_6_i);
MULT MULT647 (clk,temp_b2_18_3_r,temp_b2_18_3_i,temp_b2_18_7_r,temp_b2_18_7_i,temp_b2_22_3_r,temp_b2_22_3_i,temp_b2_22_7_r,temp_b2_22_7_i,temp_m3_18_3_r,temp_m3_18_3_i,temp_m3_18_7_r,temp_m3_18_7_i,temp_m3_22_3_r,temp_m3_22_3_i,temp_m3_22_7_r,temp_m3_22_7_i,`W8_real,`W8_imag,`W4_real,`W4_imag,`W12_real,`W12_imag);
butterfly butterfly647 (clk,temp_m3_18_3_r,temp_m3_18_3_i,temp_m3_18_7_r,temp_m3_18_7_i,temp_m3_22_3_r,temp_m3_22_3_i,temp_m3_22_7_r,temp_m3_22_7_i,temp_b3_18_3_r,temp_b3_18_3_i,temp_b3_18_7_r,temp_b3_18_7_i,temp_b3_22_3_r,temp_b3_22_3_i,temp_b3_22_7_r,temp_b3_22_7_i);
MULT MULT648 (clk,temp_b2_18_4_r,temp_b2_18_4_i,temp_b2_18_8_r,temp_b2_18_8_i,temp_b2_22_4_r,temp_b2_22_4_i,temp_b2_22_8_r,temp_b2_22_8_i,temp_m3_18_4_r,temp_m3_18_4_i,temp_m3_18_8_r,temp_m3_18_8_i,temp_m3_22_4_r,temp_m3_22_4_i,temp_m3_22_8_r,temp_m3_22_8_i,`W12_real,`W12_imag,`W4_real,`W4_imag,`W16_real,`W16_imag);
butterfly butterfly648 (clk,temp_m3_18_4_r,temp_m3_18_4_i,temp_m3_18_8_r,temp_m3_18_8_i,temp_m3_22_4_r,temp_m3_22_4_i,temp_m3_22_8_r,temp_m3_22_8_i,temp_b3_18_4_r,temp_b3_18_4_i,temp_b3_18_8_r,temp_b3_18_8_i,temp_b3_22_4_r,temp_b3_22_4_i,temp_b3_22_8_r,temp_b3_22_8_i);
MULT MULT649 (clk,temp_b2_19_1_r,temp_b2_19_1_i,temp_b2_19_5_r,temp_b2_19_5_i,temp_b2_23_1_r,temp_b2_23_1_i,temp_b2_23_5_r,temp_b2_23_5_i,temp_m3_19_1_r,temp_m3_19_1_i,temp_m3_19_5_r,temp_m3_19_5_i,temp_m3_23_1_r,temp_m3_23_1_i,temp_m3_23_5_r,temp_m3_23_5_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly649 (clk,temp_m3_19_1_r,temp_m3_19_1_i,temp_m3_19_5_r,temp_m3_19_5_i,temp_m3_23_1_r,temp_m3_23_1_i,temp_m3_23_5_r,temp_m3_23_5_i,temp_b3_19_1_r,temp_b3_19_1_i,temp_b3_19_5_r,temp_b3_19_5_i,temp_b3_23_1_r,temp_b3_23_1_i,temp_b3_23_5_r,temp_b3_23_5_i);
MULT MULT650 (clk,temp_b2_19_2_r,temp_b2_19_2_i,temp_b2_19_6_r,temp_b2_19_6_i,temp_b2_23_2_r,temp_b2_23_2_i,temp_b2_23_6_r,temp_b2_23_6_i,temp_m3_19_2_r,temp_m3_19_2_i,temp_m3_19_6_r,temp_m3_19_6_i,temp_m3_23_2_r,temp_m3_23_2_i,temp_m3_23_6_r,temp_m3_23_6_i,`W4_real,`W4_imag,`W8_real,`W8_imag,`W12_real,`W12_imag);
butterfly butterfly650 (clk,temp_m3_19_2_r,temp_m3_19_2_i,temp_m3_19_6_r,temp_m3_19_6_i,temp_m3_23_2_r,temp_m3_23_2_i,temp_m3_23_6_r,temp_m3_23_6_i,temp_b3_19_2_r,temp_b3_19_2_i,temp_b3_19_6_r,temp_b3_19_6_i,temp_b3_23_2_r,temp_b3_23_2_i,temp_b3_23_6_r,temp_b3_23_6_i);
MULT MULT651 (clk,temp_b2_19_3_r,temp_b2_19_3_i,temp_b2_19_7_r,temp_b2_19_7_i,temp_b2_23_3_r,temp_b2_23_3_i,temp_b2_23_7_r,temp_b2_23_7_i,temp_m3_19_3_r,temp_m3_19_3_i,temp_m3_19_7_r,temp_m3_19_7_i,temp_m3_23_3_r,temp_m3_23_3_i,temp_m3_23_7_r,temp_m3_23_7_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly651 (clk,temp_m3_19_3_r,temp_m3_19_3_i,temp_m3_19_7_r,temp_m3_19_7_i,temp_m3_23_3_r,temp_m3_23_3_i,temp_m3_23_7_r,temp_m3_23_7_i,temp_b3_19_3_r,temp_b3_19_3_i,temp_b3_19_7_r,temp_b3_19_7_i,temp_b3_23_3_r,temp_b3_23_3_i,temp_b3_23_7_r,temp_b3_23_7_i);
MULT MULT652 (clk,temp_b2_19_4_r,temp_b2_19_4_i,temp_b2_19_8_r,temp_b2_19_8_i,temp_b2_23_4_r,temp_b2_23_4_i,temp_b2_23_8_r,temp_b2_23_8_i,temp_m3_19_4_r,temp_m3_19_4_i,temp_m3_19_8_r,temp_m3_19_8_i,temp_m3_23_4_r,temp_m3_23_4_i,temp_m3_23_8_r,temp_m3_23_8_i,`W12_real,`W12_imag,`W8_real,`W8_imag,`W20_real,`W20_imag);
butterfly butterfly652 (clk,temp_m3_19_4_r,temp_m3_19_4_i,temp_m3_19_8_r,temp_m3_19_8_i,temp_m3_23_4_r,temp_m3_23_4_i,temp_m3_23_8_r,temp_m3_23_8_i,temp_b3_19_4_r,temp_b3_19_4_i,temp_b3_19_8_r,temp_b3_19_8_i,temp_b3_23_4_r,temp_b3_23_4_i,temp_b3_23_8_r,temp_b3_23_8_i);
MULT MULT653 (clk,temp_b2_20_1_r,temp_b2_20_1_i,temp_b2_20_5_r,temp_b2_20_5_i,temp_b2_24_1_r,temp_b2_24_1_i,temp_b2_24_5_r,temp_b2_24_5_i,temp_m3_20_1_r,temp_m3_20_1_i,temp_m3_20_5_r,temp_m3_20_5_i,temp_m3_24_1_r,temp_m3_24_1_i,temp_m3_24_5_r,temp_m3_24_5_i,`W0_real,`W0_imag,`W12_real,`W12_imag,`W12_real,`W12_imag);
butterfly butterfly653 (clk,temp_m3_20_1_r,temp_m3_20_1_i,temp_m3_20_5_r,temp_m3_20_5_i,temp_m3_24_1_r,temp_m3_24_1_i,temp_m3_24_5_r,temp_m3_24_5_i,temp_b3_20_1_r,temp_b3_20_1_i,temp_b3_20_5_r,temp_b3_20_5_i,temp_b3_24_1_r,temp_b3_24_1_i,temp_b3_24_5_r,temp_b3_24_5_i);
MULT MULT654 (clk,temp_b2_20_2_r,temp_b2_20_2_i,temp_b2_20_6_r,temp_b2_20_6_i,temp_b2_24_2_r,temp_b2_24_2_i,temp_b2_24_6_r,temp_b2_24_6_i,temp_m3_20_2_r,temp_m3_20_2_i,temp_m3_20_6_r,temp_m3_20_6_i,temp_m3_24_2_r,temp_m3_24_2_i,temp_m3_24_6_r,temp_m3_24_6_i,`W4_real,`W4_imag,`W12_real,`W12_imag,`W16_real,`W16_imag);
butterfly butterfly654 (clk,temp_m3_20_2_r,temp_m3_20_2_i,temp_m3_20_6_r,temp_m3_20_6_i,temp_m3_24_2_r,temp_m3_24_2_i,temp_m3_24_6_r,temp_m3_24_6_i,temp_b3_20_2_r,temp_b3_20_2_i,temp_b3_20_6_r,temp_b3_20_6_i,temp_b3_24_2_r,temp_b3_24_2_i,temp_b3_24_6_r,temp_b3_24_6_i);
MULT MULT655 (clk,temp_b2_20_3_r,temp_b2_20_3_i,temp_b2_20_7_r,temp_b2_20_7_i,temp_b2_24_3_r,temp_b2_24_3_i,temp_b2_24_7_r,temp_b2_24_7_i,temp_m3_20_3_r,temp_m3_20_3_i,temp_m3_20_7_r,temp_m3_20_7_i,temp_m3_24_3_r,temp_m3_24_3_i,temp_m3_24_7_r,temp_m3_24_7_i,`W8_real,`W8_imag,`W12_real,`W12_imag,`W20_real,`W20_imag);
butterfly butterfly655 (clk,temp_m3_20_3_r,temp_m3_20_3_i,temp_m3_20_7_r,temp_m3_20_7_i,temp_m3_24_3_r,temp_m3_24_3_i,temp_m3_24_7_r,temp_m3_24_7_i,temp_b3_20_3_r,temp_b3_20_3_i,temp_b3_20_7_r,temp_b3_20_7_i,temp_b3_24_3_r,temp_b3_24_3_i,temp_b3_24_7_r,temp_b3_24_7_i);
MULT MULT656 (clk,temp_b2_20_4_r,temp_b2_20_4_i,temp_b2_20_8_r,temp_b2_20_8_i,temp_b2_24_4_r,temp_b2_24_4_i,temp_b2_24_8_r,temp_b2_24_8_i,temp_m3_20_4_r,temp_m3_20_4_i,temp_m3_20_8_r,temp_m3_20_8_i,temp_m3_24_4_r,temp_m3_24_4_i,temp_m3_24_8_r,temp_m3_24_8_i,`W12_real,`W12_imag,`W12_real,`W12_imag,`W24_real,`W24_imag);
butterfly butterfly656 (clk,temp_m3_20_4_r,temp_m3_20_4_i,temp_m3_20_8_r,temp_m3_20_8_i,temp_m3_24_4_r,temp_m3_24_4_i,temp_m3_24_8_r,temp_m3_24_8_i,temp_b3_20_4_r,temp_b3_20_4_i,temp_b3_20_8_r,temp_b3_20_8_i,temp_b3_24_4_r,temp_b3_24_4_i,temp_b3_24_8_r,temp_b3_24_8_i);
MULT MULT657 (clk,temp_b2_17_9_r,temp_b2_17_9_i,temp_b2_17_13_r,temp_b2_17_13_i,temp_b2_21_9_r,temp_b2_21_9_i,temp_b2_21_13_r,temp_b2_21_13_i,temp_m3_17_9_r,temp_m3_17_9_i,temp_m3_17_13_r,temp_m3_17_13_i,temp_m3_21_9_r,temp_m3_21_9_i,temp_m3_21_13_r,temp_m3_21_13_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly657 (clk,temp_m3_17_9_r,temp_m3_17_9_i,temp_m3_17_13_r,temp_m3_17_13_i,temp_m3_21_9_r,temp_m3_21_9_i,temp_m3_21_13_r,temp_m3_21_13_i,temp_b3_17_9_r,temp_b3_17_9_i,temp_b3_17_13_r,temp_b3_17_13_i,temp_b3_21_9_r,temp_b3_21_9_i,temp_b3_21_13_r,temp_b3_21_13_i);
MULT MULT658 (clk,temp_b2_17_10_r,temp_b2_17_10_i,temp_b2_17_14_r,temp_b2_17_14_i,temp_b2_21_10_r,temp_b2_21_10_i,temp_b2_21_14_r,temp_b2_21_14_i,temp_m3_17_10_r,temp_m3_17_10_i,temp_m3_17_14_r,temp_m3_17_14_i,temp_m3_21_10_r,temp_m3_21_10_i,temp_m3_21_14_r,temp_m3_21_14_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly658 (clk,temp_m3_17_10_r,temp_m3_17_10_i,temp_m3_17_14_r,temp_m3_17_14_i,temp_m3_21_10_r,temp_m3_21_10_i,temp_m3_21_14_r,temp_m3_21_14_i,temp_b3_17_10_r,temp_b3_17_10_i,temp_b3_17_14_r,temp_b3_17_14_i,temp_b3_21_10_r,temp_b3_21_10_i,temp_b3_21_14_r,temp_b3_21_14_i);
MULT MULT659 (clk,temp_b2_17_11_r,temp_b2_17_11_i,temp_b2_17_15_r,temp_b2_17_15_i,temp_b2_21_11_r,temp_b2_21_11_i,temp_b2_21_15_r,temp_b2_21_15_i,temp_m3_17_11_r,temp_m3_17_11_i,temp_m3_17_15_r,temp_m3_17_15_i,temp_m3_21_11_r,temp_m3_21_11_i,temp_m3_21_15_r,temp_m3_21_15_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly659 (clk,temp_m3_17_11_r,temp_m3_17_11_i,temp_m3_17_15_r,temp_m3_17_15_i,temp_m3_21_11_r,temp_m3_21_11_i,temp_m3_21_15_r,temp_m3_21_15_i,temp_b3_17_11_r,temp_b3_17_11_i,temp_b3_17_15_r,temp_b3_17_15_i,temp_b3_21_11_r,temp_b3_21_11_i,temp_b3_21_15_r,temp_b3_21_15_i);
MULT MULT660 (clk,temp_b2_17_12_r,temp_b2_17_12_i,temp_b2_17_16_r,temp_b2_17_16_i,temp_b2_21_12_r,temp_b2_21_12_i,temp_b2_21_16_r,temp_b2_21_16_i,temp_m3_17_12_r,temp_m3_17_12_i,temp_m3_17_16_r,temp_m3_17_16_i,temp_m3_21_12_r,temp_m3_21_12_i,temp_m3_21_16_r,temp_m3_21_16_i,`W12_real,`W12_imag,`W0_real,`W0_imag,`W12_real,`W12_imag);
butterfly butterfly660 (clk,temp_m3_17_12_r,temp_m3_17_12_i,temp_m3_17_16_r,temp_m3_17_16_i,temp_m3_21_12_r,temp_m3_21_12_i,temp_m3_21_16_r,temp_m3_21_16_i,temp_b3_17_12_r,temp_b3_17_12_i,temp_b3_17_16_r,temp_b3_17_16_i,temp_b3_21_12_r,temp_b3_21_12_i,temp_b3_21_16_r,temp_b3_21_16_i);
MULT MULT661 (clk,temp_b2_18_9_r,temp_b2_18_9_i,temp_b2_18_13_r,temp_b2_18_13_i,temp_b2_22_9_r,temp_b2_22_9_i,temp_b2_22_13_r,temp_b2_22_13_i,temp_m3_18_9_r,temp_m3_18_9_i,temp_m3_18_13_r,temp_m3_18_13_i,temp_m3_22_9_r,temp_m3_22_9_i,temp_m3_22_13_r,temp_m3_22_13_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly661 (clk,temp_m3_18_9_r,temp_m3_18_9_i,temp_m3_18_13_r,temp_m3_18_13_i,temp_m3_22_9_r,temp_m3_22_9_i,temp_m3_22_13_r,temp_m3_22_13_i,temp_b3_18_9_r,temp_b3_18_9_i,temp_b3_18_13_r,temp_b3_18_13_i,temp_b3_22_9_r,temp_b3_22_9_i,temp_b3_22_13_r,temp_b3_22_13_i);
MULT MULT662 (clk,temp_b2_18_10_r,temp_b2_18_10_i,temp_b2_18_14_r,temp_b2_18_14_i,temp_b2_22_10_r,temp_b2_22_10_i,temp_b2_22_14_r,temp_b2_22_14_i,temp_m3_18_10_r,temp_m3_18_10_i,temp_m3_18_14_r,temp_m3_18_14_i,temp_m3_22_10_r,temp_m3_22_10_i,temp_m3_22_14_r,temp_m3_22_14_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly662 (clk,temp_m3_18_10_r,temp_m3_18_10_i,temp_m3_18_14_r,temp_m3_18_14_i,temp_m3_22_10_r,temp_m3_22_10_i,temp_m3_22_14_r,temp_m3_22_14_i,temp_b3_18_10_r,temp_b3_18_10_i,temp_b3_18_14_r,temp_b3_18_14_i,temp_b3_22_10_r,temp_b3_22_10_i,temp_b3_22_14_r,temp_b3_22_14_i);
MULT MULT663 (clk,temp_b2_18_11_r,temp_b2_18_11_i,temp_b2_18_15_r,temp_b2_18_15_i,temp_b2_22_11_r,temp_b2_22_11_i,temp_b2_22_15_r,temp_b2_22_15_i,temp_m3_18_11_r,temp_m3_18_11_i,temp_m3_18_15_r,temp_m3_18_15_i,temp_m3_22_11_r,temp_m3_22_11_i,temp_m3_22_15_r,temp_m3_22_15_i,`W8_real,`W8_imag,`W4_real,`W4_imag,`W12_real,`W12_imag);
butterfly butterfly663 (clk,temp_m3_18_11_r,temp_m3_18_11_i,temp_m3_18_15_r,temp_m3_18_15_i,temp_m3_22_11_r,temp_m3_22_11_i,temp_m3_22_15_r,temp_m3_22_15_i,temp_b3_18_11_r,temp_b3_18_11_i,temp_b3_18_15_r,temp_b3_18_15_i,temp_b3_22_11_r,temp_b3_22_11_i,temp_b3_22_15_r,temp_b3_22_15_i);
MULT MULT664 (clk,temp_b2_18_12_r,temp_b2_18_12_i,temp_b2_18_16_r,temp_b2_18_16_i,temp_b2_22_12_r,temp_b2_22_12_i,temp_b2_22_16_r,temp_b2_22_16_i,temp_m3_18_12_r,temp_m3_18_12_i,temp_m3_18_16_r,temp_m3_18_16_i,temp_m3_22_12_r,temp_m3_22_12_i,temp_m3_22_16_r,temp_m3_22_16_i,`W12_real,`W12_imag,`W4_real,`W4_imag,`W16_real,`W16_imag);
butterfly butterfly664 (clk,temp_m3_18_12_r,temp_m3_18_12_i,temp_m3_18_16_r,temp_m3_18_16_i,temp_m3_22_12_r,temp_m3_22_12_i,temp_m3_22_16_r,temp_m3_22_16_i,temp_b3_18_12_r,temp_b3_18_12_i,temp_b3_18_16_r,temp_b3_18_16_i,temp_b3_22_12_r,temp_b3_22_12_i,temp_b3_22_16_r,temp_b3_22_16_i);
MULT MULT665 (clk,temp_b2_19_9_r,temp_b2_19_9_i,temp_b2_19_13_r,temp_b2_19_13_i,temp_b2_23_9_r,temp_b2_23_9_i,temp_b2_23_13_r,temp_b2_23_13_i,temp_m3_19_9_r,temp_m3_19_9_i,temp_m3_19_13_r,temp_m3_19_13_i,temp_m3_23_9_r,temp_m3_23_9_i,temp_m3_23_13_r,temp_m3_23_13_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly665 (clk,temp_m3_19_9_r,temp_m3_19_9_i,temp_m3_19_13_r,temp_m3_19_13_i,temp_m3_23_9_r,temp_m3_23_9_i,temp_m3_23_13_r,temp_m3_23_13_i,temp_b3_19_9_r,temp_b3_19_9_i,temp_b3_19_13_r,temp_b3_19_13_i,temp_b3_23_9_r,temp_b3_23_9_i,temp_b3_23_13_r,temp_b3_23_13_i);
MULT MULT666 (clk,temp_b2_19_10_r,temp_b2_19_10_i,temp_b2_19_14_r,temp_b2_19_14_i,temp_b2_23_10_r,temp_b2_23_10_i,temp_b2_23_14_r,temp_b2_23_14_i,temp_m3_19_10_r,temp_m3_19_10_i,temp_m3_19_14_r,temp_m3_19_14_i,temp_m3_23_10_r,temp_m3_23_10_i,temp_m3_23_14_r,temp_m3_23_14_i,`W4_real,`W4_imag,`W8_real,`W8_imag,`W12_real,`W12_imag);
butterfly butterfly666 (clk,temp_m3_19_10_r,temp_m3_19_10_i,temp_m3_19_14_r,temp_m3_19_14_i,temp_m3_23_10_r,temp_m3_23_10_i,temp_m3_23_14_r,temp_m3_23_14_i,temp_b3_19_10_r,temp_b3_19_10_i,temp_b3_19_14_r,temp_b3_19_14_i,temp_b3_23_10_r,temp_b3_23_10_i,temp_b3_23_14_r,temp_b3_23_14_i);
MULT MULT667 (clk,temp_b2_19_11_r,temp_b2_19_11_i,temp_b2_19_15_r,temp_b2_19_15_i,temp_b2_23_11_r,temp_b2_23_11_i,temp_b2_23_15_r,temp_b2_23_15_i,temp_m3_19_11_r,temp_m3_19_11_i,temp_m3_19_15_r,temp_m3_19_15_i,temp_m3_23_11_r,temp_m3_23_11_i,temp_m3_23_15_r,temp_m3_23_15_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly667 (clk,temp_m3_19_11_r,temp_m3_19_11_i,temp_m3_19_15_r,temp_m3_19_15_i,temp_m3_23_11_r,temp_m3_23_11_i,temp_m3_23_15_r,temp_m3_23_15_i,temp_b3_19_11_r,temp_b3_19_11_i,temp_b3_19_15_r,temp_b3_19_15_i,temp_b3_23_11_r,temp_b3_23_11_i,temp_b3_23_15_r,temp_b3_23_15_i);
MULT MULT668 (clk,temp_b2_19_12_r,temp_b2_19_12_i,temp_b2_19_16_r,temp_b2_19_16_i,temp_b2_23_12_r,temp_b2_23_12_i,temp_b2_23_16_r,temp_b2_23_16_i,temp_m3_19_12_r,temp_m3_19_12_i,temp_m3_19_16_r,temp_m3_19_16_i,temp_m3_23_12_r,temp_m3_23_12_i,temp_m3_23_16_r,temp_m3_23_16_i,`W12_real,`W12_imag,`W8_real,`W8_imag,`W20_real,`W20_imag);
butterfly butterfly668 (clk,temp_m3_19_12_r,temp_m3_19_12_i,temp_m3_19_16_r,temp_m3_19_16_i,temp_m3_23_12_r,temp_m3_23_12_i,temp_m3_23_16_r,temp_m3_23_16_i,temp_b3_19_12_r,temp_b3_19_12_i,temp_b3_19_16_r,temp_b3_19_16_i,temp_b3_23_12_r,temp_b3_23_12_i,temp_b3_23_16_r,temp_b3_23_16_i);
MULT MULT669 (clk,temp_b2_20_9_r,temp_b2_20_9_i,temp_b2_20_13_r,temp_b2_20_13_i,temp_b2_24_9_r,temp_b2_24_9_i,temp_b2_24_13_r,temp_b2_24_13_i,temp_m3_20_9_r,temp_m3_20_9_i,temp_m3_20_13_r,temp_m3_20_13_i,temp_m3_24_9_r,temp_m3_24_9_i,temp_m3_24_13_r,temp_m3_24_13_i,`W0_real,`W0_imag,`W12_real,`W12_imag,`W12_real,`W12_imag);
butterfly butterfly669 (clk,temp_m3_20_9_r,temp_m3_20_9_i,temp_m3_20_13_r,temp_m3_20_13_i,temp_m3_24_9_r,temp_m3_24_9_i,temp_m3_24_13_r,temp_m3_24_13_i,temp_b3_20_9_r,temp_b3_20_9_i,temp_b3_20_13_r,temp_b3_20_13_i,temp_b3_24_9_r,temp_b3_24_9_i,temp_b3_24_13_r,temp_b3_24_13_i);
MULT MULT670 (clk,temp_b2_20_10_r,temp_b2_20_10_i,temp_b2_20_14_r,temp_b2_20_14_i,temp_b2_24_10_r,temp_b2_24_10_i,temp_b2_24_14_r,temp_b2_24_14_i,temp_m3_20_10_r,temp_m3_20_10_i,temp_m3_20_14_r,temp_m3_20_14_i,temp_m3_24_10_r,temp_m3_24_10_i,temp_m3_24_14_r,temp_m3_24_14_i,`W4_real,`W4_imag,`W12_real,`W12_imag,`W16_real,`W16_imag);
butterfly butterfly670 (clk,temp_m3_20_10_r,temp_m3_20_10_i,temp_m3_20_14_r,temp_m3_20_14_i,temp_m3_24_10_r,temp_m3_24_10_i,temp_m3_24_14_r,temp_m3_24_14_i,temp_b3_20_10_r,temp_b3_20_10_i,temp_b3_20_14_r,temp_b3_20_14_i,temp_b3_24_10_r,temp_b3_24_10_i,temp_b3_24_14_r,temp_b3_24_14_i);
MULT MULT671 (clk,temp_b2_20_11_r,temp_b2_20_11_i,temp_b2_20_15_r,temp_b2_20_15_i,temp_b2_24_11_r,temp_b2_24_11_i,temp_b2_24_15_r,temp_b2_24_15_i,temp_m3_20_11_r,temp_m3_20_11_i,temp_m3_20_15_r,temp_m3_20_15_i,temp_m3_24_11_r,temp_m3_24_11_i,temp_m3_24_15_r,temp_m3_24_15_i,`W8_real,`W8_imag,`W12_real,`W12_imag,`W20_real,`W20_imag);
butterfly butterfly671 (clk,temp_m3_20_11_r,temp_m3_20_11_i,temp_m3_20_15_r,temp_m3_20_15_i,temp_m3_24_11_r,temp_m3_24_11_i,temp_m3_24_15_r,temp_m3_24_15_i,temp_b3_20_11_r,temp_b3_20_11_i,temp_b3_20_15_r,temp_b3_20_15_i,temp_b3_24_11_r,temp_b3_24_11_i,temp_b3_24_15_r,temp_b3_24_15_i);
MULT MULT672 (clk,temp_b2_20_12_r,temp_b2_20_12_i,temp_b2_20_16_r,temp_b2_20_16_i,temp_b2_24_12_r,temp_b2_24_12_i,temp_b2_24_16_r,temp_b2_24_16_i,temp_m3_20_12_r,temp_m3_20_12_i,temp_m3_20_16_r,temp_m3_20_16_i,temp_m3_24_12_r,temp_m3_24_12_i,temp_m3_24_16_r,temp_m3_24_16_i,`W12_real,`W12_imag,`W12_real,`W12_imag,`W24_real,`W24_imag);
butterfly butterfly672 (clk,temp_m3_20_12_r,temp_m3_20_12_i,temp_m3_20_16_r,temp_m3_20_16_i,temp_m3_24_12_r,temp_m3_24_12_i,temp_m3_24_16_r,temp_m3_24_16_i,temp_b3_20_12_r,temp_b3_20_12_i,temp_b3_20_16_r,temp_b3_20_16_i,temp_b3_24_12_r,temp_b3_24_12_i,temp_b3_24_16_r,temp_b3_24_16_i);
MULT MULT673 (clk,temp_b2_17_17_r,temp_b2_17_17_i,temp_b2_17_21_r,temp_b2_17_21_i,temp_b2_21_17_r,temp_b2_21_17_i,temp_b2_21_21_r,temp_b2_21_21_i,temp_m3_17_17_r,temp_m3_17_17_i,temp_m3_17_21_r,temp_m3_17_21_i,temp_m3_21_17_r,temp_m3_21_17_i,temp_m3_21_21_r,temp_m3_21_21_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly673 (clk,temp_m3_17_17_r,temp_m3_17_17_i,temp_m3_17_21_r,temp_m3_17_21_i,temp_m3_21_17_r,temp_m3_21_17_i,temp_m3_21_21_r,temp_m3_21_21_i,temp_b3_17_17_r,temp_b3_17_17_i,temp_b3_17_21_r,temp_b3_17_21_i,temp_b3_21_17_r,temp_b3_21_17_i,temp_b3_21_21_r,temp_b3_21_21_i);
MULT MULT674 (clk,temp_b2_17_18_r,temp_b2_17_18_i,temp_b2_17_22_r,temp_b2_17_22_i,temp_b2_21_18_r,temp_b2_21_18_i,temp_b2_21_22_r,temp_b2_21_22_i,temp_m3_17_18_r,temp_m3_17_18_i,temp_m3_17_22_r,temp_m3_17_22_i,temp_m3_21_18_r,temp_m3_21_18_i,temp_m3_21_22_r,temp_m3_21_22_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly674 (clk,temp_m3_17_18_r,temp_m3_17_18_i,temp_m3_17_22_r,temp_m3_17_22_i,temp_m3_21_18_r,temp_m3_21_18_i,temp_m3_21_22_r,temp_m3_21_22_i,temp_b3_17_18_r,temp_b3_17_18_i,temp_b3_17_22_r,temp_b3_17_22_i,temp_b3_21_18_r,temp_b3_21_18_i,temp_b3_21_22_r,temp_b3_21_22_i);
MULT MULT675 (clk,temp_b2_17_19_r,temp_b2_17_19_i,temp_b2_17_23_r,temp_b2_17_23_i,temp_b2_21_19_r,temp_b2_21_19_i,temp_b2_21_23_r,temp_b2_21_23_i,temp_m3_17_19_r,temp_m3_17_19_i,temp_m3_17_23_r,temp_m3_17_23_i,temp_m3_21_19_r,temp_m3_21_19_i,temp_m3_21_23_r,temp_m3_21_23_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly675 (clk,temp_m3_17_19_r,temp_m3_17_19_i,temp_m3_17_23_r,temp_m3_17_23_i,temp_m3_21_19_r,temp_m3_21_19_i,temp_m3_21_23_r,temp_m3_21_23_i,temp_b3_17_19_r,temp_b3_17_19_i,temp_b3_17_23_r,temp_b3_17_23_i,temp_b3_21_19_r,temp_b3_21_19_i,temp_b3_21_23_r,temp_b3_21_23_i);
MULT MULT676 (clk,temp_b2_17_20_r,temp_b2_17_20_i,temp_b2_17_24_r,temp_b2_17_24_i,temp_b2_21_20_r,temp_b2_21_20_i,temp_b2_21_24_r,temp_b2_21_24_i,temp_m3_17_20_r,temp_m3_17_20_i,temp_m3_17_24_r,temp_m3_17_24_i,temp_m3_21_20_r,temp_m3_21_20_i,temp_m3_21_24_r,temp_m3_21_24_i,`W12_real,`W12_imag,`W0_real,`W0_imag,`W12_real,`W12_imag);
butterfly butterfly676 (clk,temp_m3_17_20_r,temp_m3_17_20_i,temp_m3_17_24_r,temp_m3_17_24_i,temp_m3_21_20_r,temp_m3_21_20_i,temp_m3_21_24_r,temp_m3_21_24_i,temp_b3_17_20_r,temp_b3_17_20_i,temp_b3_17_24_r,temp_b3_17_24_i,temp_b3_21_20_r,temp_b3_21_20_i,temp_b3_21_24_r,temp_b3_21_24_i);
MULT MULT677 (clk,temp_b2_18_17_r,temp_b2_18_17_i,temp_b2_18_21_r,temp_b2_18_21_i,temp_b2_22_17_r,temp_b2_22_17_i,temp_b2_22_21_r,temp_b2_22_21_i,temp_m3_18_17_r,temp_m3_18_17_i,temp_m3_18_21_r,temp_m3_18_21_i,temp_m3_22_17_r,temp_m3_22_17_i,temp_m3_22_21_r,temp_m3_22_21_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly677 (clk,temp_m3_18_17_r,temp_m3_18_17_i,temp_m3_18_21_r,temp_m3_18_21_i,temp_m3_22_17_r,temp_m3_22_17_i,temp_m3_22_21_r,temp_m3_22_21_i,temp_b3_18_17_r,temp_b3_18_17_i,temp_b3_18_21_r,temp_b3_18_21_i,temp_b3_22_17_r,temp_b3_22_17_i,temp_b3_22_21_r,temp_b3_22_21_i);
MULT MULT678 (clk,temp_b2_18_18_r,temp_b2_18_18_i,temp_b2_18_22_r,temp_b2_18_22_i,temp_b2_22_18_r,temp_b2_22_18_i,temp_b2_22_22_r,temp_b2_22_22_i,temp_m3_18_18_r,temp_m3_18_18_i,temp_m3_18_22_r,temp_m3_18_22_i,temp_m3_22_18_r,temp_m3_22_18_i,temp_m3_22_22_r,temp_m3_22_22_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly678 (clk,temp_m3_18_18_r,temp_m3_18_18_i,temp_m3_18_22_r,temp_m3_18_22_i,temp_m3_22_18_r,temp_m3_22_18_i,temp_m3_22_22_r,temp_m3_22_22_i,temp_b3_18_18_r,temp_b3_18_18_i,temp_b3_18_22_r,temp_b3_18_22_i,temp_b3_22_18_r,temp_b3_22_18_i,temp_b3_22_22_r,temp_b3_22_22_i);
MULT MULT679 (clk,temp_b2_18_19_r,temp_b2_18_19_i,temp_b2_18_23_r,temp_b2_18_23_i,temp_b2_22_19_r,temp_b2_22_19_i,temp_b2_22_23_r,temp_b2_22_23_i,temp_m3_18_19_r,temp_m3_18_19_i,temp_m3_18_23_r,temp_m3_18_23_i,temp_m3_22_19_r,temp_m3_22_19_i,temp_m3_22_23_r,temp_m3_22_23_i,`W8_real,`W8_imag,`W4_real,`W4_imag,`W12_real,`W12_imag);
butterfly butterfly679 (clk,temp_m3_18_19_r,temp_m3_18_19_i,temp_m3_18_23_r,temp_m3_18_23_i,temp_m3_22_19_r,temp_m3_22_19_i,temp_m3_22_23_r,temp_m3_22_23_i,temp_b3_18_19_r,temp_b3_18_19_i,temp_b3_18_23_r,temp_b3_18_23_i,temp_b3_22_19_r,temp_b3_22_19_i,temp_b3_22_23_r,temp_b3_22_23_i);
MULT MULT680 (clk,temp_b2_18_20_r,temp_b2_18_20_i,temp_b2_18_24_r,temp_b2_18_24_i,temp_b2_22_20_r,temp_b2_22_20_i,temp_b2_22_24_r,temp_b2_22_24_i,temp_m3_18_20_r,temp_m3_18_20_i,temp_m3_18_24_r,temp_m3_18_24_i,temp_m3_22_20_r,temp_m3_22_20_i,temp_m3_22_24_r,temp_m3_22_24_i,`W12_real,`W12_imag,`W4_real,`W4_imag,`W16_real,`W16_imag);
butterfly butterfly680 (clk,temp_m3_18_20_r,temp_m3_18_20_i,temp_m3_18_24_r,temp_m3_18_24_i,temp_m3_22_20_r,temp_m3_22_20_i,temp_m3_22_24_r,temp_m3_22_24_i,temp_b3_18_20_r,temp_b3_18_20_i,temp_b3_18_24_r,temp_b3_18_24_i,temp_b3_22_20_r,temp_b3_22_20_i,temp_b3_22_24_r,temp_b3_22_24_i);
MULT MULT681 (clk,temp_b2_19_17_r,temp_b2_19_17_i,temp_b2_19_21_r,temp_b2_19_21_i,temp_b2_23_17_r,temp_b2_23_17_i,temp_b2_23_21_r,temp_b2_23_21_i,temp_m3_19_17_r,temp_m3_19_17_i,temp_m3_19_21_r,temp_m3_19_21_i,temp_m3_23_17_r,temp_m3_23_17_i,temp_m3_23_21_r,temp_m3_23_21_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly681 (clk,temp_m3_19_17_r,temp_m3_19_17_i,temp_m3_19_21_r,temp_m3_19_21_i,temp_m3_23_17_r,temp_m3_23_17_i,temp_m3_23_21_r,temp_m3_23_21_i,temp_b3_19_17_r,temp_b3_19_17_i,temp_b3_19_21_r,temp_b3_19_21_i,temp_b3_23_17_r,temp_b3_23_17_i,temp_b3_23_21_r,temp_b3_23_21_i);
MULT MULT682 (clk,temp_b2_19_18_r,temp_b2_19_18_i,temp_b2_19_22_r,temp_b2_19_22_i,temp_b2_23_18_r,temp_b2_23_18_i,temp_b2_23_22_r,temp_b2_23_22_i,temp_m3_19_18_r,temp_m3_19_18_i,temp_m3_19_22_r,temp_m3_19_22_i,temp_m3_23_18_r,temp_m3_23_18_i,temp_m3_23_22_r,temp_m3_23_22_i,`W4_real,`W4_imag,`W8_real,`W8_imag,`W12_real,`W12_imag);
butterfly butterfly682 (clk,temp_m3_19_18_r,temp_m3_19_18_i,temp_m3_19_22_r,temp_m3_19_22_i,temp_m3_23_18_r,temp_m3_23_18_i,temp_m3_23_22_r,temp_m3_23_22_i,temp_b3_19_18_r,temp_b3_19_18_i,temp_b3_19_22_r,temp_b3_19_22_i,temp_b3_23_18_r,temp_b3_23_18_i,temp_b3_23_22_r,temp_b3_23_22_i);
MULT MULT683 (clk,temp_b2_19_19_r,temp_b2_19_19_i,temp_b2_19_23_r,temp_b2_19_23_i,temp_b2_23_19_r,temp_b2_23_19_i,temp_b2_23_23_r,temp_b2_23_23_i,temp_m3_19_19_r,temp_m3_19_19_i,temp_m3_19_23_r,temp_m3_19_23_i,temp_m3_23_19_r,temp_m3_23_19_i,temp_m3_23_23_r,temp_m3_23_23_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly683 (clk,temp_m3_19_19_r,temp_m3_19_19_i,temp_m3_19_23_r,temp_m3_19_23_i,temp_m3_23_19_r,temp_m3_23_19_i,temp_m3_23_23_r,temp_m3_23_23_i,temp_b3_19_19_r,temp_b3_19_19_i,temp_b3_19_23_r,temp_b3_19_23_i,temp_b3_23_19_r,temp_b3_23_19_i,temp_b3_23_23_r,temp_b3_23_23_i);
MULT MULT684 (clk,temp_b2_19_20_r,temp_b2_19_20_i,temp_b2_19_24_r,temp_b2_19_24_i,temp_b2_23_20_r,temp_b2_23_20_i,temp_b2_23_24_r,temp_b2_23_24_i,temp_m3_19_20_r,temp_m3_19_20_i,temp_m3_19_24_r,temp_m3_19_24_i,temp_m3_23_20_r,temp_m3_23_20_i,temp_m3_23_24_r,temp_m3_23_24_i,`W12_real,`W12_imag,`W8_real,`W8_imag,`W20_real,`W20_imag);
butterfly butterfly684 (clk,temp_m3_19_20_r,temp_m3_19_20_i,temp_m3_19_24_r,temp_m3_19_24_i,temp_m3_23_20_r,temp_m3_23_20_i,temp_m3_23_24_r,temp_m3_23_24_i,temp_b3_19_20_r,temp_b3_19_20_i,temp_b3_19_24_r,temp_b3_19_24_i,temp_b3_23_20_r,temp_b3_23_20_i,temp_b3_23_24_r,temp_b3_23_24_i);
MULT MULT685 (clk,temp_b2_20_17_r,temp_b2_20_17_i,temp_b2_20_21_r,temp_b2_20_21_i,temp_b2_24_17_r,temp_b2_24_17_i,temp_b2_24_21_r,temp_b2_24_21_i,temp_m3_20_17_r,temp_m3_20_17_i,temp_m3_20_21_r,temp_m3_20_21_i,temp_m3_24_17_r,temp_m3_24_17_i,temp_m3_24_21_r,temp_m3_24_21_i,`W0_real,`W0_imag,`W12_real,`W12_imag,`W12_real,`W12_imag);
butterfly butterfly685 (clk,temp_m3_20_17_r,temp_m3_20_17_i,temp_m3_20_21_r,temp_m3_20_21_i,temp_m3_24_17_r,temp_m3_24_17_i,temp_m3_24_21_r,temp_m3_24_21_i,temp_b3_20_17_r,temp_b3_20_17_i,temp_b3_20_21_r,temp_b3_20_21_i,temp_b3_24_17_r,temp_b3_24_17_i,temp_b3_24_21_r,temp_b3_24_21_i);
MULT MULT686 (clk,temp_b2_20_18_r,temp_b2_20_18_i,temp_b2_20_22_r,temp_b2_20_22_i,temp_b2_24_18_r,temp_b2_24_18_i,temp_b2_24_22_r,temp_b2_24_22_i,temp_m3_20_18_r,temp_m3_20_18_i,temp_m3_20_22_r,temp_m3_20_22_i,temp_m3_24_18_r,temp_m3_24_18_i,temp_m3_24_22_r,temp_m3_24_22_i,`W4_real,`W4_imag,`W12_real,`W12_imag,`W16_real,`W16_imag);
butterfly butterfly686 (clk,temp_m3_20_18_r,temp_m3_20_18_i,temp_m3_20_22_r,temp_m3_20_22_i,temp_m3_24_18_r,temp_m3_24_18_i,temp_m3_24_22_r,temp_m3_24_22_i,temp_b3_20_18_r,temp_b3_20_18_i,temp_b3_20_22_r,temp_b3_20_22_i,temp_b3_24_18_r,temp_b3_24_18_i,temp_b3_24_22_r,temp_b3_24_22_i);
MULT MULT687 (clk,temp_b2_20_19_r,temp_b2_20_19_i,temp_b2_20_23_r,temp_b2_20_23_i,temp_b2_24_19_r,temp_b2_24_19_i,temp_b2_24_23_r,temp_b2_24_23_i,temp_m3_20_19_r,temp_m3_20_19_i,temp_m3_20_23_r,temp_m3_20_23_i,temp_m3_24_19_r,temp_m3_24_19_i,temp_m3_24_23_r,temp_m3_24_23_i,`W8_real,`W8_imag,`W12_real,`W12_imag,`W20_real,`W20_imag);
butterfly butterfly687 (clk,temp_m3_20_19_r,temp_m3_20_19_i,temp_m3_20_23_r,temp_m3_20_23_i,temp_m3_24_19_r,temp_m3_24_19_i,temp_m3_24_23_r,temp_m3_24_23_i,temp_b3_20_19_r,temp_b3_20_19_i,temp_b3_20_23_r,temp_b3_20_23_i,temp_b3_24_19_r,temp_b3_24_19_i,temp_b3_24_23_r,temp_b3_24_23_i);
MULT MULT688 (clk,temp_b2_20_20_r,temp_b2_20_20_i,temp_b2_20_24_r,temp_b2_20_24_i,temp_b2_24_20_r,temp_b2_24_20_i,temp_b2_24_24_r,temp_b2_24_24_i,temp_m3_20_20_r,temp_m3_20_20_i,temp_m3_20_24_r,temp_m3_20_24_i,temp_m3_24_20_r,temp_m3_24_20_i,temp_m3_24_24_r,temp_m3_24_24_i,`W12_real,`W12_imag,`W12_real,`W12_imag,`W24_real,`W24_imag);
butterfly butterfly688 (clk,temp_m3_20_20_r,temp_m3_20_20_i,temp_m3_20_24_r,temp_m3_20_24_i,temp_m3_24_20_r,temp_m3_24_20_i,temp_m3_24_24_r,temp_m3_24_24_i,temp_b3_20_20_r,temp_b3_20_20_i,temp_b3_20_24_r,temp_b3_20_24_i,temp_b3_24_20_r,temp_b3_24_20_i,temp_b3_24_24_r,temp_b3_24_24_i);
MULT MULT689 (clk,temp_b2_17_25_r,temp_b2_17_25_i,temp_b2_17_29_r,temp_b2_17_29_i,temp_b2_21_25_r,temp_b2_21_25_i,temp_b2_21_29_r,temp_b2_21_29_i,temp_m3_17_25_r,temp_m3_17_25_i,temp_m3_17_29_r,temp_m3_17_29_i,temp_m3_21_25_r,temp_m3_21_25_i,temp_m3_21_29_r,temp_m3_21_29_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly689 (clk,temp_m3_17_25_r,temp_m3_17_25_i,temp_m3_17_29_r,temp_m3_17_29_i,temp_m3_21_25_r,temp_m3_21_25_i,temp_m3_21_29_r,temp_m3_21_29_i,temp_b3_17_25_r,temp_b3_17_25_i,temp_b3_17_29_r,temp_b3_17_29_i,temp_b3_21_25_r,temp_b3_21_25_i,temp_b3_21_29_r,temp_b3_21_29_i);
MULT MULT690 (clk,temp_b2_17_26_r,temp_b2_17_26_i,temp_b2_17_30_r,temp_b2_17_30_i,temp_b2_21_26_r,temp_b2_21_26_i,temp_b2_21_30_r,temp_b2_21_30_i,temp_m3_17_26_r,temp_m3_17_26_i,temp_m3_17_30_r,temp_m3_17_30_i,temp_m3_21_26_r,temp_m3_21_26_i,temp_m3_21_30_r,temp_m3_21_30_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly690 (clk,temp_m3_17_26_r,temp_m3_17_26_i,temp_m3_17_30_r,temp_m3_17_30_i,temp_m3_21_26_r,temp_m3_21_26_i,temp_m3_21_30_r,temp_m3_21_30_i,temp_b3_17_26_r,temp_b3_17_26_i,temp_b3_17_30_r,temp_b3_17_30_i,temp_b3_21_26_r,temp_b3_21_26_i,temp_b3_21_30_r,temp_b3_21_30_i);
MULT MULT691 (clk,temp_b2_17_27_r,temp_b2_17_27_i,temp_b2_17_31_r,temp_b2_17_31_i,temp_b2_21_27_r,temp_b2_21_27_i,temp_b2_21_31_r,temp_b2_21_31_i,temp_m3_17_27_r,temp_m3_17_27_i,temp_m3_17_31_r,temp_m3_17_31_i,temp_m3_21_27_r,temp_m3_21_27_i,temp_m3_21_31_r,temp_m3_21_31_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly691 (clk,temp_m3_17_27_r,temp_m3_17_27_i,temp_m3_17_31_r,temp_m3_17_31_i,temp_m3_21_27_r,temp_m3_21_27_i,temp_m3_21_31_r,temp_m3_21_31_i,temp_b3_17_27_r,temp_b3_17_27_i,temp_b3_17_31_r,temp_b3_17_31_i,temp_b3_21_27_r,temp_b3_21_27_i,temp_b3_21_31_r,temp_b3_21_31_i);
MULT MULT692 (clk,temp_b2_17_28_r,temp_b2_17_28_i,temp_b2_17_32_r,temp_b2_17_32_i,temp_b2_21_28_r,temp_b2_21_28_i,temp_b2_21_32_r,temp_b2_21_32_i,temp_m3_17_28_r,temp_m3_17_28_i,temp_m3_17_32_r,temp_m3_17_32_i,temp_m3_21_28_r,temp_m3_21_28_i,temp_m3_21_32_r,temp_m3_21_32_i,`W12_real,`W12_imag,`W0_real,`W0_imag,`W12_real,`W12_imag);
butterfly butterfly692 (clk,temp_m3_17_28_r,temp_m3_17_28_i,temp_m3_17_32_r,temp_m3_17_32_i,temp_m3_21_28_r,temp_m3_21_28_i,temp_m3_21_32_r,temp_m3_21_32_i,temp_b3_17_28_r,temp_b3_17_28_i,temp_b3_17_32_r,temp_b3_17_32_i,temp_b3_21_28_r,temp_b3_21_28_i,temp_b3_21_32_r,temp_b3_21_32_i);
MULT MULT693 (clk,temp_b2_18_25_r,temp_b2_18_25_i,temp_b2_18_29_r,temp_b2_18_29_i,temp_b2_22_25_r,temp_b2_22_25_i,temp_b2_22_29_r,temp_b2_22_29_i,temp_m3_18_25_r,temp_m3_18_25_i,temp_m3_18_29_r,temp_m3_18_29_i,temp_m3_22_25_r,temp_m3_22_25_i,temp_m3_22_29_r,temp_m3_22_29_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly693 (clk,temp_m3_18_25_r,temp_m3_18_25_i,temp_m3_18_29_r,temp_m3_18_29_i,temp_m3_22_25_r,temp_m3_22_25_i,temp_m3_22_29_r,temp_m3_22_29_i,temp_b3_18_25_r,temp_b3_18_25_i,temp_b3_18_29_r,temp_b3_18_29_i,temp_b3_22_25_r,temp_b3_22_25_i,temp_b3_22_29_r,temp_b3_22_29_i);
MULT MULT694 (clk,temp_b2_18_26_r,temp_b2_18_26_i,temp_b2_18_30_r,temp_b2_18_30_i,temp_b2_22_26_r,temp_b2_22_26_i,temp_b2_22_30_r,temp_b2_22_30_i,temp_m3_18_26_r,temp_m3_18_26_i,temp_m3_18_30_r,temp_m3_18_30_i,temp_m3_22_26_r,temp_m3_22_26_i,temp_m3_22_30_r,temp_m3_22_30_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly694 (clk,temp_m3_18_26_r,temp_m3_18_26_i,temp_m3_18_30_r,temp_m3_18_30_i,temp_m3_22_26_r,temp_m3_22_26_i,temp_m3_22_30_r,temp_m3_22_30_i,temp_b3_18_26_r,temp_b3_18_26_i,temp_b3_18_30_r,temp_b3_18_30_i,temp_b3_22_26_r,temp_b3_22_26_i,temp_b3_22_30_r,temp_b3_22_30_i);
MULT MULT695 (clk,temp_b2_18_27_r,temp_b2_18_27_i,temp_b2_18_31_r,temp_b2_18_31_i,temp_b2_22_27_r,temp_b2_22_27_i,temp_b2_22_31_r,temp_b2_22_31_i,temp_m3_18_27_r,temp_m3_18_27_i,temp_m3_18_31_r,temp_m3_18_31_i,temp_m3_22_27_r,temp_m3_22_27_i,temp_m3_22_31_r,temp_m3_22_31_i,`W8_real,`W8_imag,`W4_real,`W4_imag,`W12_real,`W12_imag);
butterfly butterfly695 (clk,temp_m3_18_27_r,temp_m3_18_27_i,temp_m3_18_31_r,temp_m3_18_31_i,temp_m3_22_27_r,temp_m3_22_27_i,temp_m3_22_31_r,temp_m3_22_31_i,temp_b3_18_27_r,temp_b3_18_27_i,temp_b3_18_31_r,temp_b3_18_31_i,temp_b3_22_27_r,temp_b3_22_27_i,temp_b3_22_31_r,temp_b3_22_31_i);
MULT MULT696 (clk,temp_b2_18_28_r,temp_b2_18_28_i,temp_b2_18_32_r,temp_b2_18_32_i,temp_b2_22_28_r,temp_b2_22_28_i,temp_b2_22_32_r,temp_b2_22_32_i,temp_m3_18_28_r,temp_m3_18_28_i,temp_m3_18_32_r,temp_m3_18_32_i,temp_m3_22_28_r,temp_m3_22_28_i,temp_m3_22_32_r,temp_m3_22_32_i,`W12_real,`W12_imag,`W4_real,`W4_imag,`W16_real,`W16_imag);
butterfly butterfly696 (clk,temp_m3_18_28_r,temp_m3_18_28_i,temp_m3_18_32_r,temp_m3_18_32_i,temp_m3_22_28_r,temp_m3_22_28_i,temp_m3_22_32_r,temp_m3_22_32_i,temp_b3_18_28_r,temp_b3_18_28_i,temp_b3_18_32_r,temp_b3_18_32_i,temp_b3_22_28_r,temp_b3_22_28_i,temp_b3_22_32_r,temp_b3_22_32_i);
MULT MULT697 (clk,temp_b2_19_25_r,temp_b2_19_25_i,temp_b2_19_29_r,temp_b2_19_29_i,temp_b2_23_25_r,temp_b2_23_25_i,temp_b2_23_29_r,temp_b2_23_29_i,temp_m3_19_25_r,temp_m3_19_25_i,temp_m3_19_29_r,temp_m3_19_29_i,temp_m3_23_25_r,temp_m3_23_25_i,temp_m3_23_29_r,temp_m3_23_29_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly697 (clk,temp_m3_19_25_r,temp_m3_19_25_i,temp_m3_19_29_r,temp_m3_19_29_i,temp_m3_23_25_r,temp_m3_23_25_i,temp_m3_23_29_r,temp_m3_23_29_i,temp_b3_19_25_r,temp_b3_19_25_i,temp_b3_19_29_r,temp_b3_19_29_i,temp_b3_23_25_r,temp_b3_23_25_i,temp_b3_23_29_r,temp_b3_23_29_i);
MULT MULT698 (clk,temp_b2_19_26_r,temp_b2_19_26_i,temp_b2_19_30_r,temp_b2_19_30_i,temp_b2_23_26_r,temp_b2_23_26_i,temp_b2_23_30_r,temp_b2_23_30_i,temp_m3_19_26_r,temp_m3_19_26_i,temp_m3_19_30_r,temp_m3_19_30_i,temp_m3_23_26_r,temp_m3_23_26_i,temp_m3_23_30_r,temp_m3_23_30_i,`W4_real,`W4_imag,`W8_real,`W8_imag,`W12_real,`W12_imag);
butterfly butterfly698 (clk,temp_m3_19_26_r,temp_m3_19_26_i,temp_m3_19_30_r,temp_m3_19_30_i,temp_m3_23_26_r,temp_m3_23_26_i,temp_m3_23_30_r,temp_m3_23_30_i,temp_b3_19_26_r,temp_b3_19_26_i,temp_b3_19_30_r,temp_b3_19_30_i,temp_b3_23_26_r,temp_b3_23_26_i,temp_b3_23_30_r,temp_b3_23_30_i);
MULT MULT699 (clk,temp_b2_19_27_r,temp_b2_19_27_i,temp_b2_19_31_r,temp_b2_19_31_i,temp_b2_23_27_r,temp_b2_23_27_i,temp_b2_23_31_r,temp_b2_23_31_i,temp_m3_19_27_r,temp_m3_19_27_i,temp_m3_19_31_r,temp_m3_19_31_i,temp_m3_23_27_r,temp_m3_23_27_i,temp_m3_23_31_r,temp_m3_23_31_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly699 (clk,temp_m3_19_27_r,temp_m3_19_27_i,temp_m3_19_31_r,temp_m3_19_31_i,temp_m3_23_27_r,temp_m3_23_27_i,temp_m3_23_31_r,temp_m3_23_31_i,temp_b3_19_27_r,temp_b3_19_27_i,temp_b3_19_31_r,temp_b3_19_31_i,temp_b3_23_27_r,temp_b3_23_27_i,temp_b3_23_31_r,temp_b3_23_31_i);
MULT MULT700 (clk,temp_b2_19_28_r,temp_b2_19_28_i,temp_b2_19_32_r,temp_b2_19_32_i,temp_b2_23_28_r,temp_b2_23_28_i,temp_b2_23_32_r,temp_b2_23_32_i,temp_m3_19_28_r,temp_m3_19_28_i,temp_m3_19_32_r,temp_m3_19_32_i,temp_m3_23_28_r,temp_m3_23_28_i,temp_m3_23_32_r,temp_m3_23_32_i,`W12_real,`W12_imag,`W8_real,`W8_imag,`W20_real,`W20_imag);
butterfly butterfly700 (clk,temp_m3_19_28_r,temp_m3_19_28_i,temp_m3_19_32_r,temp_m3_19_32_i,temp_m3_23_28_r,temp_m3_23_28_i,temp_m3_23_32_r,temp_m3_23_32_i,temp_b3_19_28_r,temp_b3_19_28_i,temp_b3_19_32_r,temp_b3_19_32_i,temp_b3_23_28_r,temp_b3_23_28_i,temp_b3_23_32_r,temp_b3_23_32_i);
MULT MULT701 (clk,temp_b2_20_25_r,temp_b2_20_25_i,temp_b2_20_29_r,temp_b2_20_29_i,temp_b2_24_25_r,temp_b2_24_25_i,temp_b2_24_29_r,temp_b2_24_29_i,temp_m3_20_25_r,temp_m3_20_25_i,temp_m3_20_29_r,temp_m3_20_29_i,temp_m3_24_25_r,temp_m3_24_25_i,temp_m3_24_29_r,temp_m3_24_29_i,`W0_real,`W0_imag,`W12_real,`W12_imag,`W12_real,`W12_imag);
butterfly butterfly701 (clk,temp_m3_20_25_r,temp_m3_20_25_i,temp_m3_20_29_r,temp_m3_20_29_i,temp_m3_24_25_r,temp_m3_24_25_i,temp_m3_24_29_r,temp_m3_24_29_i,temp_b3_20_25_r,temp_b3_20_25_i,temp_b3_20_29_r,temp_b3_20_29_i,temp_b3_24_25_r,temp_b3_24_25_i,temp_b3_24_29_r,temp_b3_24_29_i);
MULT MULT702 (clk,temp_b2_20_26_r,temp_b2_20_26_i,temp_b2_20_30_r,temp_b2_20_30_i,temp_b2_24_26_r,temp_b2_24_26_i,temp_b2_24_30_r,temp_b2_24_30_i,temp_m3_20_26_r,temp_m3_20_26_i,temp_m3_20_30_r,temp_m3_20_30_i,temp_m3_24_26_r,temp_m3_24_26_i,temp_m3_24_30_r,temp_m3_24_30_i,`W4_real,`W4_imag,`W12_real,`W12_imag,`W16_real,`W16_imag);
butterfly butterfly702 (clk,temp_m3_20_26_r,temp_m3_20_26_i,temp_m3_20_30_r,temp_m3_20_30_i,temp_m3_24_26_r,temp_m3_24_26_i,temp_m3_24_30_r,temp_m3_24_30_i,temp_b3_20_26_r,temp_b3_20_26_i,temp_b3_20_30_r,temp_b3_20_30_i,temp_b3_24_26_r,temp_b3_24_26_i,temp_b3_24_30_r,temp_b3_24_30_i);
MULT MULT703 (clk,temp_b2_20_27_r,temp_b2_20_27_i,temp_b2_20_31_r,temp_b2_20_31_i,temp_b2_24_27_r,temp_b2_24_27_i,temp_b2_24_31_r,temp_b2_24_31_i,temp_m3_20_27_r,temp_m3_20_27_i,temp_m3_20_31_r,temp_m3_20_31_i,temp_m3_24_27_r,temp_m3_24_27_i,temp_m3_24_31_r,temp_m3_24_31_i,`W8_real,`W8_imag,`W12_real,`W12_imag,`W20_real,`W20_imag);
butterfly butterfly703 (clk,temp_m3_20_27_r,temp_m3_20_27_i,temp_m3_20_31_r,temp_m3_20_31_i,temp_m3_24_27_r,temp_m3_24_27_i,temp_m3_24_31_r,temp_m3_24_31_i,temp_b3_20_27_r,temp_b3_20_27_i,temp_b3_20_31_r,temp_b3_20_31_i,temp_b3_24_27_r,temp_b3_24_27_i,temp_b3_24_31_r,temp_b3_24_31_i);
MULT MULT704 (clk,temp_b2_20_28_r,temp_b2_20_28_i,temp_b2_20_32_r,temp_b2_20_32_i,temp_b2_24_28_r,temp_b2_24_28_i,temp_b2_24_32_r,temp_b2_24_32_i,temp_m3_20_28_r,temp_m3_20_28_i,temp_m3_20_32_r,temp_m3_20_32_i,temp_m3_24_28_r,temp_m3_24_28_i,temp_m3_24_32_r,temp_m3_24_32_i,`W12_real,`W12_imag,`W12_real,`W12_imag,`W24_real,`W24_imag);
butterfly butterfly704 (clk,temp_m3_20_28_r,temp_m3_20_28_i,temp_m3_20_32_r,temp_m3_20_32_i,temp_m3_24_28_r,temp_m3_24_28_i,temp_m3_24_32_r,temp_m3_24_32_i,temp_b3_20_28_r,temp_b3_20_28_i,temp_b3_20_32_r,temp_b3_20_32_i,temp_b3_24_28_r,temp_b3_24_28_i,temp_b3_24_32_r,temp_b3_24_32_i);
MULT MULT705 (clk,temp_b2_25_1_r,temp_b2_25_1_i,temp_b2_25_5_r,temp_b2_25_5_i,temp_b2_29_1_r,temp_b2_29_1_i,temp_b2_29_5_r,temp_b2_29_5_i,temp_m3_25_1_r,temp_m3_25_1_i,temp_m3_25_5_r,temp_m3_25_5_i,temp_m3_29_1_r,temp_m3_29_1_i,temp_m3_29_5_r,temp_m3_29_5_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly705 (clk,temp_m3_25_1_r,temp_m3_25_1_i,temp_m3_25_5_r,temp_m3_25_5_i,temp_m3_29_1_r,temp_m3_29_1_i,temp_m3_29_5_r,temp_m3_29_5_i,temp_b3_25_1_r,temp_b3_25_1_i,temp_b3_25_5_r,temp_b3_25_5_i,temp_b3_29_1_r,temp_b3_29_1_i,temp_b3_29_5_r,temp_b3_29_5_i);
MULT MULT706 (clk,temp_b2_25_2_r,temp_b2_25_2_i,temp_b2_25_6_r,temp_b2_25_6_i,temp_b2_29_2_r,temp_b2_29_2_i,temp_b2_29_6_r,temp_b2_29_6_i,temp_m3_25_2_r,temp_m3_25_2_i,temp_m3_25_6_r,temp_m3_25_6_i,temp_m3_29_2_r,temp_m3_29_2_i,temp_m3_29_6_r,temp_m3_29_6_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly706 (clk,temp_m3_25_2_r,temp_m3_25_2_i,temp_m3_25_6_r,temp_m3_25_6_i,temp_m3_29_2_r,temp_m3_29_2_i,temp_m3_29_6_r,temp_m3_29_6_i,temp_b3_25_2_r,temp_b3_25_2_i,temp_b3_25_6_r,temp_b3_25_6_i,temp_b3_29_2_r,temp_b3_29_2_i,temp_b3_29_6_r,temp_b3_29_6_i);
MULT MULT707 (clk,temp_b2_25_3_r,temp_b2_25_3_i,temp_b2_25_7_r,temp_b2_25_7_i,temp_b2_29_3_r,temp_b2_29_3_i,temp_b2_29_7_r,temp_b2_29_7_i,temp_m3_25_3_r,temp_m3_25_3_i,temp_m3_25_7_r,temp_m3_25_7_i,temp_m3_29_3_r,temp_m3_29_3_i,temp_m3_29_7_r,temp_m3_29_7_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly707 (clk,temp_m3_25_3_r,temp_m3_25_3_i,temp_m3_25_7_r,temp_m3_25_7_i,temp_m3_29_3_r,temp_m3_29_3_i,temp_m3_29_7_r,temp_m3_29_7_i,temp_b3_25_3_r,temp_b3_25_3_i,temp_b3_25_7_r,temp_b3_25_7_i,temp_b3_29_3_r,temp_b3_29_3_i,temp_b3_29_7_r,temp_b3_29_7_i);
MULT MULT708 (clk,temp_b2_25_4_r,temp_b2_25_4_i,temp_b2_25_8_r,temp_b2_25_8_i,temp_b2_29_4_r,temp_b2_29_4_i,temp_b2_29_8_r,temp_b2_29_8_i,temp_m3_25_4_r,temp_m3_25_4_i,temp_m3_25_8_r,temp_m3_25_8_i,temp_m3_29_4_r,temp_m3_29_4_i,temp_m3_29_8_r,temp_m3_29_8_i,`W12_real,`W12_imag,`W0_real,`W0_imag,`W12_real,`W12_imag);
butterfly butterfly708 (clk,temp_m3_25_4_r,temp_m3_25_4_i,temp_m3_25_8_r,temp_m3_25_8_i,temp_m3_29_4_r,temp_m3_29_4_i,temp_m3_29_8_r,temp_m3_29_8_i,temp_b3_25_4_r,temp_b3_25_4_i,temp_b3_25_8_r,temp_b3_25_8_i,temp_b3_29_4_r,temp_b3_29_4_i,temp_b3_29_8_r,temp_b3_29_8_i);
MULT MULT709 (clk,temp_b2_26_1_r,temp_b2_26_1_i,temp_b2_26_5_r,temp_b2_26_5_i,temp_b2_30_1_r,temp_b2_30_1_i,temp_b2_30_5_r,temp_b2_30_5_i,temp_m3_26_1_r,temp_m3_26_1_i,temp_m3_26_5_r,temp_m3_26_5_i,temp_m3_30_1_r,temp_m3_30_1_i,temp_m3_30_5_r,temp_m3_30_5_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly709 (clk,temp_m3_26_1_r,temp_m3_26_1_i,temp_m3_26_5_r,temp_m3_26_5_i,temp_m3_30_1_r,temp_m3_30_1_i,temp_m3_30_5_r,temp_m3_30_5_i,temp_b3_26_1_r,temp_b3_26_1_i,temp_b3_26_5_r,temp_b3_26_5_i,temp_b3_30_1_r,temp_b3_30_1_i,temp_b3_30_5_r,temp_b3_30_5_i);
MULT MULT710 (clk,temp_b2_26_2_r,temp_b2_26_2_i,temp_b2_26_6_r,temp_b2_26_6_i,temp_b2_30_2_r,temp_b2_30_2_i,temp_b2_30_6_r,temp_b2_30_6_i,temp_m3_26_2_r,temp_m3_26_2_i,temp_m3_26_6_r,temp_m3_26_6_i,temp_m3_30_2_r,temp_m3_30_2_i,temp_m3_30_6_r,temp_m3_30_6_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly710 (clk,temp_m3_26_2_r,temp_m3_26_2_i,temp_m3_26_6_r,temp_m3_26_6_i,temp_m3_30_2_r,temp_m3_30_2_i,temp_m3_30_6_r,temp_m3_30_6_i,temp_b3_26_2_r,temp_b3_26_2_i,temp_b3_26_6_r,temp_b3_26_6_i,temp_b3_30_2_r,temp_b3_30_2_i,temp_b3_30_6_r,temp_b3_30_6_i);
MULT MULT711 (clk,temp_b2_26_3_r,temp_b2_26_3_i,temp_b2_26_7_r,temp_b2_26_7_i,temp_b2_30_3_r,temp_b2_30_3_i,temp_b2_30_7_r,temp_b2_30_7_i,temp_m3_26_3_r,temp_m3_26_3_i,temp_m3_26_7_r,temp_m3_26_7_i,temp_m3_30_3_r,temp_m3_30_3_i,temp_m3_30_7_r,temp_m3_30_7_i,`W8_real,`W8_imag,`W4_real,`W4_imag,`W12_real,`W12_imag);
butterfly butterfly711 (clk,temp_m3_26_3_r,temp_m3_26_3_i,temp_m3_26_7_r,temp_m3_26_7_i,temp_m3_30_3_r,temp_m3_30_3_i,temp_m3_30_7_r,temp_m3_30_7_i,temp_b3_26_3_r,temp_b3_26_3_i,temp_b3_26_7_r,temp_b3_26_7_i,temp_b3_30_3_r,temp_b3_30_3_i,temp_b3_30_7_r,temp_b3_30_7_i);
MULT MULT712 (clk,temp_b2_26_4_r,temp_b2_26_4_i,temp_b2_26_8_r,temp_b2_26_8_i,temp_b2_30_4_r,temp_b2_30_4_i,temp_b2_30_8_r,temp_b2_30_8_i,temp_m3_26_4_r,temp_m3_26_4_i,temp_m3_26_8_r,temp_m3_26_8_i,temp_m3_30_4_r,temp_m3_30_4_i,temp_m3_30_8_r,temp_m3_30_8_i,`W12_real,`W12_imag,`W4_real,`W4_imag,`W16_real,`W16_imag);
butterfly butterfly712 (clk,temp_m3_26_4_r,temp_m3_26_4_i,temp_m3_26_8_r,temp_m3_26_8_i,temp_m3_30_4_r,temp_m3_30_4_i,temp_m3_30_8_r,temp_m3_30_8_i,temp_b3_26_4_r,temp_b3_26_4_i,temp_b3_26_8_r,temp_b3_26_8_i,temp_b3_30_4_r,temp_b3_30_4_i,temp_b3_30_8_r,temp_b3_30_8_i);
MULT MULT713 (clk,temp_b2_27_1_r,temp_b2_27_1_i,temp_b2_27_5_r,temp_b2_27_5_i,temp_b2_31_1_r,temp_b2_31_1_i,temp_b2_31_5_r,temp_b2_31_5_i,temp_m3_27_1_r,temp_m3_27_1_i,temp_m3_27_5_r,temp_m3_27_5_i,temp_m3_31_1_r,temp_m3_31_1_i,temp_m3_31_5_r,temp_m3_31_5_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly713 (clk,temp_m3_27_1_r,temp_m3_27_1_i,temp_m3_27_5_r,temp_m3_27_5_i,temp_m3_31_1_r,temp_m3_31_1_i,temp_m3_31_5_r,temp_m3_31_5_i,temp_b3_27_1_r,temp_b3_27_1_i,temp_b3_27_5_r,temp_b3_27_5_i,temp_b3_31_1_r,temp_b3_31_1_i,temp_b3_31_5_r,temp_b3_31_5_i);
MULT MULT714 (clk,temp_b2_27_2_r,temp_b2_27_2_i,temp_b2_27_6_r,temp_b2_27_6_i,temp_b2_31_2_r,temp_b2_31_2_i,temp_b2_31_6_r,temp_b2_31_6_i,temp_m3_27_2_r,temp_m3_27_2_i,temp_m3_27_6_r,temp_m3_27_6_i,temp_m3_31_2_r,temp_m3_31_2_i,temp_m3_31_6_r,temp_m3_31_6_i,`W4_real,`W4_imag,`W8_real,`W8_imag,`W12_real,`W12_imag);
butterfly butterfly714 (clk,temp_m3_27_2_r,temp_m3_27_2_i,temp_m3_27_6_r,temp_m3_27_6_i,temp_m3_31_2_r,temp_m3_31_2_i,temp_m3_31_6_r,temp_m3_31_6_i,temp_b3_27_2_r,temp_b3_27_2_i,temp_b3_27_6_r,temp_b3_27_6_i,temp_b3_31_2_r,temp_b3_31_2_i,temp_b3_31_6_r,temp_b3_31_6_i);
MULT MULT715 (clk,temp_b2_27_3_r,temp_b2_27_3_i,temp_b2_27_7_r,temp_b2_27_7_i,temp_b2_31_3_r,temp_b2_31_3_i,temp_b2_31_7_r,temp_b2_31_7_i,temp_m3_27_3_r,temp_m3_27_3_i,temp_m3_27_7_r,temp_m3_27_7_i,temp_m3_31_3_r,temp_m3_31_3_i,temp_m3_31_7_r,temp_m3_31_7_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly715 (clk,temp_m3_27_3_r,temp_m3_27_3_i,temp_m3_27_7_r,temp_m3_27_7_i,temp_m3_31_3_r,temp_m3_31_3_i,temp_m3_31_7_r,temp_m3_31_7_i,temp_b3_27_3_r,temp_b3_27_3_i,temp_b3_27_7_r,temp_b3_27_7_i,temp_b3_31_3_r,temp_b3_31_3_i,temp_b3_31_7_r,temp_b3_31_7_i);
MULT MULT716 (clk,temp_b2_27_4_r,temp_b2_27_4_i,temp_b2_27_8_r,temp_b2_27_8_i,temp_b2_31_4_r,temp_b2_31_4_i,temp_b2_31_8_r,temp_b2_31_8_i,temp_m3_27_4_r,temp_m3_27_4_i,temp_m3_27_8_r,temp_m3_27_8_i,temp_m3_31_4_r,temp_m3_31_4_i,temp_m3_31_8_r,temp_m3_31_8_i,`W12_real,`W12_imag,`W8_real,`W8_imag,`W20_real,`W20_imag);
butterfly butterfly716 (clk,temp_m3_27_4_r,temp_m3_27_4_i,temp_m3_27_8_r,temp_m3_27_8_i,temp_m3_31_4_r,temp_m3_31_4_i,temp_m3_31_8_r,temp_m3_31_8_i,temp_b3_27_4_r,temp_b3_27_4_i,temp_b3_27_8_r,temp_b3_27_8_i,temp_b3_31_4_r,temp_b3_31_4_i,temp_b3_31_8_r,temp_b3_31_8_i);
MULT MULT717 (clk,temp_b2_28_1_r,temp_b2_28_1_i,temp_b2_28_5_r,temp_b2_28_5_i,temp_b2_32_1_r,temp_b2_32_1_i,temp_b2_32_5_r,temp_b2_32_5_i,temp_m3_28_1_r,temp_m3_28_1_i,temp_m3_28_5_r,temp_m3_28_5_i,temp_m3_32_1_r,temp_m3_32_1_i,temp_m3_32_5_r,temp_m3_32_5_i,`W0_real,`W0_imag,`W12_real,`W12_imag,`W12_real,`W12_imag);
butterfly butterfly717 (clk,temp_m3_28_1_r,temp_m3_28_1_i,temp_m3_28_5_r,temp_m3_28_5_i,temp_m3_32_1_r,temp_m3_32_1_i,temp_m3_32_5_r,temp_m3_32_5_i,temp_b3_28_1_r,temp_b3_28_1_i,temp_b3_28_5_r,temp_b3_28_5_i,temp_b3_32_1_r,temp_b3_32_1_i,temp_b3_32_5_r,temp_b3_32_5_i);
MULT MULT718 (clk,temp_b2_28_2_r,temp_b2_28_2_i,temp_b2_28_6_r,temp_b2_28_6_i,temp_b2_32_2_r,temp_b2_32_2_i,temp_b2_32_6_r,temp_b2_32_6_i,temp_m3_28_2_r,temp_m3_28_2_i,temp_m3_28_6_r,temp_m3_28_6_i,temp_m3_32_2_r,temp_m3_32_2_i,temp_m3_32_6_r,temp_m3_32_6_i,`W4_real,`W4_imag,`W12_real,`W12_imag,`W16_real,`W16_imag);
butterfly butterfly718 (clk,temp_m3_28_2_r,temp_m3_28_2_i,temp_m3_28_6_r,temp_m3_28_6_i,temp_m3_32_2_r,temp_m3_32_2_i,temp_m3_32_6_r,temp_m3_32_6_i,temp_b3_28_2_r,temp_b3_28_2_i,temp_b3_28_6_r,temp_b3_28_6_i,temp_b3_32_2_r,temp_b3_32_2_i,temp_b3_32_6_r,temp_b3_32_6_i);
MULT MULT719 (clk,temp_b2_28_3_r,temp_b2_28_3_i,temp_b2_28_7_r,temp_b2_28_7_i,temp_b2_32_3_r,temp_b2_32_3_i,temp_b2_32_7_r,temp_b2_32_7_i,temp_m3_28_3_r,temp_m3_28_3_i,temp_m3_28_7_r,temp_m3_28_7_i,temp_m3_32_3_r,temp_m3_32_3_i,temp_m3_32_7_r,temp_m3_32_7_i,`W8_real,`W8_imag,`W12_real,`W12_imag,`W20_real,`W20_imag);
butterfly butterfly719 (clk,temp_m3_28_3_r,temp_m3_28_3_i,temp_m3_28_7_r,temp_m3_28_7_i,temp_m3_32_3_r,temp_m3_32_3_i,temp_m3_32_7_r,temp_m3_32_7_i,temp_b3_28_3_r,temp_b3_28_3_i,temp_b3_28_7_r,temp_b3_28_7_i,temp_b3_32_3_r,temp_b3_32_3_i,temp_b3_32_7_r,temp_b3_32_7_i);
MULT MULT720 (clk,temp_b2_28_4_r,temp_b2_28_4_i,temp_b2_28_8_r,temp_b2_28_8_i,temp_b2_32_4_r,temp_b2_32_4_i,temp_b2_32_8_r,temp_b2_32_8_i,temp_m3_28_4_r,temp_m3_28_4_i,temp_m3_28_8_r,temp_m3_28_8_i,temp_m3_32_4_r,temp_m3_32_4_i,temp_m3_32_8_r,temp_m3_32_8_i,`W12_real,`W12_imag,`W12_real,`W12_imag,`W24_real,`W24_imag);
butterfly butterfly720 (clk,temp_m3_28_4_r,temp_m3_28_4_i,temp_m3_28_8_r,temp_m3_28_8_i,temp_m3_32_4_r,temp_m3_32_4_i,temp_m3_32_8_r,temp_m3_32_8_i,temp_b3_28_4_r,temp_b3_28_4_i,temp_b3_28_8_r,temp_b3_28_8_i,temp_b3_32_4_r,temp_b3_32_4_i,temp_b3_32_8_r,temp_b3_32_8_i);
MULT MULT721 (clk,temp_b2_25_9_r,temp_b2_25_9_i,temp_b2_25_13_r,temp_b2_25_13_i,temp_b2_29_9_r,temp_b2_29_9_i,temp_b2_29_13_r,temp_b2_29_13_i,temp_m3_25_9_r,temp_m3_25_9_i,temp_m3_25_13_r,temp_m3_25_13_i,temp_m3_29_9_r,temp_m3_29_9_i,temp_m3_29_13_r,temp_m3_29_13_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly721 (clk,temp_m3_25_9_r,temp_m3_25_9_i,temp_m3_25_13_r,temp_m3_25_13_i,temp_m3_29_9_r,temp_m3_29_9_i,temp_m3_29_13_r,temp_m3_29_13_i,temp_b3_25_9_r,temp_b3_25_9_i,temp_b3_25_13_r,temp_b3_25_13_i,temp_b3_29_9_r,temp_b3_29_9_i,temp_b3_29_13_r,temp_b3_29_13_i);
MULT MULT722 (clk,temp_b2_25_10_r,temp_b2_25_10_i,temp_b2_25_14_r,temp_b2_25_14_i,temp_b2_29_10_r,temp_b2_29_10_i,temp_b2_29_14_r,temp_b2_29_14_i,temp_m3_25_10_r,temp_m3_25_10_i,temp_m3_25_14_r,temp_m3_25_14_i,temp_m3_29_10_r,temp_m3_29_10_i,temp_m3_29_14_r,temp_m3_29_14_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly722 (clk,temp_m3_25_10_r,temp_m3_25_10_i,temp_m3_25_14_r,temp_m3_25_14_i,temp_m3_29_10_r,temp_m3_29_10_i,temp_m3_29_14_r,temp_m3_29_14_i,temp_b3_25_10_r,temp_b3_25_10_i,temp_b3_25_14_r,temp_b3_25_14_i,temp_b3_29_10_r,temp_b3_29_10_i,temp_b3_29_14_r,temp_b3_29_14_i);
MULT MULT723 (clk,temp_b2_25_11_r,temp_b2_25_11_i,temp_b2_25_15_r,temp_b2_25_15_i,temp_b2_29_11_r,temp_b2_29_11_i,temp_b2_29_15_r,temp_b2_29_15_i,temp_m3_25_11_r,temp_m3_25_11_i,temp_m3_25_15_r,temp_m3_25_15_i,temp_m3_29_11_r,temp_m3_29_11_i,temp_m3_29_15_r,temp_m3_29_15_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly723 (clk,temp_m3_25_11_r,temp_m3_25_11_i,temp_m3_25_15_r,temp_m3_25_15_i,temp_m3_29_11_r,temp_m3_29_11_i,temp_m3_29_15_r,temp_m3_29_15_i,temp_b3_25_11_r,temp_b3_25_11_i,temp_b3_25_15_r,temp_b3_25_15_i,temp_b3_29_11_r,temp_b3_29_11_i,temp_b3_29_15_r,temp_b3_29_15_i);
MULT MULT724 (clk,temp_b2_25_12_r,temp_b2_25_12_i,temp_b2_25_16_r,temp_b2_25_16_i,temp_b2_29_12_r,temp_b2_29_12_i,temp_b2_29_16_r,temp_b2_29_16_i,temp_m3_25_12_r,temp_m3_25_12_i,temp_m3_25_16_r,temp_m3_25_16_i,temp_m3_29_12_r,temp_m3_29_12_i,temp_m3_29_16_r,temp_m3_29_16_i,`W12_real,`W12_imag,`W0_real,`W0_imag,`W12_real,`W12_imag);
butterfly butterfly724 (clk,temp_m3_25_12_r,temp_m3_25_12_i,temp_m3_25_16_r,temp_m3_25_16_i,temp_m3_29_12_r,temp_m3_29_12_i,temp_m3_29_16_r,temp_m3_29_16_i,temp_b3_25_12_r,temp_b3_25_12_i,temp_b3_25_16_r,temp_b3_25_16_i,temp_b3_29_12_r,temp_b3_29_12_i,temp_b3_29_16_r,temp_b3_29_16_i);
MULT MULT725 (clk,temp_b2_26_9_r,temp_b2_26_9_i,temp_b2_26_13_r,temp_b2_26_13_i,temp_b2_30_9_r,temp_b2_30_9_i,temp_b2_30_13_r,temp_b2_30_13_i,temp_m3_26_9_r,temp_m3_26_9_i,temp_m3_26_13_r,temp_m3_26_13_i,temp_m3_30_9_r,temp_m3_30_9_i,temp_m3_30_13_r,temp_m3_30_13_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly725 (clk,temp_m3_26_9_r,temp_m3_26_9_i,temp_m3_26_13_r,temp_m3_26_13_i,temp_m3_30_9_r,temp_m3_30_9_i,temp_m3_30_13_r,temp_m3_30_13_i,temp_b3_26_9_r,temp_b3_26_9_i,temp_b3_26_13_r,temp_b3_26_13_i,temp_b3_30_9_r,temp_b3_30_9_i,temp_b3_30_13_r,temp_b3_30_13_i);
MULT MULT726 (clk,temp_b2_26_10_r,temp_b2_26_10_i,temp_b2_26_14_r,temp_b2_26_14_i,temp_b2_30_10_r,temp_b2_30_10_i,temp_b2_30_14_r,temp_b2_30_14_i,temp_m3_26_10_r,temp_m3_26_10_i,temp_m3_26_14_r,temp_m3_26_14_i,temp_m3_30_10_r,temp_m3_30_10_i,temp_m3_30_14_r,temp_m3_30_14_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly726 (clk,temp_m3_26_10_r,temp_m3_26_10_i,temp_m3_26_14_r,temp_m3_26_14_i,temp_m3_30_10_r,temp_m3_30_10_i,temp_m3_30_14_r,temp_m3_30_14_i,temp_b3_26_10_r,temp_b3_26_10_i,temp_b3_26_14_r,temp_b3_26_14_i,temp_b3_30_10_r,temp_b3_30_10_i,temp_b3_30_14_r,temp_b3_30_14_i);
MULT MULT727 (clk,temp_b2_26_11_r,temp_b2_26_11_i,temp_b2_26_15_r,temp_b2_26_15_i,temp_b2_30_11_r,temp_b2_30_11_i,temp_b2_30_15_r,temp_b2_30_15_i,temp_m3_26_11_r,temp_m3_26_11_i,temp_m3_26_15_r,temp_m3_26_15_i,temp_m3_30_11_r,temp_m3_30_11_i,temp_m3_30_15_r,temp_m3_30_15_i,`W8_real,`W8_imag,`W4_real,`W4_imag,`W12_real,`W12_imag);
butterfly butterfly727 (clk,temp_m3_26_11_r,temp_m3_26_11_i,temp_m3_26_15_r,temp_m3_26_15_i,temp_m3_30_11_r,temp_m3_30_11_i,temp_m3_30_15_r,temp_m3_30_15_i,temp_b3_26_11_r,temp_b3_26_11_i,temp_b3_26_15_r,temp_b3_26_15_i,temp_b3_30_11_r,temp_b3_30_11_i,temp_b3_30_15_r,temp_b3_30_15_i);
MULT MULT728 (clk,temp_b2_26_12_r,temp_b2_26_12_i,temp_b2_26_16_r,temp_b2_26_16_i,temp_b2_30_12_r,temp_b2_30_12_i,temp_b2_30_16_r,temp_b2_30_16_i,temp_m3_26_12_r,temp_m3_26_12_i,temp_m3_26_16_r,temp_m3_26_16_i,temp_m3_30_12_r,temp_m3_30_12_i,temp_m3_30_16_r,temp_m3_30_16_i,`W12_real,`W12_imag,`W4_real,`W4_imag,`W16_real,`W16_imag);
butterfly butterfly728 (clk,temp_m3_26_12_r,temp_m3_26_12_i,temp_m3_26_16_r,temp_m3_26_16_i,temp_m3_30_12_r,temp_m3_30_12_i,temp_m3_30_16_r,temp_m3_30_16_i,temp_b3_26_12_r,temp_b3_26_12_i,temp_b3_26_16_r,temp_b3_26_16_i,temp_b3_30_12_r,temp_b3_30_12_i,temp_b3_30_16_r,temp_b3_30_16_i);
MULT MULT729 (clk,temp_b2_27_9_r,temp_b2_27_9_i,temp_b2_27_13_r,temp_b2_27_13_i,temp_b2_31_9_r,temp_b2_31_9_i,temp_b2_31_13_r,temp_b2_31_13_i,temp_m3_27_9_r,temp_m3_27_9_i,temp_m3_27_13_r,temp_m3_27_13_i,temp_m3_31_9_r,temp_m3_31_9_i,temp_m3_31_13_r,temp_m3_31_13_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly729 (clk,temp_m3_27_9_r,temp_m3_27_9_i,temp_m3_27_13_r,temp_m3_27_13_i,temp_m3_31_9_r,temp_m3_31_9_i,temp_m3_31_13_r,temp_m3_31_13_i,temp_b3_27_9_r,temp_b3_27_9_i,temp_b3_27_13_r,temp_b3_27_13_i,temp_b3_31_9_r,temp_b3_31_9_i,temp_b3_31_13_r,temp_b3_31_13_i);
MULT MULT730 (clk,temp_b2_27_10_r,temp_b2_27_10_i,temp_b2_27_14_r,temp_b2_27_14_i,temp_b2_31_10_r,temp_b2_31_10_i,temp_b2_31_14_r,temp_b2_31_14_i,temp_m3_27_10_r,temp_m3_27_10_i,temp_m3_27_14_r,temp_m3_27_14_i,temp_m3_31_10_r,temp_m3_31_10_i,temp_m3_31_14_r,temp_m3_31_14_i,`W4_real,`W4_imag,`W8_real,`W8_imag,`W12_real,`W12_imag);
butterfly butterfly730 (clk,temp_m3_27_10_r,temp_m3_27_10_i,temp_m3_27_14_r,temp_m3_27_14_i,temp_m3_31_10_r,temp_m3_31_10_i,temp_m3_31_14_r,temp_m3_31_14_i,temp_b3_27_10_r,temp_b3_27_10_i,temp_b3_27_14_r,temp_b3_27_14_i,temp_b3_31_10_r,temp_b3_31_10_i,temp_b3_31_14_r,temp_b3_31_14_i);
MULT MULT731 (clk,temp_b2_27_11_r,temp_b2_27_11_i,temp_b2_27_15_r,temp_b2_27_15_i,temp_b2_31_11_r,temp_b2_31_11_i,temp_b2_31_15_r,temp_b2_31_15_i,temp_m3_27_11_r,temp_m3_27_11_i,temp_m3_27_15_r,temp_m3_27_15_i,temp_m3_31_11_r,temp_m3_31_11_i,temp_m3_31_15_r,temp_m3_31_15_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly731 (clk,temp_m3_27_11_r,temp_m3_27_11_i,temp_m3_27_15_r,temp_m3_27_15_i,temp_m3_31_11_r,temp_m3_31_11_i,temp_m3_31_15_r,temp_m3_31_15_i,temp_b3_27_11_r,temp_b3_27_11_i,temp_b3_27_15_r,temp_b3_27_15_i,temp_b3_31_11_r,temp_b3_31_11_i,temp_b3_31_15_r,temp_b3_31_15_i);
MULT MULT732 (clk,temp_b2_27_12_r,temp_b2_27_12_i,temp_b2_27_16_r,temp_b2_27_16_i,temp_b2_31_12_r,temp_b2_31_12_i,temp_b2_31_16_r,temp_b2_31_16_i,temp_m3_27_12_r,temp_m3_27_12_i,temp_m3_27_16_r,temp_m3_27_16_i,temp_m3_31_12_r,temp_m3_31_12_i,temp_m3_31_16_r,temp_m3_31_16_i,`W12_real,`W12_imag,`W8_real,`W8_imag,`W20_real,`W20_imag);
butterfly butterfly732 (clk,temp_m3_27_12_r,temp_m3_27_12_i,temp_m3_27_16_r,temp_m3_27_16_i,temp_m3_31_12_r,temp_m3_31_12_i,temp_m3_31_16_r,temp_m3_31_16_i,temp_b3_27_12_r,temp_b3_27_12_i,temp_b3_27_16_r,temp_b3_27_16_i,temp_b3_31_12_r,temp_b3_31_12_i,temp_b3_31_16_r,temp_b3_31_16_i);
MULT MULT733 (clk,temp_b2_28_9_r,temp_b2_28_9_i,temp_b2_28_13_r,temp_b2_28_13_i,temp_b2_32_9_r,temp_b2_32_9_i,temp_b2_32_13_r,temp_b2_32_13_i,temp_m3_28_9_r,temp_m3_28_9_i,temp_m3_28_13_r,temp_m3_28_13_i,temp_m3_32_9_r,temp_m3_32_9_i,temp_m3_32_13_r,temp_m3_32_13_i,`W0_real,`W0_imag,`W12_real,`W12_imag,`W12_real,`W12_imag);
butterfly butterfly733 (clk,temp_m3_28_9_r,temp_m3_28_9_i,temp_m3_28_13_r,temp_m3_28_13_i,temp_m3_32_9_r,temp_m3_32_9_i,temp_m3_32_13_r,temp_m3_32_13_i,temp_b3_28_9_r,temp_b3_28_9_i,temp_b3_28_13_r,temp_b3_28_13_i,temp_b3_32_9_r,temp_b3_32_9_i,temp_b3_32_13_r,temp_b3_32_13_i);
MULT MULT734 (clk,temp_b2_28_10_r,temp_b2_28_10_i,temp_b2_28_14_r,temp_b2_28_14_i,temp_b2_32_10_r,temp_b2_32_10_i,temp_b2_32_14_r,temp_b2_32_14_i,temp_m3_28_10_r,temp_m3_28_10_i,temp_m3_28_14_r,temp_m3_28_14_i,temp_m3_32_10_r,temp_m3_32_10_i,temp_m3_32_14_r,temp_m3_32_14_i,`W4_real,`W4_imag,`W12_real,`W12_imag,`W16_real,`W16_imag);
butterfly butterfly734 (clk,temp_m3_28_10_r,temp_m3_28_10_i,temp_m3_28_14_r,temp_m3_28_14_i,temp_m3_32_10_r,temp_m3_32_10_i,temp_m3_32_14_r,temp_m3_32_14_i,temp_b3_28_10_r,temp_b3_28_10_i,temp_b3_28_14_r,temp_b3_28_14_i,temp_b3_32_10_r,temp_b3_32_10_i,temp_b3_32_14_r,temp_b3_32_14_i);
MULT MULT735 (clk,temp_b2_28_11_r,temp_b2_28_11_i,temp_b2_28_15_r,temp_b2_28_15_i,temp_b2_32_11_r,temp_b2_32_11_i,temp_b2_32_15_r,temp_b2_32_15_i,temp_m3_28_11_r,temp_m3_28_11_i,temp_m3_28_15_r,temp_m3_28_15_i,temp_m3_32_11_r,temp_m3_32_11_i,temp_m3_32_15_r,temp_m3_32_15_i,`W8_real,`W8_imag,`W12_real,`W12_imag,`W20_real,`W20_imag);
butterfly butterfly735 (clk,temp_m3_28_11_r,temp_m3_28_11_i,temp_m3_28_15_r,temp_m3_28_15_i,temp_m3_32_11_r,temp_m3_32_11_i,temp_m3_32_15_r,temp_m3_32_15_i,temp_b3_28_11_r,temp_b3_28_11_i,temp_b3_28_15_r,temp_b3_28_15_i,temp_b3_32_11_r,temp_b3_32_11_i,temp_b3_32_15_r,temp_b3_32_15_i);
MULT MULT736 (clk,temp_b2_28_12_r,temp_b2_28_12_i,temp_b2_28_16_r,temp_b2_28_16_i,temp_b2_32_12_r,temp_b2_32_12_i,temp_b2_32_16_r,temp_b2_32_16_i,temp_m3_28_12_r,temp_m3_28_12_i,temp_m3_28_16_r,temp_m3_28_16_i,temp_m3_32_12_r,temp_m3_32_12_i,temp_m3_32_16_r,temp_m3_32_16_i,`W12_real,`W12_imag,`W12_real,`W12_imag,`W24_real,`W24_imag);
butterfly butterfly736 (clk,temp_m3_28_12_r,temp_m3_28_12_i,temp_m3_28_16_r,temp_m3_28_16_i,temp_m3_32_12_r,temp_m3_32_12_i,temp_m3_32_16_r,temp_m3_32_16_i,temp_b3_28_12_r,temp_b3_28_12_i,temp_b3_28_16_r,temp_b3_28_16_i,temp_b3_32_12_r,temp_b3_32_12_i,temp_b3_32_16_r,temp_b3_32_16_i);
MULT MULT737 (clk,temp_b2_25_17_r,temp_b2_25_17_i,temp_b2_25_21_r,temp_b2_25_21_i,temp_b2_29_17_r,temp_b2_29_17_i,temp_b2_29_21_r,temp_b2_29_21_i,temp_m3_25_17_r,temp_m3_25_17_i,temp_m3_25_21_r,temp_m3_25_21_i,temp_m3_29_17_r,temp_m3_29_17_i,temp_m3_29_21_r,temp_m3_29_21_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly737 (clk,temp_m3_25_17_r,temp_m3_25_17_i,temp_m3_25_21_r,temp_m3_25_21_i,temp_m3_29_17_r,temp_m3_29_17_i,temp_m3_29_21_r,temp_m3_29_21_i,temp_b3_25_17_r,temp_b3_25_17_i,temp_b3_25_21_r,temp_b3_25_21_i,temp_b3_29_17_r,temp_b3_29_17_i,temp_b3_29_21_r,temp_b3_29_21_i);
MULT MULT738 (clk,temp_b2_25_18_r,temp_b2_25_18_i,temp_b2_25_22_r,temp_b2_25_22_i,temp_b2_29_18_r,temp_b2_29_18_i,temp_b2_29_22_r,temp_b2_29_22_i,temp_m3_25_18_r,temp_m3_25_18_i,temp_m3_25_22_r,temp_m3_25_22_i,temp_m3_29_18_r,temp_m3_29_18_i,temp_m3_29_22_r,temp_m3_29_22_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly738 (clk,temp_m3_25_18_r,temp_m3_25_18_i,temp_m3_25_22_r,temp_m3_25_22_i,temp_m3_29_18_r,temp_m3_29_18_i,temp_m3_29_22_r,temp_m3_29_22_i,temp_b3_25_18_r,temp_b3_25_18_i,temp_b3_25_22_r,temp_b3_25_22_i,temp_b3_29_18_r,temp_b3_29_18_i,temp_b3_29_22_r,temp_b3_29_22_i);
MULT MULT739 (clk,temp_b2_25_19_r,temp_b2_25_19_i,temp_b2_25_23_r,temp_b2_25_23_i,temp_b2_29_19_r,temp_b2_29_19_i,temp_b2_29_23_r,temp_b2_29_23_i,temp_m3_25_19_r,temp_m3_25_19_i,temp_m3_25_23_r,temp_m3_25_23_i,temp_m3_29_19_r,temp_m3_29_19_i,temp_m3_29_23_r,temp_m3_29_23_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly739 (clk,temp_m3_25_19_r,temp_m3_25_19_i,temp_m3_25_23_r,temp_m3_25_23_i,temp_m3_29_19_r,temp_m3_29_19_i,temp_m3_29_23_r,temp_m3_29_23_i,temp_b3_25_19_r,temp_b3_25_19_i,temp_b3_25_23_r,temp_b3_25_23_i,temp_b3_29_19_r,temp_b3_29_19_i,temp_b3_29_23_r,temp_b3_29_23_i);
MULT MULT740 (clk,temp_b2_25_20_r,temp_b2_25_20_i,temp_b2_25_24_r,temp_b2_25_24_i,temp_b2_29_20_r,temp_b2_29_20_i,temp_b2_29_24_r,temp_b2_29_24_i,temp_m3_25_20_r,temp_m3_25_20_i,temp_m3_25_24_r,temp_m3_25_24_i,temp_m3_29_20_r,temp_m3_29_20_i,temp_m3_29_24_r,temp_m3_29_24_i,`W12_real,`W12_imag,`W0_real,`W0_imag,`W12_real,`W12_imag);
butterfly butterfly740 (clk,temp_m3_25_20_r,temp_m3_25_20_i,temp_m3_25_24_r,temp_m3_25_24_i,temp_m3_29_20_r,temp_m3_29_20_i,temp_m3_29_24_r,temp_m3_29_24_i,temp_b3_25_20_r,temp_b3_25_20_i,temp_b3_25_24_r,temp_b3_25_24_i,temp_b3_29_20_r,temp_b3_29_20_i,temp_b3_29_24_r,temp_b3_29_24_i);
MULT MULT741 (clk,temp_b2_26_17_r,temp_b2_26_17_i,temp_b2_26_21_r,temp_b2_26_21_i,temp_b2_30_17_r,temp_b2_30_17_i,temp_b2_30_21_r,temp_b2_30_21_i,temp_m3_26_17_r,temp_m3_26_17_i,temp_m3_26_21_r,temp_m3_26_21_i,temp_m3_30_17_r,temp_m3_30_17_i,temp_m3_30_21_r,temp_m3_30_21_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly741 (clk,temp_m3_26_17_r,temp_m3_26_17_i,temp_m3_26_21_r,temp_m3_26_21_i,temp_m3_30_17_r,temp_m3_30_17_i,temp_m3_30_21_r,temp_m3_30_21_i,temp_b3_26_17_r,temp_b3_26_17_i,temp_b3_26_21_r,temp_b3_26_21_i,temp_b3_30_17_r,temp_b3_30_17_i,temp_b3_30_21_r,temp_b3_30_21_i);
MULT MULT742 (clk,temp_b2_26_18_r,temp_b2_26_18_i,temp_b2_26_22_r,temp_b2_26_22_i,temp_b2_30_18_r,temp_b2_30_18_i,temp_b2_30_22_r,temp_b2_30_22_i,temp_m3_26_18_r,temp_m3_26_18_i,temp_m3_26_22_r,temp_m3_26_22_i,temp_m3_30_18_r,temp_m3_30_18_i,temp_m3_30_22_r,temp_m3_30_22_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly742 (clk,temp_m3_26_18_r,temp_m3_26_18_i,temp_m3_26_22_r,temp_m3_26_22_i,temp_m3_30_18_r,temp_m3_30_18_i,temp_m3_30_22_r,temp_m3_30_22_i,temp_b3_26_18_r,temp_b3_26_18_i,temp_b3_26_22_r,temp_b3_26_22_i,temp_b3_30_18_r,temp_b3_30_18_i,temp_b3_30_22_r,temp_b3_30_22_i);
MULT MULT743 (clk,temp_b2_26_19_r,temp_b2_26_19_i,temp_b2_26_23_r,temp_b2_26_23_i,temp_b2_30_19_r,temp_b2_30_19_i,temp_b2_30_23_r,temp_b2_30_23_i,temp_m3_26_19_r,temp_m3_26_19_i,temp_m3_26_23_r,temp_m3_26_23_i,temp_m3_30_19_r,temp_m3_30_19_i,temp_m3_30_23_r,temp_m3_30_23_i,`W8_real,`W8_imag,`W4_real,`W4_imag,`W12_real,`W12_imag);
butterfly butterfly743 (clk,temp_m3_26_19_r,temp_m3_26_19_i,temp_m3_26_23_r,temp_m3_26_23_i,temp_m3_30_19_r,temp_m3_30_19_i,temp_m3_30_23_r,temp_m3_30_23_i,temp_b3_26_19_r,temp_b3_26_19_i,temp_b3_26_23_r,temp_b3_26_23_i,temp_b3_30_19_r,temp_b3_30_19_i,temp_b3_30_23_r,temp_b3_30_23_i);
MULT MULT744 (clk,temp_b2_26_20_r,temp_b2_26_20_i,temp_b2_26_24_r,temp_b2_26_24_i,temp_b2_30_20_r,temp_b2_30_20_i,temp_b2_30_24_r,temp_b2_30_24_i,temp_m3_26_20_r,temp_m3_26_20_i,temp_m3_26_24_r,temp_m3_26_24_i,temp_m3_30_20_r,temp_m3_30_20_i,temp_m3_30_24_r,temp_m3_30_24_i,`W12_real,`W12_imag,`W4_real,`W4_imag,`W16_real,`W16_imag);
butterfly butterfly744 (clk,temp_m3_26_20_r,temp_m3_26_20_i,temp_m3_26_24_r,temp_m3_26_24_i,temp_m3_30_20_r,temp_m3_30_20_i,temp_m3_30_24_r,temp_m3_30_24_i,temp_b3_26_20_r,temp_b3_26_20_i,temp_b3_26_24_r,temp_b3_26_24_i,temp_b3_30_20_r,temp_b3_30_20_i,temp_b3_30_24_r,temp_b3_30_24_i);
MULT MULT745 (clk,temp_b2_27_17_r,temp_b2_27_17_i,temp_b2_27_21_r,temp_b2_27_21_i,temp_b2_31_17_r,temp_b2_31_17_i,temp_b2_31_21_r,temp_b2_31_21_i,temp_m3_27_17_r,temp_m3_27_17_i,temp_m3_27_21_r,temp_m3_27_21_i,temp_m3_31_17_r,temp_m3_31_17_i,temp_m3_31_21_r,temp_m3_31_21_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly745 (clk,temp_m3_27_17_r,temp_m3_27_17_i,temp_m3_27_21_r,temp_m3_27_21_i,temp_m3_31_17_r,temp_m3_31_17_i,temp_m3_31_21_r,temp_m3_31_21_i,temp_b3_27_17_r,temp_b3_27_17_i,temp_b3_27_21_r,temp_b3_27_21_i,temp_b3_31_17_r,temp_b3_31_17_i,temp_b3_31_21_r,temp_b3_31_21_i);
MULT MULT746 (clk,temp_b2_27_18_r,temp_b2_27_18_i,temp_b2_27_22_r,temp_b2_27_22_i,temp_b2_31_18_r,temp_b2_31_18_i,temp_b2_31_22_r,temp_b2_31_22_i,temp_m3_27_18_r,temp_m3_27_18_i,temp_m3_27_22_r,temp_m3_27_22_i,temp_m3_31_18_r,temp_m3_31_18_i,temp_m3_31_22_r,temp_m3_31_22_i,`W4_real,`W4_imag,`W8_real,`W8_imag,`W12_real,`W12_imag);
butterfly butterfly746 (clk,temp_m3_27_18_r,temp_m3_27_18_i,temp_m3_27_22_r,temp_m3_27_22_i,temp_m3_31_18_r,temp_m3_31_18_i,temp_m3_31_22_r,temp_m3_31_22_i,temp_b3_27_18_r,temp_b3_27_18_i,temp_b3_27_22_r,temp_b3_27_22_i,temp_b3_31_18_r,temp_b3_31_18_i,temp_b3_31_22_r,temp_b3_31_22_i);
MULT MULT747 (clk,temp_b2_27_19_r,temp_b2_27_19_i,temp_b2_27_23_r,temp_b2_27_23_i,temp_b2_31_19_r,temp_b2_31_19_i,temp_b2_31_23_r,temp_b2_31_23_i,temp_m3_27_19_r,temp_m3_27_19_i,temp_m3_27_23_r,temp_m3_27_23_i,temp_m3_31_19_r,temp_m3_31_19_i,temp_m3_31_23_r,temp_m3_31_23_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly747 (clk,temp_m3_27_19_r,temp_m3_27_19_i,temp_m3_27_23_r,temp_m3_27_23_i,temp_m3_31_19_r,temp_m3_31_19_i,temp_m3_31_23_r,temp_m3_31_23_i,temp_b3_27_19_r,temp_b3_27_19_i,temp_b3_27_23_r,temp_b3_27_23_i,temp_b3_31_19_r,temp_b3_31_19_i,temp_b3_31_23_r,temp_b3_31_23_i);
MULT MULT748 (clk,temp_b2_27_20_r,temp_b2_27_20_i,temp_b2_27_24_r,temp_b2_27_24_i,temp_b2_31_20_r,temp_b2_31_20_i,temp_b2_31_24_r,temp_b2_31_24_i,temp_m3_27_20_r,temp_m3_27_20_i,temp_m3_27_24_r,temp_m3_27_24_i,temp_m3_31_20_r,temp_m3_31_20_i,temp_m3_31_24_r,temp_m3_31_24_i,`W12_real,`W12_imag,`W8_real,`W8_imag,`W20_real,`W20_imag);
butterfly butterfly748 (clk,temp_m3_27_20_r,temp_m3_27_20_i,temp_m3_27_24_r,temp_m3_27_24_i,temp_m3_31_20_r,temp_m3_31_20_i,temp_m3_31_24_r,temp_m3_31_24_i,temp_b3_27_20_r,temp_b3_27_20_i,temp_b3_27_24_r,temp_b3_27_24_i,temp_b3_31_20_r,temp_b3_31_20_i,temp_b3_31_24_r,temp_b3_31_24_i);
MULT MULT749 (clk,temp_b2_28_17_r,temp_b2_28_17_i,temp_b2_28_21_r,temp_b2_28_21_i,temp_b2_32_17_r,temp_b2_32_17_i,temp_b2_32_21_r,temp_b2_32_21_i,temp_m3_28_17_r,temp_m3_28_17_i,temp_m3_28_21_r,temp_m3_28_21_i,temp_m3_32_17_r,temp_m3_32_17_i,temp_m3_32_21_r,temp_m3_32_21_i,`W0_real,`W0_imag,`W12_real,`W12_imag,`W12_real,`W12_imag);
butterfly butterfly749 (clk,temp_m3_28_17_r,temp_m3_28_17_i,temp_m3_28_21_r,temp_m3_28_21_i,temp_m3_32_17_r,temp_m3_32_17_i,temp_m3_32_21_r,temp_m3_32_21_i,temp_b3_28_17_r,temp_b3_28_17_i,temp_b3_28_21_r,temp_b3_28_21_i,temp_b3_32_17_r,temp_b3_32_17_i,temp_b3_32_21_r,temp_b3_32_21_i);
MULT MULT750 (clk,temp_b2_28_18_r,temp_b2_28_18_i,temp_b2_28_22_r,temp_b2_28_22_i,temp_b2_32_18_r,temp_b2_32_18_i,temp_b2_32_22_r,temp_b2_32_22_i,temp_m3_28_18_r,temp_m3_28_18_i,temp_m3_28_22_r,temp_m3_28_22_i,temp_m3_32_18_r,temp_m3_32_18_i,temp_m3_32_22_r,temp_m3_32_22_i,`W4_real,`W4_imag,`W12_real,`W12_imag,`W16_real,`W16_imag);
butterfly butterfly750 (clk,temp_m3_28_18_r,temp_m3_28_18_i,temp_m3_28_22_r,temp_m3_28_22_i,temp_m3_32_18_r,temp_m3_32_18_i,temp_m3_32_22_r,temp_m3_32_22_i,temp_b3_28_18_r,temp_b3_28_18_i,temp_b3_28_22_r,temp_b3_28_22_i,temp_b3_32_18_r,temp_b3_32_18_i,temp_b3_32_22_r,temp_b3_32_22_i);
MULT MULT751 (clk,temp_b2_28_19_r,temp_b2_28_19_i,temp_b2_28_23_r,temp_b2_28_23_i,temp_b2_32_19_r,temp_b2_32_19_i,temp_b2_32_23_r,temp_b2_32_23_i,temp_m3_28_19_r,temp_m3_28_19_i,temp_m3_28_23_r,temp_m3_28_23_i,temp_m3_32_19_r,temp_m3_32_19_i,temp_m3_32_23_r,temp_m3_32_23_i,`W8_real,`W8_imag,`W12_real,`W12_imag,`W20_real,`W20_imag);
butterfly butterfly751 (clk,temp_m3_28_19_r,temp_m3_28_19_i,temp_m3_28_23_r,temp_m3_28_23_i,temp_m3_32_19_r,temp_m3_32_19_i,temp_m3_32_23_r,temp_m3_32_23_i,temp_b3_28_19_r,temp_b3_28_19_i,temp_b3_28_23_r,temp_b3_28_23_i,temp_b3_32_19_r,temp_b3_32_19_i,temp_b3_32_23_r,temp_b3_32_23_i);
MULT MULT752 (clk,temp_b2_28_20_r,temp_b2_28_20_i,temp_b2_28_24_r,temp_b2_28_24_i,temp_b2_32_20_r,temp_b2_32_20_i,temp_b2_32_24_r,temp_b2_32_24_i,temp_m3_28_20_r,temp_m3_28_20_i,temp_m3_28_24_r,temp_m3_28_24_i,temp_m3_32_20_r,temp_m3_32_20_i,temp_m3_32_24_r,temp_m3_32_24_i,`W12_real,`W12_imag,`W12_real,`W12_imag,`W24_real,`W24_imag);
butterfly butterfly752 (clk,temp_m3_28_20_r,temp_m3_28_20_i,temp_m3_28_24_r,temp_m3_28_24_i,temp_m3_32_20_r,temp_m3_32_20_i,temp_m3_32_24_r,temp_m3_32_24_i,temp_b3_28_20_r,temp_b3_28_20_i,temp_b3_28_24_r,temp_b3_28_24_i,temp_b3_32_20_r,temp_b3_32_20_i,temp_b3_32_24_r,temp_b3_32_24_i);
MULT MULT753 (clk,temp_b2_25_25_r,temp_b2_25_25_i,temp_b2_25_29_r,temp_b2_25_29_i,temp_b2_29_25_r,temp_b2_29_25_i,temp_b2_29_29_r,temp_b2_29_29_i,temp_m3_25_25_r,temp_m3_25_25_i,temp_m3_25_29_r,temp_m3_25_29_i,temp_m3_29_25_r,temp_m3_29_25_i,temp_m3_29_29_r,temp_m3_29_29_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly753 (clk,temp_m3_25_25_r,temp_m3_25_25_i,temp_m3_25_29_r,temp_m3_25_29_i,temp_m3_29_25_r,temp_m3_29_25_i,temp_m3_29_29_r,temp_m3_29_29_i,temp_b3_25_25_r,temp_b3_25_25_i,temp_b3_25_29_r,temp_b3_25_29_i,temp_b3_29_25_r,temp_b3_29_25_i,temp_b3_29_29_r,temp_b3_29_29_i);
MULT MULT754 (clk,temp_b2_25_26_r,temp_b2_25_26_i,temp_b2_25_30_r,temp_b2_25_30_i,temp_b2_29_26_r,temp_b2_29_26_i,temp_b2_29_30_r,temp_b2_29_30_i,temp_m3_25_26_r,temp_m3_25_26_i,temp_m3_25_30_r,temp_m3_25_30_i,temp_m3_29_26_r,temp_m3_29_26_i,temp_m3_29_30_r,temp_m3_29_30_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly754 (clk,temp_m3_25_26_r,temp_m3_25_26_i,temp_m3_25_30_r,temp_m3_25_30_i,temp_m3_29_26_r,temp_m3_29_26_i,temp_m3_29_30_r,temp_m3_29_30_i,temp_b3_25_26_r,temp_b3_25_26_i,temp_b3_25_30_r,temp_b3_25_30_i,temp_b3_29_26_r,temp_b3_29_26_i,temp_b3_29_30_r,temp_b3_29_30_i);
MULT MULT755 (clk,temp_b2_25_27_r,temp_b2_25_27_i,temp_b2_25_31_r,temp_b2_25_31_i,temp_b2_29_27_r,temp_b2_29_27_i,temp_b2_29_31_r,temp_b2_29_31_i,temp_m3_25_27_r,temp_m3_25_27_i,temp_m3_25_31_r,temp_m3_25_31_i,temp_m3_29_27_r,temp_m3_29_27_i,temp_m3_29_31_r,temp_m3_29_31_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly755 (clk,temp_m3_25_27_r,temp_m3_25_27_i,temp_m3_25_31_r,temp_m3_25_31_i,temp_m3_29_27_r,temp_m3_29_27_i,temp_m3_29_31_r,temp_m3_29_31_i,temp_b3_25_27_r,temp_b3_25_27_i,temp_b3_25_31_r,temp_b3_25_31_i,temp_b3_29_27_r,temp_b3_29_27_i,temp_b3_29_31_r,temp_b3_29_31_i);
MULT MULT756 (clk,temp_b2_25_28_r,temp_b2_25_28_i,temp_b2_25_32_r,temp_b2_25_32_i,temp_b2_29_28_r,temp_b2_29_28_i,temp_b2_29_32_r,temp_b2_29_32_i,temp_m3_25_28_r,temp_m3_25_28_i,temp_m3_25_32_r,temp_m3_25_32_i,temp_m3_29_28_r,temp_m3_29_28_i,temp_m3_29_32_r,temp_m3_29_32_i,`W12_real,`W12_imag,`W0_real,`W0_imag,`W12_real,`W12_imag);
butterfly butterfly756 (clk,temp_m3_25_28_r,temp_m3_25_28_i,temp_m3_25_32_r,temp_m3_25_32_i,temp_m3_29_28_r,temp_m3_29_28_i,temp_m3_29_32_r,temp_m3_29_32_i,temp_b3_25_28_r,temp_b3_25_28_i,temp_b3_25_32_r,temp_b3_25_32_i,temp_b3_29_28_r,temp_b3_29_28_i,temp_b3_29_32_r,temp_b3_29_32_i);
MULT MULT757 (clk,temp_b2_26_25_r,temp_b2_26_25_i,temp_b2_26_29_r,temp_b2_26_29_i,temp_b2_30_25_r,temp_b2_30_25_i,temp_b2_30_29_r,temp_b2_30_29_i,temp_m3_26_25_r,temp_m3_26_25_i,temp_m3_26_29_r,temp_m3_26_29_i,temp_m3_30_25_r,temp_m3_30_25_i,temp_m3_30_29_r,temp_m3_30_29_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly757 (clk,temp_m3_26_25_r,temp_m3_26_25_i,temp_m3_26_29_r,temp_m3_26_29_i,temp_m3_30_25_r,temp_m3_30_25_i,temp_m3_30_29_r,temp_m3_30_29_i,temp_b3_26_25_r,temp_b3_26_25_i,temp_b3_26_29_r,temp_b3_26_29_i,temp_b3_30_25_r,temp_b3_30_25_i,temp_b3_30_29_r,temp_b3_30_29_i);
MULT MULT758 (clk,temp_b2_26_26_r,temp_b2_26_26_i,temp_b2_26_30_r,temp_b2_26_30_i,temp_b2_30_26_r,temp_b2_30_26_i,temp_b2_30_30_r,temp_b2_30_30_i,temp_m3_26_26_r,temp_m3_26_26_i,temp_m3_26_30_r,temp_m3_26_30_i,temp_m3_30_26_r,temp_m3_30_26_i,temp_m3_30_30_r,temp_m3_30_30_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly758 (clk,temp_m3_26_26_r,temp_m3_26_26_i,temp_m3_26_30_r,temp_m3_26_30_i,temp_m3_30_26_r,temp_m3_30_26_i,temp_m3_30_30_r,temp_m3_30_30_i,temp_b3_26_26_r,temp_b3_26_26_i,temp_b3_26_30_r,temp_b3_26_30_i,temp_b3_30_26_r,temp_b3_30_26_i,temp_b3_30_30_r,temp_b3_30_30_i);
MULT MULT759 (clk,temp_b2_26_27_r,temp_b2_26_27_i,temp_b2_26_31_r,temp_b2_26_31_i,temp_b2_30_27_r,temp_b2_30_27_i,temp_b2_30_31_r,temp_b2_30_31_i,temp_m3_26_27_r,temp_m3_26_27_i,temp_m3_26_31_r,temp_m3_26_31_i,temp_m3_30_27_r,temp_m3_30_27_i,temp_m3_30_31_r,temp_m3_30_31_i,`W8_real,`W8_imag,`W4_real,`W4_imag,`W12_real,`W12_imag);
butterfly butterfly759 (clk,temp_m3_26_27_r,temp_m3_26_27_i,temp_m3_26_31_r,temp_m3_26_31_i,temp_m3_30_27_r,temp_m3_30_27_i,temp_m3_30_31_r,temp_m3_30_31_i,temp_b3_26_27_r,temp_b3_26_27_i,temp_b3_26_31_r,temp_b3_26_31_i,temp_b3_30_27_r,temp_b3_30_27_i,temp_b3_30_31_r,temp_b3_30_31_i);
MULT MULT760 (clk,temp_b2_26_28_r,temp_b2_26_28_i,temp_b2_26_32_r,temp_b2_26_32_i,temp_b2_30_28_r,temp_b2_30_28_i,temp_b2_30_32_r,temp_b2_30_32_i,temp_m3_26_28_r,temp_m3_26_28_i,temp_m3_26_32_r,temp_m3_26_32_i,temp_m3_30_28_r,temp_m3_30_28_i,temp_m3_30_32_r,temp_m3_30_32_i,`W12_real,`W12_imag,`W4_real,`W4_imag,`W16_real,`W16_imag);
butterfly butterfly760 (clk,temp_m3_26_28_r,temp_m3_26_28_i,temp_m3_26_32_r,temp_m3_26_32_i,temp_m3_30_28_r,temp_m3_30_28_i,temp_m3_30_32_r,temp_m3_30_32_i,temp_b3_26_28_r,temp_b3_26_28_i,temp_b3_26_32_r,temp_b3_26_32_i,temp_b3_30_28_r,temp_b3_30_28_i,temp_b3_30_32_r,temp_b3_30_32_i);
MULT MULT761 (clk,temp_b2_27_25_r,temp_b2_27_25_i,temp_b2_27_29_r,temp_b2_27_29_i,temp_b2_31_25_r,temp_b2_31_25_i,temp_b2_31_29_r,temp_b2_31_29_i,temp_m3_27_25_r,temp_m3_27_25_i,temp_m3_27_29_r,temp_m3_27_29_i,temp_m3_31_25_r,temp_m3_31_25_i,temp_m3_31_29_r,temp_m3_31_29_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly761 (clk,temp_m3_27_25_r,temp_m3_27_25_i,temp_m3_27_29_r,temp_m3_27_29_i,temp_m3_31_25_r,temp_m3_31_25_i,temp_m3_31_29_r,temp_m3_31_29_i,temp_b3_27_25_r,temp_b3_27_25_i,temp_b3_27_29_r,temp_b3_27_29_i,temp_b3_31_25_r,temp_b3_31_25_i,temp_b3_31_29_r,temp_b3_31_29_i);
MULT MULT762 (clk,temp_b2_27_26_r,temp_b2_27_26_i,temp_b2_27_30_r,temp_b2_27_30_i,temp_b2_31_26_r,temp_b2_31_26_i,temp_b2_31_30_r,temp_b2_31_30_i,temp_m3_27_26_r,temp_m3_27_26_i,temp_m3_27_30_r,temp_m3_27_30_i,temp_m3_31_26_r,temp_m3_31_26_i,temp_m3_31_30_r,temp_m3_31_30_i,`W4_real,`W4_imag,`W8_real,`W8_imag,`W12_real,`W12_imag);
butterfly butterfly762 (clk,temp_m3_27_26_r,temp_m3_27_26_i,temp_m3_27_30_r,temp_m3_27_30_i,temp_m3_31_26_r,temp_m3_31_26_i,temp_m3_31_30_r,temp_m3_31_30_i,temp_b3_27_26_r,temp_b3_27_26_i,temp_b3_27_30_r,temp_b3_27_30_i,temp_b3_31_26_r,temp_b3_31_26_i,temp_b3_31_30_r,temp_b3_31_30_i);
MULT MULT763 (clk,temp_b2_27_27_r,temp_b2_27_27_i,temp_b2_27_31_r,temp_b2_27_31_i,temp_b2_31_27_r,temp_b2_31_27_i,temp_b2_31_31_r,temp_b2_31_31_i,temp_m3_27_27_r,temp_m3_27_27_i,temp_m3_27_31_r,temp_m3_27_31_i,temp_m3_31_27_r,temp_m3_31_27_i,temp_m3_31_31_r,temp_m3_31_31_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly763 (clk,temp_m3_27_27_r,temp_m3_27_27_i,temp_m3_27_31_r,temp_m3_27_31_i,temp_m3_31_27_r,temp_m3_31_27_i,temp_m3_31_31_r,temp_m3_31_31_i,temp_b3_27_27_r,temp_b3_27_27_i,temp_b3_27_31_r,temp_b3_27_31_i,temp_b3_31_27_r,temp_b3_31_27_i,temp_b3_31_31_r,temp_b3_31_31_i);
MULT MULT764 (clk,temp_b2_27_28_r,temp_b2_27_28_i,temp_b2_27_32_r,temp_b2_27_32_i,temp_b2_31_28_r,temp_b2_31_28_i,temp_b2_31_32_r,temp_b2_31_32_i,temp_m3_27_28_r,temp_m3_27_28_i,temp_m3_27_32_r,temp_m3_27_32_i,temp_m3_31_28_r,temp_m3_31_28_i,temp_m3_31_32_r,temp_m3_31_32_i,`W12_real,`W12_imag,`W8_real,`W8_imag,`W20_real,`W20_imag);
butterfly butterfly764 (clk,temp_m3_27_28_r,temp_m3_27_28_i,temp_m3_27_32_r,temp_m3_27_32_i,temp_m3_31_28_r,temp_m3_31_28_i,temp_m3_31_32_r,temp_m3_31_32_i,temp_b3_27_28_r,temp_b3_27_28_i,temp_b3_27_32_r,temp_b3_27_32_i,temp_b3_31_28_r,temp_b3_31_28_i,temp_b3_31_32_r,temp_b3_31_32_i);
MULT MULT765 (clk,temp_b2_28_25_r,temp_b2_28_25_i,temp_b2_28_29_r,temp_b2_28_29_i,temp_b2_32_25_r,temp_b2_32_25_i,temp_b2_32_29_r,temp_b2_32_29_i,temp_m3_28_25_r,temp_m3_28_25_i,temp_m3_28_29_r,temp_m3_28_29_i,temp_m3_32_25_r,temp_m3_32_25_i,temp_m3_32_29_r,temp_m3_32_29_i,`W0_real,`W0_imag,`W12_real,`W12_imag,`W12_real,`W12_imag);
butterfly butterfly765 (clk,temp_m3_28_25_r,temp_m3_28_25_i,temp_m3_28_29_r,temp_m3_28_29_i,temp_m3_32_25_r,temp_m3_32_25_i,temp_m3_32_29_r,temp_m3_32_29_i,temp_b3_28_25_r,temp_b3_28_25_i,temp_b3_28_29_r,temp_b3_28_29_i,temp_b3_32_25_r,temp_b3_32_25_i,temp_b3_32_29_r,temp_b3_32_29_i);
MULT MULT766 (clk,temp_b2_28_26_r,temp_b2_28_26_i,temp_b2_28_30_r,temp_b2_28_30_i,temp_b2_32_26_r,temp_b2_32_26_i,temp_b2_32_30_r,temp_b2_32_30_i,temp_m3_28_26_r,temp_m3_28_26_i,temp_m3_28_30_r,temp_m3_28_30_i,temp_m3_32_26_r,temp_m3_32_26_i,temp_m3_32_30_r,temp_m3_32_30_i,`W4_real,`W4_imag,`W12_real,`W12_imag,`W16_real,`W16_imag);
butterfly butterfly766 (clk,temp_m3_28_26_r,temp_m3_28_26_i,temp_m3_28_30_r,temp_m3_28_30_i,temp_m3_32_26_r,temp_m3_32_26_i,temp_m3_32_30_r,temp_m3_32_30_i,temp_b3_28_26_r,temp_b3_28_26_i,temp_b3_28_30_r,temp_b3_28_30_i,temp_b3_32_26_r,temp_b3_32_26_i,temp_b3_32_30_r,temp_b3_32_30_i);
MULT MULT767 (clk,temp_b2_28_27_r,temp_b2_28_27_i,temp_b2_28_31_r,temp_b2_28_31_i,temp_b2_32_27_r,temp_b2_32_27_i,temp_b2_32_31_r,temp_b2_32_31_i,temp_m3_28_27_r,temp_m3_28_27_i,temp_m3_28_31_r,temp_m3_28_31_i,temp_m3_32_27_r,temp_m3_32_27_i,temp_m3_32_31_r,temp_m3_32_31_i,`W8_real,`W8_imag,`W12_real,`W12_imag,`W20_real,`W20_imag);
butterfly butterfly767 (clk,temp_m3_28_27_r,temp_m3_28_27_i,temp_m3_28_31_r,temp_m3_28_31_i,temp_m3_32_27_r,temp_m3_32_27_i,temp_m3_32_31_r,temp_m3_32_31_i,temp_b3_28_27_r,temp_b3_28_27_i,temp_b3_28_31_r,temp_b3_28_31_i,temp_b3_32_27_r,temp_b3_32_27_i,temp_b3_32_31_r,temp_b3_32_31_i);
MULT MULT768 (clk,temp_b2_28_28_r,temp_b2_28_28_i,temp_b2_28_32_r,temp_b2_28_32_i,temp_b2_32_28_r,temp_b2_32_28_i,temp_b2_32_32_r,temp_b2_32_32_i,temp_m3_28_28_r,temp_m3_28_28_i,temp_m3_28_32_r,temp_m3_28_32_i,temp_m3_32_28_r,temp_m3_32_28_i,temp_m3_32_32_r,temp_m3_32_32_i,`W12_real,`W12_imag,`W12_real,`W12_imag,`W24_real,`W24_imag);
butterfly butterfly768 (clk,temp_m3_28_28_r,temp_m3_28_28_i,temp_m3_28_32_r,temp_m3_28_32_i,temp_m3_32_28_r,temp_m3_32_28_i,temp_m3_32_32_r,temp_m3_32_32_i,temp_b3_28_28_r,temp_b3_28_28_i,temp_b3_28_32_r,temp_b3_28_32_i,temp_b3_32_28_r,temp_b3_32_28_i,temp_b3_32_32_r,temp_b3_32_32_i);
MULT MULT769 (clk,temp_b3_1_1_r,temp_b3_1_1_i,temp_b3_1_9_r,temp_b3_1_9_i,temp_b3_9_1_r,temp_b3_9_1_i,temp_b3_9_9_r,temp_b3_9_9_i,temp_m4_1_1_r,temp_m4_1_1_i,temp_m4_1_9_r,temp_m4_1_9_i,temp_m4_9_1_r,temp_m4_9_1_i,temp_m4_9_9_r,temp_m4_9_9_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly769 (clk,temp_m4_1_1_r,temp_m4_1_1_i,temp_m4_1_9_r,temp_m4_1_9_i,temp_m4_9_1_r,temp_m4_9_1_i,temp_m4_9_9_r,temp_m4_9_9_i,temp_b4_1_1_r,temp_b4_1_1_i,temp_b4_1_9_r,temp_b4_1_9_i,temp_b4_9_1_r,temp_b4_9_1_i,temp_b4_9_9_r,temp_b4_9_9_i);
MULT MULT770 (clk,temp_b3_1_2_r,temp_b3_1_2_i,temp_b3_1_10_r,temp_b3_1_10_i,temp_b3_9_2_r,temp_b3_9_2_i,temp_b3_9_10_r,temp_b3_9_10_i,temp_m4_1_2_r,temp_m4_1_2_i,temp_m4_1_10_r,temp_m4_1_10_i,temp_m4_9_2_r,temp_m4_9_2_i,temp_m4_9_10_r,temp_m4_9_10_i,`W2_real,`W2_imag,`W0_real,`W0_imag,`W2_real,`W2_imag);
butterfly butterfly770 (clk,temp_m4_1_2_r,temp_m4_1_2_i,temp_m4_1_10_r,temp_m4_1_10_i,temp_m4_9_2_r,temp_m4_9_2_i,temp_m4_9_10_r,temp_m4_9_10_i,temp_b4_1_2_r,temp_b4_1_2_i,temp_b4_1_10_r,temp_b4_1_10_i,temp_b4_9_2_r,temp_b4_9_2_i,temp_b4_9_10_r,temp_b4_9_10_i);
MULT MULT771 (clk,temp_b3_1_3_r,temp_b3_1_3_i,temp_b3_1_11_r,temp_b3_1_11_i,temp_b3_9_3_r,temp_b3_9_3_i,temp_b3_9_11_r,temp_b3_9_11_i,temp_m4_1_3_r,temp_m4_1_3_i,temp_m4_1_11_r,temp_m4_1_11_i,temp_m4_9_3_r,temp_m4_9_3_i,temp_m4_9_11_r,temp_m4_9_11_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly771 (clk,temp_m4_1_3_r,temp_m4_1_3_i,temp_m4_1_11_r,temp_m4_1_11_i,temp_m4_9_3_r,temp_m4_9_3_i,temp_m4_9_11_r,temp_m4_9_11_i,temp_b4_1_3_r,temp_b4_1_3_i,temp_b4_1_11_r,temp_b4_1_11_i,temp_b4_9_3_r,temp_b4_9_3_i,temp_b4_9_11_r,temp_b4_9_11_i);
MULT MULT772 (clk,temp_b3_1_4_r,temp_b3_1_4_i,temp_b3_1_12_r,temp_b3_1_12_i,temp_b3_9_4_r,temp_b3_9_4_i,temp_b3_9_12_r,temp_b3_9_12_i,temp_m4_1_4_r,temp_m4_1_4_i,temp_m4_1_12_r,temp_m4_1_12_i,temp_m4_9_4_r,temp_m4_9_4_i,temp_m4_9_12_r,temp_m4_9_12_i,`W6_real,`W6_imag,`W0_real,`W0_imag,`W6_real,`W6_imag);
butterfly butterfly772 (clk,temp_m4_1_4_r,temp_m4_1_4_i,temp_m4_1_12_r,temp_m4_1_12_i,temp_m4_9_4_r,temp_m4_9_4_i,temp_m4_9_12_r,temp_m4_9_12_i,temp_b4_1_4_r,temp_b4_1_4_i,temp_b4_1_12_r,temp_b4_1_12_i,temp_b4_9_4_r,temp_b4_9_4_i,temp_b4_9_12_r,temp_b4_9_12_i);
MULT MULT773 (clk,temp_b3_1_5_r,temp_b3_1_5_i,temp_b3_1_13_r,temp_b3_1_13_i,temp_b3_9_5_r,temp_b3_9_5_i,temp_b3_9_13_r,temp_b3_9_13_i,temp_m4_1_5_r,temp_m4_1_5_i,temp_m4_1_13_r,temp_m4_1_13_i,temp_m4_9_5_r,temp_m4_9_5_i,temp_m4_9_13_r,temp_m4_9_13_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly773 (clk,temp_m4_1_5_r,temp_m4_1_5_i,temp_m4_1_13_r,temp_m4_1_13_i,temp_m4_9_5_r,temp_m4_9_5_i,temp_m4_9_13_r,temp_m4_9_13_i,temp_b4_1_5_r,temp_b4_1_5_i,temp_b4_1_13_r,temp_b4_1_13_i,temp_b4_9_5_r,temp_b4_9_5_i,temp_b4_9_13_r,temp_b4_9_13_i);
MULT MULT774 (clk,temp_b3_1_6_r,temp_b3_1_6_i,temp_b3_1_14_r,temp_b3_1_14_i,temp_b3_9_6_r,temp_b3_9_6_i,temp_b3_9_14_r,temp_b3_9_14_i,temp_m4_1_6_r,temp_m4_1_6_i,temp_m4_1_14_r,temp_m4_1_14_i,temp_m4_9_6_r,temp_m4_9_6_i,temp_m4_9_14_r,temp_m4_9_14_i,`W10_real,`W10_imag,`W0_real,`W0_imag,`W10_real,`W10_imag);
butterfly butterfly774 (clk,temp_m4_1_6_r,temp_m4_1_6_i,temp_m4_1_14_r,temp_m4_1_14_i,temp_m4_9_6_r,temp_m4_9_6_i,temp_m4_9_14_r,temp_m4_9_14_i,temp_b4_1_6_r,temp_b4_1_6_i,temp_b4_1_14_r,temp_b4_1_14_i,temp_b4_9_6_r,temp_b4_9_6_i,temp_b4_9_14_r,temp_b4_9_14_i);
MULT MULT775 (clk,temp_b3_1_7_r,temp_b3_1_7_i,temp_b3_1_15_r,temp_b3_1_15_i,temp_b3_9_7_r,temp_b3_9_7_i,temp_b3_9_15_r,temp_b3_9_15_i,temp_m4_1_7_r,temp_m4_1_7_i,temp_m4_1_15_r,temp_m4_1_15_i,temp_m4_9_7_r,temp_m4_9_7_i,temp_m4_9_15_r,temp_m4_9_15_i,`W12_real,`W12_imag,`W0_real,`W0_imag,`W12_real,`W12_imag);
butterfly butterfly775 (clk,temp_m4_1_7_r,temp_m4_1_7_i,temp_m4_1_15_r,temp_m4_1_15_i,temp_m4_9_7_r,temp_m4_9_7_i,temp_m4_9_15_r,temp_m4_9_15_i,temp_b4_1_7_r,temp_b4_1_7_i,temp_b4_1_15_r,temp_b4_1_15_i,temp_b4_9_7_r,temp_b4_9_7_i,temp_b4_9_15_r,temp_b4_9_15_i);
MULT MULT776 (clk,temp_b3_1_8_r,temp_b3_1_8_i,temp_b3_1_16_r,temp_b3_1_16_i,temp_b3_9_8_r,temp_b3_9_8_i,temp_b3_9_16_r,temp_b3_9_16_i,temp_m4_1_8_r,temp_m4_1_8_i,temp_m4_1_16_r,temp_m4_1_16_i,temp_m4_9_8_r,temp_m4_9_8_i,temp_m4_9_16_r,temp_m4_9_16_i,`W14_real,`W14_imag,`W0_real,`W0_imag,`W14_real,`W14_imag);
butterfly butterfly776 (clk,temp_m4_1_8_r,temp_m4_1_8_i,temp_m4_1_16_r,temp_m4_1_16_i,temp_m4_9_8_r,temp_m4_9_8_i,temp_m4_9_16_r,temp_m4_9_16_i,temp_b4_1_8_r,temp_b4_1_8_i,temp_b4_1_16_r,temp_b4_1_16_i,temp_b4_9_8_r,temp_b4_9_8_i,temp_b4_9_16_r,temp_b4_9_16_i);
MULT MULT777 (clk,temp_b3_2_1_r,temp_b3_2_1_i,temp_b3_2_9_r,temp_b3_2_9_i,temp_b3_10_1_r,temp_b3_10_1_i,temp_b3_10_9_r,temp_b3_10_9_i,temp_m4_2_1_r,temp_m4_2_1_i,temp_m4_2_9_r,temp_m4_2_9_i,temp_m4_10_1_r,temp_m4_10_1_i,temp_m4_10_9_r,temp_m4_10_9_i,`W0_real,`W0_imag,`W2_real,`W2_imag,`W2_real,`W2_imag);
butterfly butterfly777 (clk,temp_m4_2_1_r,temp_m4_2_1_i,temp_m4_2_9_r,temp_m4_2_9_i,temp_m4_10_1_r,temp_m4_10_1_i,temp_m4_10_9_r,temp_m4_10_9_i,temp_b4_2_1_r,temp_b4_2_1_i,temp_b4_2_9_r,temp_b4_2_9_i,temp_b4_10_1_r,temp_b4_10_1_i,temp_b4_10_9_r,temp_b4_10_9_i);
MULT MULT778 (clk,temp_b3_2_2_r,temp_b3_2_2_i,temp_b3_2_10_r,temp_b3_2_10_i,temp_b3_10_2_r,temp_b3_10_2_i,temp_b3_10_10_r,temp_b3_10_10_i,temp_m4_2_2_r,temp_m4_2_2_i,temp_m4_2_10_r,temp_m4_2_10_i,temp_m4_10_2_r,temp_m4_10_2_i,temp_m4_10_10_r,temp_m4_10_10_i,`W2_real,`W2_imag,`W2_real,`W2_imag,`W4_real,`W4_imag);
butterfly butterfly778 (clk,temp_m4_2_2_r,temp_m4_2_2_i,temp_m4_2_10_r,temp_m4_2_10_i,temp_m4_10_2_r,temp_m4_10_2_i,temp_m4_10_10_r,temp_m4_10_10_i,temp_b4_2_2_r,temp_b4_2_2_i,temp_b4_2_10_r,temp_b4_2_10_i,temp_b4_10_2_r,temp_b4_10_2_i,temp_b4_10_10_r,temp_b4_10_10_i);
MULT MULT779 (clk,temp_b3_2_3_r,temp_b3_2_3_i,temp_b3_2_11_r,temp_b3_2_11_i,temp_b3_10_3_r,temp_b3_10_3_i,temp_b3_10_11_r,temp_b3_10_11_i,temp_m4_2_3_r,temp_m4_2_3_i,temp_m4_2_11_r,temp_m4_2_11_i,temp_m4_10_3_r,temp_m4_10_3_i,temp_m4_10_11_r,temp_m4_10_11_i,`W4_real,`W4_imag,`W2_real,`W2_imag,`W6_real,`W6_imag);
butterfly butterfly779 (clk,temp_m4_2_3_r,temp_m4_2_3_i,temp_m4_2_11_r,temp_m4_2_11_i,temp_m4_10_3_r,temp_m4_10_3_i,temp_m4_10_11_r,temp_m4_10_11_i,temp_b4_2_3_r,temp_b4_2_3_i,temp_b4_2_11_r,temp_b4_2_11_i,temp_b4_10_3_r,temp_b4_10_3_i,temp_b4_10_11_r,temp_b4_10_11_i);
MULT MULT780 (clk,temp_b3_2_4_r,temp_b3_2_4_i,temp_b3_2_12_r,temp_b3_2_12_i,temp_b3_10_4_r,temp_b3_10_4_i,temp_b3_10_12_r,temp_b3_10_12_i,temp_m4_2_4_r,temp_m4_2_4_i,temp_m4_2_12_r,temp_m4_2_12_i,temp_m4_10_4_r,temp_m4_10_4_i,temp_m4_10_12_r,temp_m4_10_12_i,`W6_real,`W6_imag,`W2_real,`W2_imag,`W8_real,`W8_imag);
butterfly butterfly780 (clk,temp_m4_2_4_r,temp_m4_2_4_i,temp_m4_2_12_r,temp_m4_2_12_i,temp_m4_10_4_r,temp_m4_10_4_i,temp_m4_10_12_r,temp_m4_10_12_i,temp_b4_2_4_r,temp_b4_2_4_i,temp_b4_2_12_r,temp_b4_2_12_i,temp_b4_10_4_r,temp_b4_10_4_i,temp_b4_10_12_r,temp_b4_10_12_i);
MULT MULT781 (clk,temp_b3_2_5_r,temp_b3_2_5_i,temp_b3_2_13_r,temp_b3_2_13_i,temp_b3_10_5_r,temp_b3_10_5_i,temp_b3_10_13_r,temp_b3_10_13_i,temp_m4_2_5_r,temp_m4_2_5_i,temp_m4_2_13_r,temp_m4_2_13_i,temp_m4_10_5_r,temp_m4_10_5_i,temp_m4_10_13_r,temp_m4_10_13_i,`W8_real,`W8_imag,`W2_real,`W2_imag,`W10_real,`W10_imag);
butterfly butterfly781 (clk,temp_m4_2_5_r,temp_m4_2_5_i,temp_m4_2_13_r,temp_m4_2_13_i,temp_m4_10_5_r,temp_m4_10_5_i,temp_m4_10_13_r,temp_m4_10_13_i,temp_b4_2_5_r,temp_b4_2_5_i,temp_b4_2_13_r,temp_b4_2_13_i,temp_b4_10_5_r,temp_b4_10_5_i,temp_b4_10_13_r,temp_b4_10_13_i);
MULT MULT782 (clk,temp_b3_2_6_r,temp_b3_2_6_i,temp_b3_2_14_r,temp_b3_2_14_i,temp_b3_10_6_r,temp_b3_10_6_i,temp_b3_10_14_r,temp_b3_10_14_i,temp_m4_2_6_r,temp_m4_2_6_i,temp_m4_2_14_r,temp_m4_2_14_i,temp_m4_10_6_r,temp_m4_10_6_i,temp_m4_10_14_r,temp_m4_10_14_i,`W10_real,`W10_imag,`W2_real,`W2_imag,`W12_real,`W12_imag);
butterfly butterfly782 (clk,temp_m4_2_6_r,temp_m4_2_6_i,temp_m4_2_14_r,temp_m4_2_14_i,temp_m4_10_6_r,temp_m4_10_6_i,temp_m4_10_14_r,temp_m4_10_14_i,temp_b4_2_6_r,temp_b4_2_6_i,temp_b4_2_14_r,temp_b4_2_14_i,temp_b4_10_6_r,temp_b4_10_6_i,temp_b4_10_14_r,temp_b4_10_14_i);
MULT MULT783 (clk,temp_b3_2_7_r,temp_b3_2_7_i,temp_b3_2_15_r,temp_b3_2_15_i,temp_b3_10_7_r,temp_b3_10_7_i,temp_b3_10_15_r,temp_b3_10_15_i,temp_m4_2_7_r,temp_m4_2_7_i,temp_m4_2_15_r,temp_m4_2_15_i,temp_m4_10_7_r,temp_m4_10_7_i,temp_m4_10_15_r,temp_m4_10_15_i,`W12_real,`W12_imag,`W2_real,`W2_imag,`W14_real,`W14_imag);
butterfly butterfly783 (clk,temp_m4_2_7_r,temp_m4_2_7_i,temp_m4_2_15_r,temp_m4_2_15_i,temp_m4_10_7_r,temp_m4_10_7_i,temp_m4_10_15_r,temp_m4_10_15_i,temp_b4_2_7_r,temp_b4_2_7_i,temp_b4_2_15_r,temp_b4_2_15_i,temp_b4_10_7_r,temp_b4_10_7_i,temp_b4_10_15_r,temp_b4_10_15_i);
MULT MULT784 (clk,temp_b3_2_8_r,temp_b3_2_8_i,temp_b3_2_16_r,temp_b3_2_16_i,temp_b3_10_8_r,temp_b3_10_8_i,temp_b3_10_16_r,temp_b3_10_16_i,temp_m4_2_8_r,temp_m4_2_8_i,temp_m4_2_16_r,temp_m4_2_16_i,temp_m4_10_8_r,temp_m4_10_8_i,temp_m4_10_16_r,temp_m4_10_16_i,`W14_real,`W14_imag,`W2_real,`W2_imag,`W16_real,`W16_imag);
butterfly butterfly784 (clk,temp_m4_2_8_r,temp_m4_2_8_i,temp_m4_2_16_r,temp_m4_2_16_i,temp_m4_10_8_r,temp_m4_10_8_i,temp_m4_10_16_r,temp_m4_10_16_i,temp_b4_2_8_r,temp_b4_2_8_i,temp_b4_2_16_r,temp_b4_2_16_i,temp_b4_10_8_r,temp_b4_10_8_i,temp_b4_10_16_r,temp_b4_10_16_i);
MULT MULT785 (clk,temp_b3_3_1_r,temp_b3_3_1_i,temp_b3_3_9_r,temp_b3_3_9_i,temp_b3_11_1_r,temp_b3_11_1_i,temp_b3_11_9_r,temp_b3_11_9_i,temp_m4_3_1_r,temp_m4_3_1_i,temp_m4_3_9_r,temp_m4_3_9_i,temp_m4_11_1_r,temp_m4_11_1_i,temp_m4_11_9_r,temp_m4_11_9_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly785 (clk,temp_m4_3_1_r,temp_m4_3_1_i,temp_m4_3_9_r,temp_m4_3_9_i,temp_m4_11_1_r,temp_m4_11_1_i,temp_m4_11_9_r,temp_m4_11_9_i,temp_b4_3_1_r,temp_b4_3_1_i,temp_b4_3_9_r,temp_b4_3_9_i,temp_b4_11_1_r,temp_b4_11_1_i,temp_b4_11_9_r,temp_b4_11_9_i);
MULT MULT786 (clk,temp_b3_3_2_r,temp_b3_3_2_i,temp_b3_3_10_r,temp_b3_3_10_i,temp_b3_11_2_r,temp_b3_11_2_i,temp_b3_11_10_r,temp_b3_11_10_i,temp_m4_3_2_r,temp_m4_3_2_i,temp_m4_3_10_r,temp_m4_3_10_i,temp_m4_11_2_r,temp_m4_11_2_i,temp_m4_11_10_r,temp_m4_11_10_i,`W2_real,`W2_imag,`W4_real,`W4_imag,`W6_real,`W6_imag);
butterfly butterfly786 (clk,temp_m4_3_2_r,temp_m4_3_2_i,temp_m4_3_10_r,temp_m4_3_10_i,temp_m4_11_2_r,temp_m4_11_2_i,temp_m4_11_10_r,temp_m4_11_10_i,temp_b4_3_2_r,temp_b4_3_2_i,temp_b4_3_10_r,temp_b4_3_10_i,temp_b4_11_2_r,temp_b4_11_2_i,temp_b4_11_10_r,temp_b4_11_10_i);
MULT MULT787 (clk,temp_b3_3_3_r,temp_b3_3_3_i,temp_b3_3_11_r,temp_b3_3_11_i,temp_b3_11_3_r,temp_b3_11_3_i,temp_b3_11_11_r,temp_b3_11_11_i,temp_m4_3_3_r,temp_m4_3_3_i,temp_m4_3_11_r,temp_m4_3_11_i,temp_m4_11_3_r,temp_m4_11_3_i,temp_m4_11_11_r,temp_m4_11_11_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly787 (clk,temp_m4_3_3_r,temp_m4_3_3_i,temp_m4_3_11_r,temp_m4_3_11_i,temp_m4_11_3_r,temp_m4_11_3_i,temp_m4_11_11_r,temp_m4_11_11_i,temp_b4_3_3_r,temp_b4_3_3_i,temp_b4_3_11_r,temp_b4_3_11_i,temp_b4_11_3_r,temp_b4_11_3_i,temp_b4_11_11_r,temp_b4_11_11_i);
MULT MULT788 (clk,temp_b3_3_4_r,temp_b3_3_4_i,temp_b3_3_12_r,temp_b3_3_12_i,temp_b3_11_4_r,temp_b3_11_4_i,temp_b3_11_12_r,temp_b3_11_12_i,temp_m4_3_4_r,temp_m4_3_4_i,temp_m4_3_12_r,temp_m4_3_12_i,temp_m4_11_4_r,temp_m4_11_4_i,temp_m4_11_12_r,temp_m4_11_12_i,`W6_real,`W6_imag,`W4_real,`W4_imag,`W10_real,`W10_imag);
butterfly butterfly788 (clk,temp_m4_3_4_r,temp_m4_3_4_i,temp_m4_3_12_r,temp_m4_3_12_i,temp_m4_11_4_r,temp_m4_11_4_i,temp_m4_11_12_r,temp_m4_11_12_i,temp_b4_3_4_r,temp_b4_3_4_i,temp_b4_3_12_r,temp_b4_3_12_i,temp_b4_11_4_r,temp_b4_11_4_i,temp_b4_11_12_r,temp_b4_11_12_i);
MULT MULT789 (clk,temp_b3_3_5_r,temp_b3_3_5_i,temp_b3_3_13_r,temp_b3_3_13_i,temp_b3_11_5_r,temp_b3_11_5_i,temp_b3_11_13_r,temp_b3_11_13_i,temp_m4_3_5_r,temp_m4_3_5_i,temp_m4_3_13_r,temp_m4_3_13_i,temp_m4_11_5_r,temp_m4_11_5_i,temp_m4_11_13_r,temp_m4_11_13_i,`W8_real,`W8_imag,`W4_real,`W4_imag,`W12_real,`W12_imag);
butterfly butterfly789 (clk,temp_m4_3_5_r,temp_m4_3_5_i,temp_m4_3_13_r,temp_m4_3_13_i,temp_m4_11_5_r,temp_m4_11_5_i,temp_m4_11_13_r,temp_m4_11_13_i,temp_b4_3_5_r,temp_b4_3_5_i,temp_b4_3_13_r,temp_b4_3_13_i,temp_b4_11_5_r,temp_b4_11_5_i,temp_b4_11_13_r,temp_b4_11_13_i);
MULT MULT790 (clk,temp_b3_3_6_r,temp_b3_3_6_i,temp_b3_3_14_r,temp_b3_3_14_i,temp_b3_11_6_r,temp_b3_11_6_i,temp_b3_11_14_r,temp_b3_11_14_i,temp_m4_3_6_r,temp_m4_3_6_i,temp_m4_3_14_r,temp_m4_3_14_i,temp_m4_11_6_r,temp_m4_11_6_i,temp_m4_11_14_r,temp_m4_11_14_i,`W10_real,`W10_imag,`W4_real,`W4_imag,`W14_real,`W14_imag);
butterfly butterfly790 (clk,temp_m4_3_6_r,temp_m4_3_6_i,temp_m4_3_14_r,temp_m4_3_14_i,temp_m4_11_6_r,temp_m4_11_6_i,temp_m4_11_14_r,temp_m4_11_14_i,temp_b4_3_6_r,temp_b4_3_6_i,temp_b4_3_14_r,temp_b4_3_14_i,temp_b4_11_6_r,temp_b4_11_6_i,temp_b4_11_14_r,temp_b4_11_14_i);
MULT MULT791 (clk,temp_b3_3_7_r,temp_b3_3_7_i,temp_b3_3_15_r,temp_b3_3_15_i,temp_b3_11_7_r,temp_b3_11_7_i,temp_b3_11_15_r,temp_b3_11_15_i,temp_m4_3_7_r,temp_m4_3_7_i,temp_m4_3_15_r,temp_m4_3_15_i,temp_m4_11_7_r,temp_m4_11_7_i,temp_m4_11_15_r,temp_m4_11_15_i,`W12_real,`W12_imag,`W4_real,`W4_imag,`W16_real,`W16_imag);
butterfly butterfly791 (clk,temp_m4_3_7_r,temp_m4_3_7_i,temp_m4_3_15_r,temp_m4_3_15_i,temp_m4_11_7_r,temp_m4_11_7_i,temp_m4_11_15_r,temp_m4_11_15_i,temp_b4_3_7_r,temp_b4_3_7_i,temp_b4_3_15_r,temp_b4_3_15_i,temp_b4_11_7_r,temp_b4_11_7_i,temp_b4_11_15_r,temp_b4_11_15_i);
MULT MULT792 (clk,temp_b3_3_8_r,temp_b3_3_8_i,temp_b3_3_16_r,temp_b3_3_16_i,temp_b3_11_8_r,temp_b3_11_8_i,temp_b3_11_16_r,temp_b3_11_16_i,temp_m4_3_8_r,temp_m4_3_8_i,temp_m4_3_16_r,temp_m4_3_16_i,temp_m4_11_8_r,temp_m4_11_8_i,temp_m4_11_16_r,temp_m4_11_16_i,`W14_real,`W14_imag,`W4_real,`W4_imag,`W18_real,`W18_imag);
butterfly butterfly792 (clk,temp_m4_3_8_r,temp_m4_3_8_i,temp_m4_3_16_r,temp_m4_3_16_i,temp_m4_11_8_r,temp_m4_11_8_i,temp_m4_11_16_r,temp_m4_11_16_i,temp_b4_3_8_r,temp_b4_3_8_i,temp_b4_3_16_r,temp_b4_3_16_i,temp_b4_11_8_r,temp_b4_11_8_i,temp_b4_11_16_r,temp_b4_11_16_i);
MULT MULT793 (clk,temp_b3_4_1_r,temp_b3_4_1_i,temp_b3_4_9_r,temp_b3_4_9_i,temp_b3_12_1_r,temp_b3_12_1_i,temp_b3_12_9_r,temp_b3_12_9_i,temp_m4_4_1_r,temp_m4_4_1_i,temp_m4_4_9_r,temp_m4_4_9_i,temp_m4_12_1_r,temp_m4_12_1_i,temp_m4_12_9_r,temp_m4_12_9_i,`W0_real,`W0_imag,`W6_real,`W6_imag,`W6_real,`W6_imag);
butterfly butterfly793 (clk,temp_m4_4_1_r,temp_m4_4_1_i,temp_m4_4_9_r,temp_m4_4_9_i,temp_m4_12_1_r,temp_m4_12_1_i,temp_m4_12_9_r,temp_m4_12_9_i,temp_b4_4_1_r,temp_b4_4_1_i,temp_b4_4_9_r,temp_b4_4_9_i,temp_b4_12_1_r,temp_b4_12_1_i,temp_b4_12_9_r,temp_b4_12_9_i);
MULT MULT794 (clk,temp_b3_4_2_r,temp_b3_4_2_i,temp_b3_4_10_r,temp_b3_4_10_i,temp_b3_12_2_r,temp_b3_12_2_i,temp_b3_12_10_r,temp_b3_12_10_i,temp_m4_4_2_r,temp_m4_4_2_i,temp_m4_4_10_r,temp_m4_4_10_i,temp_m4_12_2_r,temp_m4_12_2_i,temp_m4_12_10_r,temp_m4_12_10_i,`W2_real,`W2_imag,`W6_real,`W6_imag,`W8_real,`W8_imag);
butterfly butterfly794 (clk,temp_m4_4_2_r,temp_m4_4_2_i,temp_m4_4_10_r,temp_m4_4_10_i,temp_m4_12_2_r,temp_m4_12_2_i,temp_m4_12_10_r,temp_m4_12_10_i,temp_b4_4_2_r,temp_b4_4_2_i,temp_b4_4_10_r,temp_b4_4_10_i,temp_b4_12_2_r,temp_b4_12_2_i,temp_b4_12_10_r,temp_b4_12_10_i);
MULT MULT795 (clk,temp_b3_4_3_r,temp_b3_4_3_i,temp_b3_4_11_r,temp_b3_4_11_i,temp_b3_12_3_r,temp_b3_12_3_i,temp_b3_12_11_r,temp_b3_12_11_i,temp_m4_4_3_r,temp_m4_4_3_i,temp_m4_4_11_r,temp_m4_4_11_i,temp_m4_12_3_r,temp_m4_12_3_i,temp_m4_12_11_r,temp_m4_12_11_i,`W4_real,`W4_imag,`W6_real,`W6_imag,`W10_real,`W10_imag);
butterfly butterfly795 (clk,temp_m4_4_3_r,temp_m4_4_3_i,temp_m4_4_11_r,temp_m4_4_11_i,temp_m4_12_3_r,temp_m4_12_3_i,temp_m4_12_11_r,temp_m4_12_11_i,temp_b4_4_3_r,temp_b4_4_3_i,temp_b4_4_11_r,temp_b4_4_11_i,temp_b4_12_3_r,temp_b4_12_3_i,temp_b4_12_11_r,temp_b4_12_11_i);
MULT MULT796 (clk,temp_b3_4_4_r,temp_b3_4_4_i,temp_b3_4_12_r,temp_b3_4_12_i,temp_b3_12_4_r,temp_b3_12_4_i,temp_b3_12_12_r,temp_b3_12_12_i,temp_m4_4_4_r,temp_m4_4_4_i,temp_m4_4_12_r,temp_m4_4_12_i,temp_m4_12_4_r,temp_m4_12_4_i,temp_m4_12_12_r,temp_m4_12_12_i,`W6_real,`W6_imag,`W6_real,`W6_imag,`W12_real,`W12_imag);
butterfly butterfly796 (clk,temp_m4_4_4_r,temp_m4_4_4_i,temp_m4_4_12_r,temp_m4_4_12_i,temp_m4_12_4_r,temp_m4_12_4_i,temp_m4_12_12_r,temp_m4_12_12_i,temp_b4_4_4_r,temp_b4_4_4_i,temp_b4_4_12_r,temp_b4_4_12_i,temp_b4_12_4_r,temp_b4_12_4_i,temp_b4_12_12_r,temp_b4_12_12_i);
MULT MULT797 (clk,temp_b3_4_5_r,temp_b3_4_5_i,temp_b3_4_13_r,temp_b3_4_13_i,temp_b3_12_5_r,temp_b3_12_5_i,temp_b3_12_13_r,temp_b3_12_13_i,temp_m4_4_5_r,temp_m4_4_5_i,temp_m4_4_13_r,temp_m4_4_13_i,temp_m4_12_5_r,temp_m4_12_5_i,temp_m4_12_13_r,temp_m4_12_13_i,`W8_real,`W8_imag,`W6_real,`W6_imag,`W14_real,`W14_imag);
butterfly butterfly797 (clk,temp_m4_4_5_r,temp_m4_4_5_i,temp_m4_4_13_r,temp_m4_4_13_i,temp_m4_12_5_r,temp_m4_12_5_i,temp_m4_12_13_r,temp_m4_12_13_i,temp_b4_4_5_r,temp_b4_4_5_i,temp_b4_4_13_r,temp_b4_4_13_i,temp_b4_12_5_r,temp_b4_12_5_i,temp_b4_12_13_r,temp_b4_12_13_i);
MULT MULT798 (clk,temp_b3_4_6_r,temp_b3_4_6_i,temp_b3_4_14_r,temp_b3_4_14_i,temp_b3_12_6_r,temp_b3_12_6_i,temp_b3_12_14_r,temp_b3_12_14_i,temp_m4_4_6_r,temp_m4_4_6_i,temp_m4_4_14_r,temp_m4_4_14_i,temp_m4_12_6_r,temp_m4_12_6_i,temp_m4_12_14_r,temp_m4_12_14_i,`W10_real,`W10_imag,`W6_real,`W6_imag,`W16_real,`W16_imag);
butterfly butterfly798 (clk,temp_m4_4_6_r,temp_m4_4_6_i,temp_m4_4_14_r,temp_m4_4_14_i,temp_m4_12_6_r,temp_m4_12_6_i,temp_m4_12_14_r,temp_m4_12_14_i,temp_b4_4_6_r,temp_b4_4_6_i,temp_b4_4_14_r,temp_b4_4_14_i,temp_b4_12_6_r,temp_b4_12_6_i,temp_b4_12_14_r,temp_b4_12_14_i);
MULT MULT799 (clk,temp_b3_4_7_r,temp_b3_4_7_i,temp_b3_4_15_r,temp_b3_4_15_i,temp_b3_12_7_r,temp_b3_12_7_i,temp_b3_12_15_r,temp_b3_12_15_i,temp_m4_4_7_r,temp_m4_4_7_i,temp_m4_4_15_r,temp_m4_4_15_i,temp_m4_12_7_r,temp_m4_12_7_i,temp_m4_12_15_r,temp_m4_12_15_i,`W12_real,`W12_imag,`W6_real,`W6_imag,`W18_real,`W18_imag);
butterfly butterfly799 (clk,temp_m4_4_7_r,temp_m4_4_7_i,temp_m4_4_15_r,temp_m4_4_15_i,temp_m4_12_7_r,temp_m4_12_7_i,temp_m4_12_15_r,temp_m4_12_15_i,temp_b4_4_7_r,temp_b4_4_7_i,temp_b4_4_15_r,temp_b4_4_15_i,temp_b4_12_7_r,temp_b4_12_7_i,temp_b4_12_15_r,temp_b4_12_15_i);
MULT MULT800 (clk,temp_b3_4_8_r,temp_b3_4_8_i,temp_b3_4_16_r,temp_b3_4_16_i,temp_b3_12_8_r,temp_b3_12_8_i,temp_b3_12_16_r,temp_b3_12_16_i,temp_m4_4_8_r,temp_m4_4_8_i,temp_m4_4_16_r,temp_m4_4_16_i,temp_m4_12_8_r,temp_m4_12_8_i,temp_m4_12_16_r,temp_m4_12_16_i,`W14_real,`W14_imag,`W6_real,`W6_imag,`W20_real,`W20_imag);
butterfly butterfly800 (clk,temp_m4_4_8_r,temp_m4_4_8_i,temp_m4_4_16_r,temp_m4_4_16_i,temp_m4_12_8_r,temp_m4_12_8_i,temp_m4_12_16_r,temp_m4_12_16_i,temp_b4_4_8_r,temp_b4_4_8_i,temp_b4_4_16_r,temp_b4_4_16_i,temp_b4_12_8_r,temp_b4_12_8_i,temp_b4_12_16_r,temp_b4_12_16_i);
MULT MULT801 (clk,temp_b3_5_1_r,temp_b3_5_1_i,temp_b3_5_9_r,temp_b3_5_9_i,temp_b3_13_1_r,temp_b3_13_1_i,temp_b3_13_9_r,temp_b3_13_9_i,temp_m4_5_1_r,temp_m4_5_1_i,temp_m4_5_9_r,temp_m4_5_9_i,temp_m4_13_1_r,temp_m4_13_1_i,temp_m4_13_9_r,temp_m4_13_9_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly801 (clk,temp_m4_5_1_r,temp_m4_5_1_i,temp_m4_5_9_r,temp_m4_5_9_i,temp_m4_13_1_r,temp_m4_13_1_i,temp_m4_13_9_r,temp_m4_13_9_i,temp_b4_5_1_r,temp_b4_5_1_i,temp_b4_5_9_r,temp_b4_5_9_i,temp_b4_13_1_r,temp_b4_13_1_i,temp_b4_13_9_r,temp_b4_13_9_i);
MULT MULT802 (clk,temp_b3_5_2_r,temp_b3_5_2_i,temp_b3_5_10_r,temp_b3_5_10_i,temp_b3_13_2_r,temp_b3_13_2_i,temp_b3_13_10_r,temp_b3_13_10_i,temp_m4_5_2_r,temp_m4_5_2_i,temp_m4_5_10_r,temp_m4_5_10_i,temp_m4_13_2_r,temp_m4_13_2_i,temp_m4_13_10_r,temp_m4_13_10_i,`W2_real,`W2_imag,`W8_real,`W8_imag,`W10_real,`W10_imag);
butterfly butterfly802 (clk,temp_m4_5_2_r,temp_m4_5_2_i,temp_m4_5_10_r,temp_m4_5_10_i,temp_m4_13_2_r,temp_m4_13_2_i,temp_m4_13_10_r,temp_m4_13_10_i,temp_b4_5_2_r,temp_b4_5_2_i,temp_b4_5_10_r,temp_b4_5_10_i,temp_b4_13_2_r,temp_b4_13_2_i,temp_b4_13_10_r,temp_b4_13_10_i);
MULT MULT803 (clk,temp_b3_5_3_r,temp_b3_5_3_i,temp_b3_5_11_r,temp_b3_5_11_i,temp_b3_13_3_r,temp_b3_13_3_i,temp_b3_13_11_r,temp_b3_13_11_i,temp_m4_5_3_r,temp_m4_5_3_i,temp_m4_5_11_r,temp_m4_5_11_i,temp_m4_13_3_r,temp_m4_13_3_i,temp_m4_13_11_r,temp_m4_13_11_i,`W4_real,`W4_imag,`W8_real,`W8_imag,`W12_real,`W12_imag);
butterfly butterfly803 (clk,temp_m4_5_3_r,temp_m4_5_3_i,temp_m4_5_11_r,temp_m4_5_11_i,temp_m4_13_3_r,temp_m4_13_3_i,temp_m4_13_11_r,temp_m4_13_11_i,temp_b4_5_3_r,temp_b4_5_3_i,temp_b4_5_11_r,temp_b4_5_11_i,temp_b4_13_3_r,temp_b4_13_3_i,temp_b4_13_11_r,temp_b4_13_11_i);
MULT MULT804 (clk,temp_b3_5_4_r,temp_b3_5_4_i,temp_b3_5_12_r,temp_b3_5_12_i,temp_b3_13_4_r,temp_b3_13_4_i,temp_b3_13_12_r,temp_b3_13_12_i,temp_m4_5_4_r,temp_m4_5_4_i,temp_m4_5_12_r,temp_m4_5_12_i,temp_m4_13_4_r,temp_m4_13_4_i,temp_m4_13_12_r,temp_m4_13_12_i,`W6_real,`W6_imag,`W8_real,`W8_imag,`W14_real,`W14_imag);
butterfly butterfly804 (clk,temp_m4_5_4_r,temp_m4_5_4_i,temp_m4_5_12_r,temp_m4_5_12_i,temp_m4_13_4_r,temp_m4_13_4_i,temp_m4_13_12_r,temp_m4_13_12_i,temp_b4_5_4_r,temp_b4_5_4_i,temp_b4_5_12_r,temp_b4_5_12_i,temp_b4_13_4_r,temp_b4_13_4_i,temp_b4_13_12_r,temp_b4_13_12_i);
MULT MULT805 (clk,temp_b3_5_5_r,temp_b3_5_5_i,temp_b3_5_13_r,temp_b3_5_13_i,temp_b3_13_5_r,temp_b3_13_5_i,temp_b3_13_13_r,temp_b3_13_13_i,temp_m4_5_5_r,temp_m4_5_5_i,temp_m4_5_13_r,temp_m4_5_13_i,temp_m4_13_5_r,temp_m4_13_5_i,temp_m4_13_13_r,temp_m4_13_13_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly805 (clk,temp_m4_5_5_r,temp_m4_5_5_i,temp_m4_5_13_r,temp_m4_5_13_i,temp_m4_13_5_r,temp_m4_13_5_i,temp_m4_13_13_r,temp_m4_13_13_i,temp_b4_5_5_r,temp_b4_5_5_i,temp_b4_5_13_r,temp_b4_5_13_i,temp_b4_13_5_r,temp_b4_13_5_i,temp_b4_13_13_r,temp_b4_13_13_i);
MULT MULT806 (clk,temp_b3_5_6_r,temp_b3_5_6_i,temp_b3_5_14_r,temp_b3_5_14_i,temp_b3_13_6_r,temp_b3_13_6_i,temp_b3_13_14_r,temp_b3_13_14_i,temp_m4_5_6_r,temp_m4_5_6_i,temp_m4_5_14_r,temp_m4_5_14_i,temp_m4_13_6_r,temp_m4_13_6_i,temp_m4_13_14_r,temp_m4_13_14_i,`W10_real,`W10_imag,`W8_real,`W8_imag,`W18_real,`W18_imag);
butterfly butterfly806 (clk,temp_m4_5_6_r,temp_m4_5_6_i,temp_m4_5_14_r,temp_m4_5_14_i,temp_m4_13_6_r,temp_m4_13_6_i,temp_m4_13_14_r,temp_m4_13_14_i,temp_b4_5_6_r,temp_b4_5_6_i,temp_b4_5_14_r,temp_b4_5_14_i,temp_b4_13_6_r,temp_b4_13_6_i,temp_b4_13_14_r,temp_b4_13_14_i);
MULT MULT807 (clk,temp_b3_5_7_r,temp_b3_5_7_i,temp_b3_5_15_r,temp_b3_5_15_i,temp_b3_13_7_r,temp_b3_13_7_i,temp_b3_13_15_r,temp_b3_13_15_i,temp_m4_5_7_r,temp_m4_5_7_i,temp_m4_5_15_r,temp_m4_5_15_i,temp_m4_13_7_r,temp_m4_13_7_i,temp_m4_13_15_r,temp_m4_13_15_i,`W12_real,`W12_imag,`W8_real,`W8_imag,`W20_real,`W20_imag);
butterfly butterfly807 (clk,temp_m4_5_7_r,temp_m4_5_7_i,temp_m4_5_15_r,temp_m4_5_15_i,temp_m4_13_7_r,temp_m4_13_7_i,temp_m4_13_15_r,temp_m4_13_15_i,temp_b4_5_7_r,temp_b4_5_7_i,temp_b4_5_15_r,temp_b4_5_15_i,temp_b4_13_7_r,temp_b4_13_7_i,temp_b4_13_15_r,temp_b4_13_15_i);
MULT MULT808 (clk,temp_b3_5_8_r,temp_b3_5_8_i,temp_b3_5_16_r,temp_b3_5_16_i,temp_b3_13_8_r,temp_b3_13_8_i,temp_b3_13_16_r,temp_b3_13_16_i,temp_m4_5_8_r,temp_m4_5_8_i,temp_m4_5_16_r,temp_m4_5_16_i,temp_m4_13_8_r,temp_m4_13_8_i,temp_m4_13_16_r,temp_m4_13_16_i,`W14_real,`W14_imag,`W8_real,`W8_imag,`W22_real,`W22_imag);
butterfly butterfly808 (clk,temp_m4_5_8_r,temp_m4_5_8_i,temp_m4_5_16_r,temp_m4_5_16_i,temp_m4_13_8_r,temp_m4_13_8_i,temp_m4_13_16_r,temp_m4_13_16_i,temp_b4_5_8_r,temp_b4_5_8_i,temp_b4_5_16_r,temp_b4_5_16_i,temp_b4_13_8_r,temp_b4_13_8_i,temp_b4_13_16_r,temp_b4_13_16_i);
MULT MULT809 (clk,temp_b3_6_1_r,temp_b3_6_1_i,temp_b3_6_9_r,temp_b3_6_9_i,temp_b3_14_1_r,temp_b3_14_1_i,temp_b3_14_9_r,temp_b3_14_9_i,temp_m4_6_1_r,temp_m4_6_1_i,temp_m4_6_9_r,temp_m4_6_9_i,temp_m4_14_1_r,temp_m4_14_1_i,temp_m4_14_9_r,temp_m4_14_9_i,`W0_real,`W0_imag,`W10_real,`W10_imag,`W10_real,`W10_imag);
butterfly butterfly809 (clk,temp_m4_6_1_r,temp_m4_6_1_i,temp_m4_6_9_r,temp_m4_6_9_i,temp_m4_14_1_r,temp_m4_14_1_i,temp_m4_14_9_r,temp_m4_14_9_i,temp_b4_6_1_r,temp_b4_6_1_i,temp_b4_6_9_r,temp_b4_6_9_i,temp_b4_14_1_r,temp_b4_14_1_i,temp_b4_14_9_r,temp_b4_14_9_i);
MULT MULT810 (clk,temp_b3_6_2_r,temp_b3_6_2_i,temp_b3_6_10_r,temp_b3_6_10_i,temp_b3_14_2_r,temp_b3_14_2_i,temp_b3_14_10_r,temp_b3_14_10_i,temp_m4_6_2_r,temp_m4_6_2_i,temp_m4_6_10_r,temp_m4_6_10_i,temp_m4_14_2_r,temp_m4_14_2_i,temp_m4_14_10_r,temp_m4_14_10_i,`W2_real,`W2_imag,`W10_real,`W10_imag,`W12_real,`W12_imag);
butterfly butterfly810 (clk,temp_m4_6_2_r,temp_m4_6_2_i,temp_m4_6_10_r,temp_m4_6_10_i,temp_m4_14_2_r,temp_m4_14_2_i,temp_m4_14_10_r,temp_m4_14_10_i,temp_b4_6_2_r,temp_b4_6_2_i,temp_b4_6_10_r,temp_b4_6_10_i,temp_b4_14_2_r,temp_b4_14_2_i,temp_b4_14_10_r,temp_b4_14_10_i);
MULT MULT811 (clk,temp_b3_6_3_r,temp_b3_6_3_i,temp_b3_6_11_r,temp_b3_6_11_i,temp_b3_14_3_r,temp_b3_14_3_i,temp_b3_14_11_r,temp_b3_14_11_i,temp_m4_6_3_r,temp_m4_6_3_i,temp_m4_6_11_r,temp_m4_6_11_i,temp_m4_14_3_r,temp_m4_14_3_i,temp_m4_14_11_r,temp_m4_14_11_i,`W4_real,`W4_imag,`W10_real,`W10_imag,`W14_real,`W14_imag);
butterfly butterfly811 (clk,temp_m4_6_3_r,temp_m4_6_3_i,temp_m4_6_11_r,temp_m4_6_11_i,temp_m4_14_3_r,temp_m4_14_3_i,temp_m4_14_11_r,temp_m4_14_11_i,temp_b4_6_3_r,temp_b4_6_3_i,temp_b4_6_11_r,temp_b4_6_11_i,temp_b4_14_3_r,temp_b4_14_3_i,temp_b4_14_11_r,temp_b4_14_11_i);
MULT MULT812 (clk,temp_b3_6_4_r,temp_b3_6_4_i,temp_b3_6_12_r,temp_b3_6_12_i,temp_b3_14_4_r,temp_b3_14_4_i,temp_b3_14_12_r,temp_b3_14_12_i,temp_m4_6_4_r,temp_m4_6_4_i,temp_m4_6_12_r,temp_m4_6_12_i,temp_m4_14_4_r,temp_m4_14_4_i,temp_m4_14_12_r,temp_m4_14_12_i,`W6_real,`W6_imag,`W10_real,`W10_imag,`W16_real,`W16_imag);
butterfly butterfly812 (clk,temp_m4_6_4_r,temp_m4_6_4_i,temp_m4_6_12_r,temp_m4_6_12_i,temp_m4_14_4_r,temp_m4_14_4_i,temp_m4_14_12_r,temp_m4_14_12_i,temp_b4_6_4_r,temp_b4_6_4_i,temp_b4_6_12_r,temp_b4_6_12_i,temp_b4_14_4_r,temp_b4_14_4_i,temp_b4_14_12_r,temp_b4_14_12_i);
MULT MULT813 (clk,temp_b3_6_5_r,temp_b3_6_5_i,temp_b3_6_13_r,temp_b3_6_13_i,temp_b3_14_5_r,temp_b3_14_5_i,temp_b3_14_13_r,temp_b3_14_13_i,temp_m4_6_5_r,temp_m4_6_5_i,temp_m4_6_13_r,temp_m4_6_13_i,temp_m4_14_5_r,temp_m4_14_5_i,temp_m4_14_13_r,temp_m4_14_13_i,`W8_real,`W8_imag,`W10_real,`W10_imag,`W18_real,`W18_imag);
butterfly butterfly813 (clk,temp_m4_6_5_r,temp_m4_6_5_i,temp_m4_6_13_r,temp_m4_6_13_i,temp_m4_14_5_r,temp_m4_14_5_i,temp_m4_14_13_r,temp_m4_14_13_i,temp_b4_6_5_r,temp_b4_6_5_i,temp_b4_6_13_r,temp_b4_6_13_i,temp_b4_14_5_r,temp_b4_14_5_i,temp_b4_14_13_r,temp_b4_14_13_i);
MULT MULT814 (clk,temp_b3_6_6_r,temp_b3_6_6_i,temp_b3_6_14_r,temp_b3_6_14_i,temp_b3_14_6_r,temp_b3_14_6_i,temp_b3_14_14_r,temp_b3_14_14_i,temp_m4_6_6_r,temp_m4_6_6_i,temp_m4_6_14_r,temp_m4_6_14_i,temp_m4_14_6_r,temp_m4_14_6_i,temp_m4_14_14_r,temp_m4_14_14_i,`W10_real,`W10_imag,`W10_real,`W10_imag,`W20_real,`W20_imag);
butterfly butterfly814 (clk,temp_m4_6_6_r,temp_m4_6_6_i,temp_m4_6_14_r,temp_m4_6_14_i,temp_m4_14_6_r,temp_m4_14_6_i,temp_m4_14_14_r,temp_m4_14_14_i,temp_b4_6_6_r,temp_b4_6_6_i,temp_b4_6_14_r,temp_b4_6_14_i,temp_b4_14_6_r,temp_b4_14_6_i,temp_b4_14_14_r,temp_b4_14_14_i);
MULT MULT815 (clk,temp_b3_6_7_r,temp_b3_6_7_i,temp_b3_6_15_r,temp_b3_6_15_i,temp_b3_14_7_r,temp_b3_14_7_i,temp_b3_14_15_r,temp_b3_14_15_i,temp_m4_6_7_r,temp_m4_6_7_i,temp_m4_6_15_r,temp_m4_6_15_i,temp_m4_14_7_r,temp_m4_14_7_i,temp_m4_14_15_r,temp_m4_14_15_i,`W12_real,`W12_imag,`W10_real,`W10_imag,`W22_real,`W22_imag);
butterfly butterfly815 (clk,temp_m4_6_7_r,temp_m4_6_7_i,temp_m4_6_15_r,temp_m4_6_15_i,temp_m4_14_7_r,temp_m4_14_7_i,temp_m4_14_15_r,temp_m4_14_15_i,temp_b4_6_7_r,temp_b4_6_7_i,temp_b4_6_15_r,temp_b4_6_15_i,temp_b4_14_7_r,temp_b4_14_7_i,temp_b4_14_15_r,temp_b4_14_15_i);
MULT MULT816 (clk,temp_b3_6_8_r,temp_b3_6_8_i,temp_b3_6_16_r,temp_b3_6_16_i,temp_b3_14_8_r,temp_b3_14_8_i,temp_b3_14_16_r,temp_b3_14_16_i,temp_m4_6_8_r,temp_m4_6_8_i,temp_m4_6_16_r,temp_m4_6_16_i,temp_m4_14_8_r,temp_m4_14_8_i,temp_m4_14_16_r,temp_m4_14_16_i,`W14_real,`W14_imag,`W10_real,`W10_imag,`W24_real,`W24_imag);
butterfly butterfly816 (clk,temp_m4_6_8_r,temp_m4_6_8_i,temp_m4_6_16_r,temp_m4_6_16_i,temp_m4_14_8_r,temp_m4_14_8_i,temp_m4_14_16_r,temp_m4_14_16_i,temp_b4_6_8_r,temp_b4_6_8_i,temp_b4_6_16_r,temp_b4_6_16_i,temp_b4_14_8_r,temp_b4_14_8_i,temp_b4_14_16_r,temp_b4_14_16_i);
MULT MULT817 (clk,temp_b3_7_1_r,temp_b3_7_1_i,temp_b3_7_9_r,temp_b3_7_9_i,temp_b3_15_1_r,temp_b3_15_1_i,temp_b3_15_9_r,temp_b3_15_9_i,temp_m4_7_1_r,temp_m4_7_1_i,temp_m4_7_9_r,temp_m4_7_9_i,temp_m4_15_1_r,temp_m4_15_1_i,temp_m4_15_9_r,temp_m4_15_9_i,`W0_real,`W0_imag,`W12_real,`W12_imag,`W12_real,`W12_imag);
butterfly butterfly817 (clk,temp_m4_7_1_r,temp_m4_7_1_i,temp_m4_7_9_r,temp_m4_7_9_i,temp_m4_15_1_r,temp_m4_15_1_i,temp_m4_15_9_r,temp_m4_15_9_i,temp_b4_7_1_r,temp_b4_7_1_i,temp_b4_7_9_r,temp_b4_7_9_i,temp_b4_15_1_r,temp_b4_15_1_i,temp_b4_15_9_r,temp_b4_15_9_i);
MULT MULT818 (clk,temp_b3_7_2_r,temp_b3_7_2_i,temp_b3_7_10_r,temp_b3_7_10_i,temp_b3_15_2_r,temp_b3_15_2_i,temp_b3_15_10_r,temp_b3_15_10_i,temp_m4_7_2_r,temp_m4_7_2_i,temp_m4_7_10_r,temp_m4_7_10_i,temp_m4_15_2_r,temp_m4_15_2_i,temp_m4_15_10_r,temp_m4_15_10_i,`W2_real,`W2_imag,`W12_real,`W12_imag,`W14_real,`W14_imag);
butterfly butterfly818 (clk,temp_m4_7_2_r,temp_m4_7_2_i,temp_m4_7_10_r,temp_m4_7_10_i,temp_m4_15_2_r,temp_m4_15_2_i,temp_m4_15_10_r,temp_m4_15_10_i,temp_b4_7_2_r,temp_b4_7_2_i,temp_b4_7_10_r,temp_b4_7_10_i,temp_b4_15_2_r,temp_b4_15_2_i,temp_b4_15_10_r,temp_b4_15_10_i);
MULT MULT819 (clk,temp_b3_7_3_r,temp_b3_7_3_i,temp_b3_7_11_r,temp_b3_7_11_i,temp_b3_15_3_r,temp_b3_15_3_i,temp_b3_15_11_r,temp_b3_15_11_i,temp_m4_7_3_r,temp_m4_7_3_i,temp_m4_7_11_r,temp_m4_7_11_i,temp_m4_15_3_r,temp_m4_15_3_i,temp_m4_15_11_r,temp_m4_15_11_i,`W4_real,`W4_imag,`W12_real,`W12_imag,`W16_real,`W16_imag);
butterfly butterfly819 (clk,temp_m4_7_3_r,temp_m4_7_3_i,temp_m4_7_11_r,temp_m4_7_11_i,temp_m4_15_3_r,temp_m4_15_3_i,temp_m4_15_11_r,temp_m4_15_11_i,temp_b4_7_3_r,temp_b4_7_3_i,temp_b4_7_11_r,temp_b4_7_11_i,temp_b4_15_3_r,temp_b4_15_3_i,temp_b4_15_11_r,temp_b4_15_11_i);
MULT MULT820 (clk,temp_b3_7_4_r,temp_b3_7_4_i,temp_b3_7_12_r,temp_b3_7_12_i,temp_b3_15_4_r,temp_b3_15_4_i,temp_b3_15_12_r,temp_b3_15_12_i,temp_m4_7_4_r,temp_m4_7_4_i,temp_m4_7_12_r,temp_m4_7_12_i,temp_m4_15_4_r,temp_m4_15_4_i,temp_m4_15_12_r,temp_m4_15_12_i,`W6_real,`W6_imag,`W12_real,`W12_imag,`W18_real,`W18_imag);
butterfly butterfly820 (clk,temp_m4_7_4_r,temp_m4_7_4_i,temp_m4_7_12_r,temp_m4_7_12_i,temp_m4_15_4_r,temp_m4_15_4_i,temp_m4_15_12_r,temp_m4_15_12_i,temp_b4_7_4_r,temp_b4_7_4_i,temp_b4_7_12_r,temp_b4_7_12_i,temp_b4_15_4_r,temp_b4_15_4_i,temp_b4_15_12_r,temp_b4_15_12_i);
MULT MULT821 (clk,temp_b3_7_5_r,temp_b3_7_5_i,temp_b3_7_13_r,temp_b3_7_13_i,temp_b3_15_5_r,temp_b3_15_5_i,temp_b3_15_13_r,temp_b3_15_13_i,temp_m4_7_5_r,temp_m4_7_5_i,temp_m4_7_13_r,temp_m4_7_13_i,temp_m4_15_5_r,temp_m4_15_5_i,temp_m4_15_13_r,temp_m4_15_13_i,`W8_real,`W8_imag,`W12_real,`W12_imag,`W20_real,`W20_imag);
butterfly butterfly821 (clk,temp_m4_7_5_r,temp_m4_7_5_i,temp_m4_7_13_r,temp_m4_7_13_i,temp_m4_15_5_r,temp_m4_15_5_i,temp_m4_15_13_r,temp_m4_15_13_i,temp_b4_7_5_r,temp_b4_7_5_i,temp_b4_7_13_r,temp_b4_7_13_i,temp_b4_15_5_r,temp_b4_15_5_i,temp_b4_15_13_r,temp_b4_15_13_i);
MULT MULT822 (clk,temp_b3_7_6_r,temp_b3_7_6_i,temp_b3_7_14_r,temp_b3_7_14_i,temp_b3_15_6_r,temp_b3_15_6_i,temp_b3_15_14_r,temp_b3_15_14_i,temp_m4_7_6_r,temp_m4_7_6_i,temp_m4_7_14_r,temp_m4_7_14_i,temp_m4_15_6_r,temp_m4_15_6_i,temp_m4_15_14_r,temp_m4_15_14_i,`W10_real,`W10_imag,`W12_real,`W12_imag,`W22_real,`W22_imag);
butterfly butterfly822 (clk,temp_m4_7_6_r,temp_m4_7_6_i,temp_m4_7_14_r,temp_m4_7_14_i,temp_m4_15_6_r,temp_m4_15_6_i,temp_m4_15_14_r,temp_m4_15_14_i,temp_b4_7_6_r,temp_b4_7_6_i,temp_b4_7_14_r,temp_b4_7_14_i,temp_b4_15_6_r,temp_b4_15_6_i,temp_b4_15_14_r,temp_b4_15_14_i);
MULT MULT823 (clk,temp_b3_7_7_r,temp_b3_7_7_i,temp_b3_7_15_r,temp_b3_7_15_i,temp_b3_15_7_r,temp_b3_15_7_i,temp_b3_15_15_r,temp_b3_15_15_i,temp_m4_7_7_r,temp_m4_7_7_i,temp_m4_7_15_r,temp_m4_7_15_i,temp_m4_15_7_r,temp_m4_15_7_i,temp_m4_15_15_r,temp_m4_15_15_i,`W12_real,`W12_imag,`W12_real,`W12_imag,`W24_real,`W24_imag);
butterfly butterfly823 (clk,temp_m4_7_7_r,temp_m4_7_7_i,temp_m4_7_15_r,temp_m4_7_15_i,temp_m4_15_7_r,temp_m4_15_7_i,temp_m4_15_15_r,temp_m4_15_15_i,temp_b4_7_7_r,temp_b4_7_7_i,temp_b4_7_15_r,temp_b4_7_15_i,temp_b4_15_7_r,temp_b4_15_7_i,temp_b4_15_15_r,temp_b4_15_15_i);
MULT MULT824 (clk,temp_b3_7_8_r,temp_b3_7_8_i,temp_b3_7_16_r,temp_b3_7_16_i,temp_b3_15_8_r,temp_b3_15_8_i,temp_b3_15_16_r,temp_b3_15_16_i,temp_m4_7_8_r,temp_m4_7_8_i,temp_m4_7_16_r,temp_m4_7_16_i,temp_m4_15_8_r,temp_m4_15_8_i,temp_m4_15_16_r,temp_m4_15_16_i,`W14_real,`W14_imag,`W12_real,`W12_imag,`W26_real,`W26_imag);
butterfly butterfly824 (clk,temp_m4_7_8_r,temp_m4_7_8_i,temp_m4_7_16_r,temp_m4_7_16_i,temp_m4_15_8_r,temp_m4_15_8_i,temp_m4_15_16_r,temp_m4_15_16_i,temp_b4_7_8_r,temp_b4_7_8_i,temp_b4_7_16_r,temp_b4_7_16_i,temp_b4_15_8_r,temp_b4_15_8_i,temp_b4_15_16_r,temp_b4_15_16_i);
MULT MULT825 (clk,temp_b3_8_1_r,temp_b3_8_1_i,temp_b3_8_9_r,temp_b3_8_9_i,temp_b3_16_1_r,temp_b3_16_1_i,temp_b3_16_9_r,temp_b3_16_9_i,temp_m4_8_1_r,temp_m4_8_1_i,temp_m4_8_9_r,temp_m4_8_9_i,temp_m4_16_1_r,temp_m4_16_1_i,temp_m4_16_9_r,temp_m4_16_9_i,`W0_real,`W0_imag,`W14_real,`W14_imag,`W14_real,`W14_imag);
butterfly butterfly825 (clk,temp_m4_8_1_r,temp_m4_8_1_i,temp_m4_8_9_r,temp_m4_8_9_i,temp_m4_16_1_r,temp_m4_16_1_i,temp_m4_16_9_r,temp_m4_16_9_i,temp_b4_8_1_r,temp_b4_8_1_i,temp_b4_8_9_r,temp_b4_8_9_i,temp_b4_16_1_r,temp_b4_16_1_i,temp_b4_16_9_r,temp_b4_16_9_i);
MULT MULT826 (clk,temp_b3_8_2_r,temp_b3_8_2_i,temp_b3_8_10_r,temp_b3_8_10_i,temp_b3_16_2_r,temp_b3_16_2_i,temp_b3_16_10_r,temp_b3_16_10_i,temp_m4_8_2_r,temp_m4_8_2_i,temp_m4_8_10_r,temp_m4_8_10_i,temp_m4_16_2_r,temp_m4_16_2_i,temp_m4_16_10_r,temp_m4_16_10_i,`W2_real,`W2_imag,`W14_real,`W14_imag,`W16_real,`W16_imag);
butterfly butterfly826 (clk,temp_m4_8_2_r,temp_m4_8_2_i,temp_m4_8_10_r,temp_m4_8_10_i,temp_m4_16_2_r,temp_m4_16_2_i,temp_m4_16_10_r,temp_m4_16_10_i,temp_b4_8_2_r,temp_b4_8_2_i,temp_b4_8_10_r,temp_b4_8_10_i,temp_b4_16_2_r,temp_b4_16_2_i,temp_b4_16_10_r,temp_b4_16_10_i);
MULT MULT827 (clk,temp_b3_8_3_r,temp_b3_8_3_i,temp_b3_8_11_r,temp_b3_8_11_i,temp_b3_16_3_r,temp_b3_16_3_i,temp_b3_16_11_r,temp_b3_16_11_i,temp_m4_8_3_r,temp_m4_8_3_i,temp_m4_8_11_r,temp_m4_8_11_i,temp_m4_16_3_r,temp_m4_16_3_i,temp_m4_16_11_r,temp_m4_16_11_i,`W4_real,`W4_imag,`W14_real,`W14_imag,`W18_real,`W18_imag);
butterfly butterfly827 (clk,temp_m4_8_3_r,temp_m4_8_3_i,temp_m4_8_11_r,temp_m4_8_11_i,temp_m4_16_3_r,temp_m4_16_3_i,temp_m4_16_11_r,temp_m4_16_11_i,temp_b4_8_3_r,temp_b4_8_3_i,temp_b4_8_11_r,temp_b4_8_11_i,temp_b4_16_3_r,temp_b4_16_3_i,temp_b4_16_11_r,temp_b4_16_11_i);
MULT MULT828 (clk,temp_b3_8_4_r,temp_b3_8_4_i,temp_b3_8_12_r,temp_b3_8_12_i,temp_b3_16_4_r,temp_b3_16_4_i,temp_b3_16_12_r,temp_b3_16_12_i,temp_m4_8_4_r,temp_m4_8_4_i,temp_m4_8_12_r,temp_m4_8_12_i,temp_m4_16_4_r,temp_m4_16_4_i,temp_m4_16_12_r,temp_m4_16_12_i,`W6_real,`W6_imag,`W14_real,`W14_imag,`W20_real,`W20_imag);
butterfly butterfly828 (clk,temp_m4_8_4_r,temp_m4_8_4_i,temp_m4_8_12_r,temp_m4_8_12_i,temp_m4_16_4_r,temp_m4_16_4_i,temp_m4_16_12_r,temp_m4_16_12_i,temp_b4_8_4_r,temp_b4_8_4_i,temp_b4_8_12_r,temp_b4_8_12_i,temp_b4_16_4_r,temp_b4_16_4_i,temp_b4_16_12_r,temp_b4_16_12_i);
MULT MULT829 (clk,temp_b3_8_5_r,temp_b3_8_5_i,temp_b3_8_13_r,temp_b3_8_13_i,temp_b3_16_5_r,temp_b3_16_5_i,temp_b3_16_13_r,temp_b3_16_13_i,temp_m4_8_5_r,temp_m4_8_5_i,temp_m4_8_13_r,temp_m4_8_13_i,temp_m4_16_5_r,temp_m4_16_5_i,temp_m4_16_13_r,temp_m4_16_13_i,`W8_real,`W8_imag,`W14_real,`W14_imag,`W22_real,`W22_imag);
butterfly butterfly829 (clk,temp_m4_8_5_r,temp_m4_8_5_i,temp_m4_8_13_r,temp_m4_8_13_i,temp_m4_16_5_r,temp_m4_16_5_i,temp_m4_16_13_r,temp_m4_16_13_i,temp_b4_8_5_r,temp_b4_8_5_i,temp_b4_8_13_r,temp_b4_8_13_i,temp_b4_16_5_r,temp_b4_16_5_i,temp_b4_16_13_r,temp_b4_16_13_i);
MULT MULT830 (clk,temp_b3_8_6_r,temp_b3_8_6_i,temp_b3_8_14_r,temp_b3_8_14_i,temp_b3_16_6_r,temp_b3_16_6_i,temp_b3_16_14_r,temp_b3_16_14_i,temp_m4_8_6_r,temp_m4_8_6_i,temp_m4_8_14_r,temp_m4_8_14_i,temp_m4_16_6_r,temp_m4_16_6_i,temp_m4_16_14_r,temp_m4_16_14_i,`W10_real,`W10_imag,`W14_real,`W14_imag,`W24_real,`W24_imag);
butterfly butterfly830 (clk,temp_m4_8_6_r,temp_m4_8_6_i,temp_m4_8_14_r,temp_m4_8_14_i,temp_m4_16_6_r,temp_m4_16_6_i,temp_m4_16_14_r,temp_m4_16_14_i,temp_b4_8_6_r,temp_b4_8_6_i,temp_b4_8_14_r,temp_b4_8_14_i,temp_b4_16_6_r,temp_b4_16_6_i,temp_b4_16_14_r,temp_b4_16_14_i);
MULT MULT831 (clk,temp_b3_8_7_r,temp_b3_8_7_i,temp_b3_8_15_r,temp_b3_8_15_i,temp_b3_16_7_r,temp_b3_16_7_i,temp_b3_16_15_r,temp_b3_16_15_i,temp_m4_8_7_r,temp_m4_8_7_i,temp_m4_8_15_r,temp_m4_8_15_i,temp_m4_16_7_r,temp_m4_16_7_i,temp_m4_16_15_r,temp_m4_16_15_i,`W12_real,`W12_imag,`W14_real,`W14_imag,`W26_real,`W26_imag);
butterfly butterfly831 (clk,temp_m4_8_7_r,temp_m4_8_7_i,temp_m4_8_15_r,temp_m4_8_15_i,temp_m4_16_7_r,temp_m4_16_7_i,temp_m4_16_15_r,temp_m4_16_15_i,temp_b4_8_7_r,temp_b4_8_7_i,temp_b4_8_15_r,temp_b4_8_15_i,temp_b4_16_7_r,temp_b4_16_7_i,temp_b4_16_15_r,temp_b4_16_15_i);
MULT MULT832 (clk,temp_b3_8_8_r,temp_b3_8_8_i,temp_b3_8_16_r,temp_b3_8_16_i,temp_b3_16_8_r,temp_b3_16_8_i,temp_b3_16_16_r,temp_b3_16_16_i,temp_m4_8_8_r,temp_m4_8_8_i,temp_m4_8_16_r,temp_m4_8_16_i,temp_m4_16_8_r,temp_m4_16_8_i,temp_m4_16_16_r,temp_m4_16_16_i,`W14_real,`W14_imag,`W14_real,`W14_imag,`W28_real,`W28_imag);
butterfly butterfly832 (clk,temp_m4_8_8_r,temp_m4_8_8_i,temp_m4_8_16_r,temp_m4_8_16_i,temp_m4_16_8_r,temp_m4_16_8_i,temp_m4_16_16_r,temp_m4_16_16_i,temp_b4_8_8_r,temp_b4_8_8_i,temp_b4_8_16_r,temp_b4_8_16_i,temp_b4_16_8_r,temp_b4_16_8_i,temp_b4_16_16_r,temp_b4_16_16_i);
MULT MULT833 (clk,temp_b3_1_17_r,temp_b3_1_17_i,temp_b3_1_25_r,temp_b3_1_25_i,temp_b3_9_17_r,temp_b3_9_17_i,temp_b3_9_25_r,temp_b3_9_25_i,temp_m4_1_17_r,temp_m4_1_17_i,temp_m4_1_25_r,temp_m4_1_25_i,temp_m4_9_17_r,temp_m4_9_17_i,temp_m4_9_25_r,temp_m4_9_25_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly833 (clk,temp_m4_1_17_r,temp_m4_1_17_i,temp_m4_1_25_r,temp_m4_1_25_i,temp_m4_9_17_r,temp_m4_9_17_i,temp_m4_9_25_r,temp_m4_9_25_i,temp_b4_1_17_r,temp_b4_1_17_i,temp_b4_1_25_r,temp_b4_1_25_i,temp_b4_9_17_r,temp_b4_9_17_i,temp_b4_9_25_r,temp_b4_9_25_i);
MULT MULT834 (clk,temp_b3_1_18_r,temp_b3_1_18_i,temp_b3_1_26_r,temp_b3_1_26_i,temp_b3_9_18_r,temp_b3_9_18_i,temp_b3_9_26_r,temp_b3_9_26_i,temp_m4_1_18_r,temp_m4_1_18_i,temp_m4_1_26_r,temp_m4_1_26_i,temp_m4_9_18_r,temp_m4_9_18_i,temp_m4_9_26_r,temp_m4_9_26_i,`W2_real,`W2_imag,`W0_real,`W0_imag,`W2_real,`W2_imag);
butterfly butterfly834 (clk,temp_m4_1_18_r,temp_m4_1_18_i,temp_m4_1_26_r,temp_m4_1_26_i,temp_m4_9_18_r,temp_m4_9_18_i,temp_m4_9_26_r,temp_m4_9_26_i,temp_b4_1_18_r,temp_b4_1_18_i,temp_b4_1_26_r,temp_b4_1_26_i,temp_b4_9_18_r,temp_b4_9_18_i,temp_b4_9_26_r,temp_b4_9_26_i);
MULT MULT835 (clk,temp_b3_1_19_r,temp_b3_1_19_i,temp_b3_1_27_r,temp_b3_1_27_i,temp_b3_9_19_r,temp_b3_9_19_i,temp_b3_9_27_r,temp_b3_9_27_i,temp_m4_1_19_r,temp_m4_1_19_i,temp_m4_1_27_r,temp_m4_1_27_i,temp_m4_9_19_r,temp_m4_9_19_i,temp_m4_9_27_r,temp_m4_9_27_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly835 (clk,temp_m4_1_19_r,temp_m4_1_19_i,temp_m4_1_27_r,temp_m4_1_27_i,temp_m4_9_19_r,temp_m4_9_19_i,temp_m4_9_27_r,temp_m4_9_27_i,temp_b4_1_19_r,temp_b4_1_19_i,temp_b4_1_27_r,temp_b4_1_27_i,temp_b4_9_19_r,temp_b4_9_19_i,temp_b4_9_27_r,temp_b4_9_27_i);
MULT MULT836 (clk,temp_b3_1_20_r,temp_b3_1_20_i,temp_b3_1_28_r,temp_b3_1_28_i,temp_b3_9_20_r,temp_b3_9_20_i,temp_b3_9_28_r,temp_b3_9_28_i,temp_m4_1_20_r,temp_m4_1_20_i,temp_m4_1_28_r,temp_m4_1_28_i,temp_m4_9_20_r,temp_m4_9_20_i,temp_m4_9_28_r,temp_m4_9_28_i,`W6_real,`W6_imag,`W0_real,`W0_imag,`W6_real,`W6_imag);
butterfly butterfly836 (clk,temp_m4_1_20_r,temp_m4_1_20_i,temp_m4_1_28_r,temp_m4_1_28_i,temp_m4_9_20_r,temp_m4_9_20_i,temp_m4_9_28_r,temp_m4_9_28_i,temp_b4_1_20_r,temp_b4_1_20_i,temp_b4_1_28_r,temp_b4_1_28_i,temp_b4_9_20_r,temp_b4_9_20_i,temp_b4_9_28_r,temp_b4_9_28_i);
MULT MULT837 (clk,temp_b3_1_21_r,temp_b3_1_21_i,temp_b3_1_29_r,temp_b3_1_29_i,temp_b3_9_21_r,temp_b3_9_21_i,temp_b3_9_29_r,temp_b3_9_29_i,temp_m4_1_21_r,temp_m4_1_21_i,temp_m4_1_29_r,temp_m4_1_29_i,temp_m4_9_21_r,temp_m4_9_21_i,temp_m4_9_29_r,temp_m4_9_29_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly837 (clk,temp_m4_1_21_r,temp_m4_1_21_i,temp_m4_1_29_r,temp_m4_1_29_i,temp_m4_9_21_r,temp_m4_9_21_i,temp_m4_9_29_r,temp_m4_9_29_i,temp_b4_1_21_r,temp_b4_1_21_i,temp_b4_1_29_r,temp_b4_1_29_i,temp_b4_9_21_r,temp_b4_9_21_i,temp_b4_9_29_r,temp_b4_9_29_i);
MULT MULT838 (clk,temp_b3_1_22_r,temp_b3_1_22_i,temp_b3_1_30_r,temp_b3_1_30_i,temp_b3_9_22_r,temp_b3_9_22_i,temp_b3_9_30_r,temp_b3_9_30_i,temp_m4_1_22_r,temp_m4_1_22_i,temp_m4_1_30_r,temp_m4_1_30_i,temp_m4_9_22_r,temp_m4_9_22_i,temp_m4_9_30_r,temp_m4_9_30_i,`W10_real,`W10_imag,`W0_real,`W0_imag,`W10_real,`W10_imag);
butterfly butterfly838 (clk,temp_m4_1_22_r,temp_m4_1_22_i,temp_m4_1_30_r,temp_m4_1_30_i,temp_m4_9_22_r,temp_m4_9_22_i,temp_m4_9_30_r,temp_m4_9_30_i,temp_b4_1_22_r,temp_b4_1_22_i,temp_b4_1_30_r,temp_b4_1_30_i,temp_b4_9_22_r,temp_b4_9_22_i,temp_b4_9_30_r,temp_b4_9_30_i);
MULT MULT839 (clk,temp_b3_1_23_r,temp_b3_1_23_i,temp_b3_1_31_r,temp_b3_1_31_i,temp_b3_9_23_r,temp_b3_9_23_i,temp_b3_9_31_r,temp_b3_9_31_i,temp_m4_1_23_r,temp_m4_1_23_i,temp_m4_1_31_r,temp_m4_1_31_i,temp_m4_9_23_r,temp_m4_9_23_i,temp_m4_9_31_r,temp_m4_9_31_i,`W12_real,`W12_imag,`W0_real,`W0_imag,`W12_real,`W12_imag);
butterfly butterfly839 (clk,temp_m4_1_23_r,temp_m4_1_23_i,temp_m4_1_31_r,temp_m4_1_31_i,temp_m4_9_23_r,temp_m4_9_23_i,temp_m4_9_31_r,temp_m4_9_31_i,temp_b4_1_23_r,temp_b4_1_23_i,temp_b4_1_31_r,temp_b4_1_31_i,temp_b4_9_23_r,temp_b4_9_23_i,temp_b4_9_31_r,temp_b4_9_31_i);
MULT MULT840 (clk,temp_b3_1_24_r,temp_b3_1_24_i,temp_b3_1_32_r,temp_b3_1_32_i,temp_b3_9_24_r,temp_b3_9_24_i,temp_b3_9_32_r,temp_b3_9_32_i,temp_m4_1_24_r,temp_m4_1_24_i,temp_m4_1_32_r,temp_m4_1_32_i,temp_m4_9_24_r,temp_m4_9_24_i,temp_m4_9_32_r,temp_m4_9_32_i,`W14_real,`W14_imag,`W0_real,`W0_imag,`W14_real,`W14_imag);
butterfly butterfly840 (clk,temp_m4_1_24_r,temp_m4_1_24_i,temp_m4_1_32_r,temp_m4_1_32_i,temp_m4_9_24_r,temp_m4_9_24_i,temp_m4_9_32_r,temp_m4_9_32_i,temp_b4_1_24_r,temp_b4_1_24_i,temp_b4_1_32_r,temp_b4_1_32_i,temp_b4_9_24_r,temp_b4_9_24_i,temp_b4_9_32_r,temp_b4_9_32_i);
MULT MULT841 (clk,temp_b3_2_17_r,temp_b3_2_17_i,temp_b3_2_25_r,temp_b3_2_25_i,temp_b3_10_17_r,temp_b3_10_17_i,temp_b3_10_25_r,temp_b3_10_25_i,temp_m4_2_17_r,temp_m4_2_17_i,temp_m4_2_25_r,temp_m4_2_25_i,temp_m4_10_17_r,temp_m4_10_17_i,temp_m4_10_25_r,temp_m4_10_25_i,`W0_real,`W0_imag,`W2_real,`W2_imag,`W2_real,`W2_imag);
butterfly butterfly841 (clk,temp_m4_2_17_r,temp_m4_2_17_i,temp_m4_2_25_r,temp_m4_2_25_i,temp_m4_10_17_r,temp_m4_10_17_i,temp_m4_10_25_r,temp_m4_10_25_i,temp_b4_2_17_r,temp_b4_2_17_i,temp_b4_2_25_r,temp_b4_2_25_i,temp_b4_10_17_r,temp_b4_10_17_i,temp_b4_10_25_r,temp_b4_10_25_i);
MULT MULT842 (clk,temp_b3_2_18_r,temp_b3_2_18_i,temp_b3_2_26_r,temp_b3_2_26_i,temp_b3_10_18_r,temp_b3_10_18_i,temp_b3_10_26_r,temp_b3_10_26_i,temp_m4_2_18_r,temp_m4_2_18_i,temp_m4_2_26_r,temp_m4_2_26_i,temp_m4_10_18_r,temp_m4_10_18_i,temp_m4_10_26_r,temp_m4_10_26_i,`W2_real,`W2_imag,`W2_real,`W2_imag,`W4_real,`W4_imag);
butterfly butterfly842 (clk,temp_m4_2_18_r,temp_m4_2_18_i,temp_m4_2_26_r,temp_m4_2_26_i,temp_m4_10_18_r,temp_m4_10_18_i,temp_m4_10_26_r,temp_m4_10_26_i,temp_b4_2_18_r,temp_b4_2_18_i,temp_b4_2_26_r,temp_b4_2_26_i,temp_b4_10_18_r,temp_b4_10_18_i,temp_b4_10_26_r,temp_b4_10_26_i);
MULT MULT843 (clk,temp_b3_2_19_r,temp_b3_2_19_i,temp_b3_2_27_r,temp_b3_2_27_i,temp_b3_10_19_r,temp_b3_10_19_i,temp_b3_10_27_r,temp_b3_10_27_i,temp_m4_2_19_r,temp_m4_2_19_i,temp_m4_2_27_r,temp_m4_2_27_i,temp_m4_10_19_r,temp_m4_10_19_i,temp_m4_10_27_r,temp_m4_10_27_i,`W4_real,`W4_imag,`W2_real,`W2_imag,`W6_real,`W6_imag);
butterfly butterfly843 (clk,temp_m4_2_19_r,temp_m4_2_19_i,temp_m4_2_27_r,temp_m4_2_27_i,temp_m4_10_19_r,temp_m4_10_19_i,temp_m4_10_27_r,temp_m4_10_27_i,temp_b4_2_19_r,temp_b4_2_19_i,temp_b4_2_27_r,temp_b4_2_27_i,temp_b4_10_19_r,temp_b4_10_19_i,temp_b4_10_27_r,temp_b4_10_27_i);
MULT MULT844 (clk,temp_b3_2_20_r,temp_b3_2_20_i,temp_b3_2_28_r,temp_b3_2_28_i,temp_b3_10_20_r,temp_b3_10_20_i,temp_b3_10_28_r,temp_b3_10_28_i,temp_m4_2_20_r,temp_m4_2_20_i,temp_m4_2_28_r,temp_m4_2_28_i,temp_m4_10_20_r,temp_m4_10_20_i,temp_m4_10_28_r,temp_m4_10_28_i,`W6_real,`W6_imag,`W2_real,`W2_imag,`W8_real,`W8_imag);
butterfly butterfly844 (clk,temp_m4_2_20_r,temp_m4_2_20_i,temp_m4_2_28_r,temp_m4_2_28_i,temp_m4_10_20_r,temp_m4_10_20_i,temp_m4_10_28_r,temp_m4_10_28_i,temp_b4_2_20_r,temp_b4_2_20_i,temp_b4_2_28_r,temp_b4_2_28_i,temp_b4_10_20_r,temp_b4_10_20_i,temp_b4_10_28_r,temp_b4_10_28_i);
MULT MULT845 (clk,temp_b3_2_21_r,temp_b3_2_21_i,temp_b3_2_29_r,temp_b3_2_29_i,temp_b3_10_21_r,temp_b3_10_21_i,temp_b3_10_29_r,temp_b3_10_29_i,temp_m4_2_21_r,temp_m4_2_21_i,temp_m4_2_29_r,temp_m4_2_29_i,temp_m4_10_21_r,temp_m4_10_21_i,temp_m4_10_29_r,temp_m4_10_29_i,`W8_real,`W8_imag,`W2_real,`W2_imag,`W10_real,`W10_imag);
butterfly butterfly845 (clk,temp_m4_2_21_r,temp_m4_2_21_i,temp_m4_2_29_r,temp_m4_2_29_i,temp_m4_10_21_r,temp_m4_10_21_i,temp_m4_10_29_r,temp_m4_10_29_i,temp_b4_2_21_r,temp_b4_2_21_i,temp_b4_2_29_r,temp_b4_2_29_i,temp_b4_10_21_r,temp_b4_10_21_i,temp_b4_10_29_r,temp_b4_10_29_i);
MULT MULT846 (clk,temp_b3_2_22_r,temp_b3_2_22_i,temp_b3_2_30_r,temp_b3_2_30_i,temp_b3_10_22_r,temp_b3_10_22_i,temp_b3_10_30_r,temp_b3_10_30_i,temp_m4_2_22_r,temp_m4_2_22_i,temp_m4_2_30_r,temp_m4_2_30_i,temp_m4_10_22_r,temp_m4_10_22_i,temp_m4_10_30_r,temp_m4_10_30_i,`W10_real,`W10_imag,`W2_real,`W2_imag,`W12_real,`W12_imag);
butterfly butterfly846 (clk,temp_m4_2_22_r,temp_m4_2_22_i,temp_m4_2_30_r,temp_m4_2_30_i,temp_m4_10_22_r,temp_m4_10_22_i,temp_m4_10_30_r,temp_m4_10_30_i,temp_b4_2_22_r,temp_b4_2_22_i,temp_b4_2_30_r,temp_b4_2_30_i,temp_b4_10_22_r,temp_b4_10_22_i,temp_b4_10_30_r,temp_b4_10_30_i);
MULT MULT847 (clk,temp_b3_2_23_r,temp_b3_2_23_i,temp_b3_2_31_r,temp_b3_2_31_i,temp_b3_10_23_r,temp_b3_10_23_i,temp_b3_10_31_r,temp_b3_10_31_i,temp_m4_2_23_r,temp_m4_2_23_i,temp_m4_2_31_r,temp_m4_2_31_i,temp_m4_10_23_r,temp_m4_10_23_i,temp_m4_10_31_r,temp_m4_10_31_i,`W12_real,`W12_imag,`W2_real,`W2_imag,`W14_real,`W14_imag);
butterfly butterfly847 (clk,temp_m4_2_23_r,temp_m4_2_23_i,temp_m4_2_31_r,temp_m4_2_31_i,temp_m4_10_23_r,temp_m4_10_23_i,temp_m4_10_31_r,temp_m4_10_31_i,temp_b4_2_23_r,temp_b4_2_23_i,temp_b4_2_31_r,temp_b4_2_31_i,temp_b4_10_23_r,temp_b4_10_23_i,temp_b4_10_31_r,temp_b4_10_31_i);
MULT MULT848 (clk,temp_b3_2_24_r,temp_b3_2_24_i,temp_b3_2_32_r,temp_b3_2_32_i,temp_b3_10_24_r,temp_b3_10_24_i,temp_b3_10_32_r,temp_b3_10_32_i,temp_m4_2_24_r,temp_m4_2_24_i,temp_m4_2_32_r,temp_m4_2_32_i,temp_m4_10_24_r,temp_m4_10_24_i,temp_m4_10_32_r,temp_m4_10_32_i,`W14_real,`W14_imag,`W2_real,`W2_imag,`W16_real,`W16_imag);
butterfly butterfly848 (clk,temp_m4_2_24_r,temp_m4_2_24_i,temp_m4_2_32_r,temp_m4_2_32_i,temp_m4_10_24_r,temp_m4_10_24_i,temp_m4_10_32_r,temp_m4_10_32_i,temp_b4_2_24_r,temp_b4_2_24_i,temp_b4_2_32_r,temp_b4_2_32_i,temp_b4_10_24_r,temp_b4_10_24_i,temp_b4_10_32_r,temp_b4_10_32_i);
MULT MULT849 (clk,temp_b3_3_17_r,temp_b3_3_17_i,temp_b3_3_25_r,temp_b3_3_25_i,temp_b3_11_17_r,temp_b3_11_17_i,temp_b3_11_25_r,temp_b3_11_25_i,temp_m4_3_17_r,temp_m4_3_17_i,temp_m4_3_25_r,temp_m4_3_25_i,temp_m4_11_17_r,temp_m4_11_17_i,temp_m4_11_25_r,temp_m4_11_25_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly849 (clk,temp_m4_3_17_r,temp_m4_3_17_i,temp_m4_3_25_r,temp_m4_3_25_i,temp_m4_11_17_r,temp_m4_11_17_i,temp_m4_11_25_r,temp_m4_11_25_i,temp_b4_3_17_r,temp_b4_3_17_i,temp_b4_3_25_r,temp_b4_3_25_i,temp_b4_11_17_r,temp_b4_11_17_i,temp_b4_11_25_r,temp_b4_11_25_i);
MULT MULT850 (clk,temp_b3_3_18_r,temp_b3_3_18_i,temp_b3_3_26_r,temp_b3_3_26_i,temp_b3_11_18_r,temp_b3_11_18_i,temp_b3_11_26_r,temp_b3_11_26_i,temp_m4_3_18_r,temp_m4_3_18_i,temp_m4_3_26_r,temp_m4_3_26_i,temp_m4_11_18_r,temp_m4_11_18_i,temp_m4_11_26_r,temp_m4_11_26_i,`W2_real,`W2_imag,`W4_real,`W4_imag,`W6_real,`W6_imag);
butterfly butterfly850 (clk,temp_m4_3_18_r,temp_m4_3_18_i,temp_m4_3_26_r,temp_m4_3_26_i,temp_m4_11_18_r,temp_m4_11_18_i,temp_m4_11_26_r,temp_m4_11_26_i,temp_b4_3_18_r,temp_b4_3_18_i,temp_b4_3_26_r,temp_b4_3_26_i,temp_b4_11_18_r,temp_b4_11_18_i,temp_b4_11_26_r,temp_b4_11_26_i);
MULT MULT851 (clk,temp_b3_3_19_r,temp_b3_3_19_i,temp_b3_3_27_r,temp_b3_3_27_i,temp_b3_11_19_r,temp_b3_11_19_i,temp_b3_11_27_r,temp_b3_11_27_i,temp_m4_3_19_r,temp_m4_3_19_i,temp_m4_3_27_r,temp_m4_3_27_i,temp_m4_11_19_r,temp_m4_11_19_i,temp_m4_11_27_r,temp_m4_11_27_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly851 (clk,temp_m4_3_19_r,temp_m4_3_19_i,temp_m4_3_27_r,temp_m4_3_27_i,temp_m4_11_19_r,temp_m4_11_19_i,temp_m4_11_27_r,temp_m4_11_27_i,temp_b4_3_19_r,temp_b4_3_19_i,temp_b4_3_27_r,temp_b4_3_27_i,temp_b4_11_19_r,temp_b4_11_19_i,temp_b4_11_27_r,temp_b4_11_27_i);
MULT MULT852 (clk,temp_b3_3_20_r,temp_b3_3_20_i,temp_b3_3_28_r,temp_b3_3_28_i,temp_b3_11_20_r,temp_b3_11_20_i,temp_b3_11_28_r,temp_b3_11_28_i,temp_m4_3_20_r,temp_m4_3_20_i,temp_m4_3_28_r,temp_m4_3_28_i,temp_m4_11_20_r,temp_m4_11_20_i,temp_m4_11_28_r,temp_m4_11_28_i,`W6_real,`W6_imag,`W4_real,`W4_imag,`W10_real,`W10_imag);
butterfly butterfly852 (clk,temp_m4_3_20_r,temp_m4_3_20_i,temp_m4_3_28_r,temp_m4_3_28_i,temp_m4_11_20_r,temp_m4_11_20_i,temp_m4_11_28_r,temp_m4_11_28_i,temp_b4_3_20_r,temp_b4_3_20_i,temp_b4_3_28_r,temp_b4_3_28_i,temp_b4_11_20_r,temp_b4_11_20_i,temp_b4_11_28_r,temp_b4_11_28_i);
MULT MULT853 (clk,temp_b3_3_21_r,temp_b3_3_21_i,temp_b3_3_29_r,temp_b3_3_29_i,temp_b3_11_21_r,temp_b3_11_21_i,temp_b3_11_29_r,temp_b3_11_29_i,temp_m4_3_21_r,temp_m4_3_21_i,temp_m4_3_29_r,temp_m4_3_29_i,temp_m4_11_21_r,temp_m4_11_21_i,temp_m4_11_29_r,temp_m4_11_29_i,`W8_real,`W8_imag,`W4_real,`W4_imag,`W12_real,`W12_imag);
butterfly butterfly853 (clk,temp_m4_3_21_r,temp_m4_3_21_i,temp_m4_3_29_r,temp_m4_3_29_i,temp_m4_11_21_r,temp_m4_11_21_i,temp_m4_11_29_r,temp_m4_11_29_i,temp_b4_3_21_r,temp_b4_3_21_i,temp_b4_3_29_r,temp_b4_3_29_i,temp_b4_11_21_r,temp_b4_11_21_i,temp_b4_11_29_r,temp_b4_11_29_i);
MULT MULT854 (clk,temp_b3_3_22_r,temp_b3_3_22_i,temp_b3_3_30_r,temp_b3_3_30_i,temp_b3_11_22_r,temp_b3_11_22_i,temp_b3_11_30_r,temp_b3_11_30_i,temp_m4_3_22_r,temp_m4_3_22_i,temp_m4_3_30_r,temp_m4_3_30_i,temp_m4_11_22_r,temp_m4_11_22_i,temp_m4_11_30_r,temp_m4_11_30_i,`W10_real,`W10_imag,`W4_real,`W4_imag,`W14_real,`W14_imag);
butterfly butterfly854 (clk,temp_m4_3_22_r,temp_m4_3_22_i,temp_m4_3_30_r,temp_m4_3_30_i,temp_m4_11_22_r,temp_m4_11_22_i,temp_m4_11_30_r,temp_m4_11_30_i,temp_b4_3_22_r,temp_b4_3_22_i,temp_b4_3_30_r,temp_b4_3_30_i,temp_b4_11_22_r,temp_b4_11_22_i,temp_b4_11_30_r,temp_b4_11_30_i);
MULT MULT855 (clk,temp_b3_3_23_r,temp_b3_3_23_i,temp_b3_3_31_r,temp_b3_3_31_i,temp_b3_11_23_r,temp_b3_11_23_i,temp_b3_11_31_r,temp_b3_11_31_i,temp_m4_3_23_r,temp_m4_3_23_i,temp_m4_3_31_r,temp_m4_3_31_i,temp_m4_11_23_r,temp_m4_11_23_i,temp_m4_11_31_r,temp_m4_11_31_i,`W12_real,`W12_imag,`W4_real,`W4_imag,`W16_real,`W16_imag);
butterfly butterfly855 (clk,temp_m4_3_23_r,temp_m4_3_23_i,temp_m4_3_31_r,temp_m4_3_31_i,temp_m4_11_23_r,temp_m4_11_23_i,temp_m4_11_31_r,temp_m4_11_31_i,temp_b4_3_23_r,temp_b4_3_23_i,temp_b4_3_31_r,temp_b4_3_31_i,temp_b4_11_23_r,temp_b4_11_23_i,temp_b4_11_31_r,temp_b4_11_31_i);
MULT MULT856 (clk,temp_b3_3_24_r,temp_b3_3_24_i,temp_b3_3_32_r,temp_b3_3_32_i,temp_b3_11_24_r,temp_b3_11_24_i,temp_b3_11_32_r,temp_b3_11_32_i,temp_m4_3_24_r,temp_m4_3_24_i,temp_m4_3_32_r,temp_m4_3_32_i,temp_m4_11_24_r,temp_m4_11_24_i,temp_m4_11_32_r,temp_m4_11_32_i,`W14_real,`W14_imag,`W4_real,`W4_imag,`W18_real,`W18_imag);
butterfly butterfly856 (clk,temp_m4_3_24_r,temp_m4_3_24_i,temp_m4_3_32_r,temp_m4_3_32_i,temp_m4_11_24_r,temp_m4_11_24_i,temp_m4_11_32_r,temp_m4_11_32_i,temp_b4_3_24_r,temp_b4_3_24_i,temp_b4_3_32_r,temp_b4_3_32_i,temp_b4_11_24_r,temp_b4_11_24_i,temp_b4_11_32_r,temp_b4_11_32_i);
MULT MULT857 (clk,temp_b3_4_17_r,temp_b3_4_17_i,temp_b3_4_25_r,temp_b3_4_25_i,temp_b3_12_17_r,temp_b3_12_17_i,temp_b3_12_25_r,temp_b3_12_25_i,temp_m4_4_17_r,temp_m4_4_17_i,temp_m4_4_25_r,temp_m4_4_25_i,temp_m4_12_17_r,temp_m4_12_17_i,temp_m4_12_25_r,temp_m4_12_25_i,`W0_real,`W0_imag,`W6_real,`W6_imag,`W6_real,`W6_imag);
butterfly butterfly857 (clk,temp_m4_4_17_r,temp_m4_4_17_i,temp_m4_4_25_r,temp_m4_4_25_i,temp_m4_12_17_r,temp_m4_12_17_i,temp_m4_12_25_r,temp_m4_12_25_i,temp_b4_4_17_r,temp_b4_4_17_i,temp_b4_4_25_r,temp_b4_4_25_i,temp_b4_12_17_r,temp_b4_12_17_i,temp_b4_12_25_r,temp_b4_12_25_i);
MULT MULT858 (clk,temp_b3_4_18_r,temp_b3_4_18_i,temp_b3_4_26_r,temp_b3_4_26_i,temp_b3_12_18_r,temp_b3_12_18_i,temp_b3_12_26_r,temp_b3_12_26_i,temp_m4_4_18_r,temp_m4_4_18_i,temp_m4_4_26_r,temp_m4_4_26_i,temp_m4_12_18_r,temp_m4_12_18_i,temp_m4_12_26_r,temp_m4_12_26_i,`W2_real,`W2_imag,`W6_real,`W6_imag,`W8_real,`W8_imag);
butterfly butterfly858 (clk,temp_m4_4_18_r,temp_m4_4_18_i,temp_m4_4_26_r,temp_m4_4_26_i,temp_m4_12_18_r,temp_m4_12_18_i,temp_m4_12_26_r,temp_m4_12_26_i,temp_b4_4_18_r,temp_b4_4_18_i,temp_b4_4_26_r,temp_b4_4_26_i,temp_b4_12_18_r,temp_b4_12_18_i,temp_b4_12_26_r,temp_b4_12_26_i);
MULT MULT859 (clk,temp_b3_4_19_r,temp_b3_4_19_i,temp_b3_4_27_r,temp_b3_4_27_i,temp_b3_12_19_r,temp_b3_12_19_i,temp_b3_12_27_r,temp_b3_12_27_i,temp_m4_4_19_r,temp_m4_4_19_i,temp_m4_4_27_r,temp_m4_4_27_i,temp_m4_12_19_r,temp_m4_12_19_i,temp_m4_12_27_r,temp_m4_12_27_i,`W4_real,`W4_imag,`W6_real,`W6_imag,`W10_real,`W10_imag);
butterfly butterfly859 (clk,temp_m4_4_19_r,temp_m4_4_19_i,temp_m4_4_27_r,temp_m4_4_27_i,temp_m4_12_19_r,temp_m4_12_19_i,temp_m4_12_27_r,temp_m4_12_27_i,temp_b4_4_19_r,temp_b4_4_19_i,temp_b4_4_27_r,temp_b4_4_27_i,temp_b4_12_19_r,temp_b4_12_19_i,temp_b4_12_27_r,temp_b4_12_27_i);
MULT MULT860 (clk,temp_b3_4_20_r,temp_b3_4_20_i,temp_b3_4_28_r,temp_b3_4_28_i,temp_b3_12_20_r,temp_b3_12_20_i,temp_b3_12_28_r,temp_b3_12_28_i,temp_m4_4_20_r,temp_m4_4_20_i,temp_m4_4_28_r,temp_m4_4_28_i,temp_m4_12_20_r,temp_m4_12_20_i,temp_m4_12_28_r,temp_m4_12_28_i,`W6_real,`W6_imag,`W6_real,`W6_imag,`W12_real,`W12_imag);
butterfly butterfly860 (clk,temp_m4_4_20_r,temp_m4_4_20_i,temp_m4_4_28_r,temp_m4_4_28_i,temp_m4_12_20_r,temp_m4_12_20_i,temp_m4_12_28_r,temp_m4_12_28_i,temp_b4_4_20_r,temp_b4_4_20_i,temp_b4_4_28_r,temp_b4_4_28_i,temp_b4_12_20_r,temp_b4_12_20_i,temp_b4_12_28_r,temp_b4_12_28_i);
MULT MULT861 (clk,temp_b3_4_21_r,temp_b3_4_21_i,temp_b3_4_29_r,temp_b3_4_29_i,temp_b3_12_21_r,temp_b3_12_21_i,temp_b3_12_29_r,temp_b3_12_29_i,temp_m4_4_21_r,temp_m4_4_21_i,temp_m4_4_29_r,temp_m4_4_29_i,temp_m4_12_21_r,temp_m4_12_21_i,temp_m4_12_29_r,temp_m4_12_29_i,`W8_real,`W8_imag,`W6_real,`W6_imag,`W14_real,`W14_imag);
butterfly butterfly861 (clk,temp_m4_4_21_r,temp_m4_4_21_i,temp_m4_4_29_r,temp_m4_4_29_i,temp_m4_12_21_r,temp_m4_12_21_i,temp_m4_12_29_r,temp_m4_12_29_i,temp_b4_4_21_r,temp_b4_4_21_i,temp_b4_4_29_r,temp_b4_4_29_i,temp_b4_12_21_r,temp_b4_12_21_i,temp_b4_12_29_r,temp_b4_12_29_i);
MULT MULT862 (clk,temp_b3_4_22_r,temp_b3_4_22_i,temp_b3_4_30_r,temp_b3_4_30_i,temp_b3_12_22_r,temp_b3_12_22_i,temp_b3_12_30_r,temp_b3_12_30_i,temp_m4_4_22_r,temp_m4_4_22_i,temp_m4_4_30_r,temp_m4_4_30_i,temp_m4_12_22_r,temp_m4_12_22_i,temp_m4_12_30_r,temp_m4_12_30_i,`W10_real,`W10_imag,`W6_real,`W6_imag,`W16_real,`W16_imag);
butterfly butterfly862 (clk,temp_m4_4_22_r,temp_m4_4_22_i,temp_m4_4_30_r,temp_m4_4_30_i,temp_m4_12_22_r,temp_m4_12_22_i,temp_m4_12_30_r,temp_m4_12_30_i,temp_b4_4_22_r,temp_b4_4_22_i,temp_b4_4_30_r,temp_b4_4_30_i,temp_b4_12_22_r,temp_b4_12_22_i,temp_b4_12_30_r,temp_b4_12_30_i);
MULT MULT863 (clk,temp_b3_4_23_r,temp_b3_4_23_i,temp_b3_4_31_r,temp_b3_4_31_i,temp_b3_12_23_r,temp_b3_12_23_i,temp_b3_12_31_r,temp_b3_12_31_i,temp_m4_4_23_r,temp_m4_4_23_i,temp_m4_4_31_r,temp_m4_4_31_i,temp_m4_12_23_r,temp_m4_12_23_i,temp_m4_12_31_r,temp_m4_12_31_i,`W12_real,`W12_imag,`W6_real,`W6_imag,`W18_real,`W18_imag);
butterfly butterfly863 (clk,temp_m4_4_23_r,temp_m4_4_23_i,temp_m4_4_31_r,temp_m4_4_31_i,temp_m4_12_23_r,temp_m4_12_23_i,temp_m4_12_31_r,temp_m4_12_31_i,temp_b4_4_23_r,temp_b4_4_23_i,temp_b4_4_31_r,temp_b4_4_31_i,temp_b4_12_23_r,temp_b4_12_23_i,temp_b4_12_31_r,temp_b4_12_31_i);
MULT MULT864 (clk,temp_b3_4_24_r,temp_b3_4_24_i,temp_b3_4_32_r,temp_b3_4_32_i,temp_b3_12_24_r,temp_b3_12_24_i,temp_b3_12_32_r,temp_b3_12_32_i,temp_m4_4_24_r,temp_m4_4_24_i,temp_m4_4_32_r,temp_m4_4_32_i,temp_m4_12_24_r,temp_m4_12_24_i,temp_m4_12_32_r,temp_m4_12_32_i,`W14_real,`W14_imag,`W6_real,`W6_imag,`W20_real,`W20_imag);
butterfly butterfly864 (clk,temp_m4_4_24_r,temp_m4_4_24_i,temp_m4_4_32_r,temp_m4_4_32_i,temp_m4_12_24_r,temp_m4_12_24_i,temp_m4_12_32_r,temp_m4_12_32_i,temp_b4_4_24_r,temp_b4_4_24_i,temp_b4_4_32_r,temp_b4_4_32_i,temp_b4_12_24_r,temp_b4_12_24_i,temp_b4_12_32_r,temp_b4_12_32_i);
MULT MULT865 (clk,temp_b3_5_17_r,temp_b3_5_17_i,temp_b3_5_25_r,temp_b3_5_25_i,temp_b3_13_17_r,temp_b3_13_17_i,temp_b3_13_25_r,temp_b3_13_25_i,temp_m4_5_17_r,temp_m4_5_17_i,temp_m4_5_25_r,temp_m4_5_25_i,temp_m4_13_17_r,temp_m4_13_17_i,temp_m4_13_25_r,temp_m4_13_25_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly865 (clk,temp_m4_5_17_r,temp_m4_5_17_i,temp_m4_5_25_r,temp_m4_5_25_i,temp_m4_13_17_r,temp_m4_13_17_i,temp_m4_13_25_r,temp_m4_13_25_i,temp_b4_5_17_r,temp_b4_5_17_i,temp_b4_5_25_r,temp_b4_5_25_i,temp_b4_13_17_r,temp_b4_13_17_i,temp_b4_13_25_r,temp_b4_13_25_i);
MULT MULT866 (clk,temp_b3_5_18_r,temp_b3_5_18_i,temp_b3_5_26_r,temp_b3_5_26_i,temp_b3_13_18_r,temp_b3_13_18_i,temp_b3_13_26_r,temp_b3_13_26_i,temp_m4_5_18_r,temp_m4_5_18_i,temp_m4_5_26_r,temp_m4_5_26_i,temp_m4_13_18_r,temp_m4_13_18_i,temp_m4_13_26_r,temp_m4_13_26_i,`W2_real,`W2_imag,`W8_real,`W8_imag,`W10_real,`W10_imag);
butterfly butterfly866 (clk,temp_m4_5_18_r,temp_m4_5_18_i,temp_m4_5_26_r,temp_m4_5_26_i,temp_m4_13_18_r,temp_m4_13_18_i,temp_m4_13_26_r,temp_m4_13_26_i,temp_b4_5_18_r,temp_b4_5_18_i,temp_b4_5_26_r,temp_b4_5_26_i,temp_b4_13_18_r,temp_b4_13_18_i,temp_b4_13_26_r,temp_b4_13_26_i);
MULT MULT867 (clk,temp_b3_5_19_r,temp_b3_5_19_i,temp_b3_5_27_r,temp_b3_5_27_i,temp_b3_13_19_r,temp_b3_13_19_i,temp_b3_13_27_r,temp_b3_13_27_i,temp_m4_5_19_r,temp_m4_5_19_i,temp_m4_5_27_r,temp_m4_5_27_i,temp_m4_13_19_r,temp_m4_13_19_i,temp_m4_13_27_r,temp_m4_13_27_i,`W4_real,`W4_imag,`W8_real,`W8_imag,`W12_real,`W12_imag);
butterfly butterfly867 (clk,temp_m4_5_19_r,temp_m4_5_19_i,temp_m4_5_27_r,temp_m4_5_27_i,temp_m4_13_19_r,temp_m4_13_19_i,temp_m4_13_27_r,temp_m4_13_27_i,temp_b4_5_19_r,temp_b4_5_19_i,temp_b4_5_27_r,temp_b4_5_27_i,temp_b4_13_19_r,temp_b4_13_19_i,temp_b4_13_27_r,temp_b4_13_27_i);
MULT MULT868 (clk,temp_b3_5_20_r,temp_b3_5_20_i,temp_b3_5_28_r,temp_b3_5_28_i,temp_b3_13_20_r,temp_b3_13_20_i,temp_b3_13_28_r,temp_b3_13_28_i,temp_m4_5_20_r,temp_m4_5_20_i,temp_m4_5_28_r,temp_m4_5_28_i,temp_m4_13_20_r,temp_m4_13_20_i,temp_m4_13_28_r,temp_m4_13_28_i,`W6_real,`W6_imag,`W8_real,`W8_imag,`W14_real,`W14_imag);
butterfly butterfly868 (clk,temp_m4_5_20_r,temp_m4_5_20_i,temp_m4_5_28_r,temp_m4_5_28_i,temp_m4_13_20_r,temp_m4_13_20_i,temp_m4_13_28_r,temp_m4_13_28_i,temp_b4_5_20_r,temp_b4_5_20_i,temp_b4_5_28_r,temp_b4_5_28_i,temp_b4_13_20_r,temp_b4_13_20_i,temp_b4_13_28_r,temp_b4_13_28_i);
MULT MULT869 (clk,temp_b3_5_21_r,temp_b3_5_21_i,temp_b3_5_29_r,temp_b3_5_29_i,temp_b3_13_21_r,temp_b3_13_21_i,temp_b3_13_29_r,temp_b3_13_29_i,temp_m4_5_21_r,temp_m4_5_21_i,temp_m4_5_29_r,temp_m4_5_29_i,temp_m4_13_21_r,temp_m4_13_21_i,temp_m4_13_29_r,temp_m4_13_29_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly869 (clk,temp_m4_5_21_r,temp_m4_5_21_i,temp_m4_5_29_r,temp_m4_5_29_i,temp_m4_13_21_r,temp_m4_13_21_i,temp_m4_13_29_r,temp_m4_13_29_i,temp_b4_5_21_r,temp_b4_5_21_i,temp_b4_5_29_r,temp_b4_5_29_i,temp_b4_13_21_r,temp_b4_13_21_i,temp_b4_13_29_r,temp_b4_13_29_i);
MULT MULT870 (clk,temp_b3_5_22_r,temp_b3_5_22_i,temp_b3_5_30_r,temp_b3_5_30_i,temp_b3_13_22_r,temp_b3_13_22_i,temp_b3_13_30_r,temp_b3_13_30_i,temp_m4_5_22_r,temp_m4_5_22_i,temp_m4_5_30_r,temp_m4_5_30_i,temp_m4_13_22_r,temp_m4_13_22_i,temp_m4_13_30_r,temp_m4_13_30_i,`W10_real,`W10_imag,`W8_real,`W8_imag,`W18_real,`W18_imag);
butterfly butterfly870 (clk,temp_m4_5_22_r,temp_m4_5_22_i,temp_m4_5_30_r,temp_m4_5_30_i,temp_m4_13_22_r,temp_m4_13_22_i,temp_m4_13_30_r,temp_m4_13_30_i,temp_b4_5_22_r,temp_b4_5_22_i,temp_b4_5_30_r,temp_b4_5_30_i,temp_b4_13_22_r,temp_b4_13_22_i,temp_b4_13_30_r,temp_b4_13_30_i);
MULT MULT871 (clk,temp_b3_5_23_r,temp_b3_5_23_i,temp_b3_5_31_r,temp_b3_5_31_i,temp_b3_13_23_r,temp_b3_13_23_i,temp_b3_13_31_r,temp_b3_13_31_i,temp_m4_5_23_r,temp_m4_5_23_i,temp_m4_5_31_r,temp_m4_5_31_i,temp_m4_13_23_r,temp_m4_13_23_i,temp_m4_13_31_r,temp_m4_13_31_i,`W12_real,`W12_imag,`W8_real,`W8_imag,`W20_real,`W20_imag);
butterfly butterfly871 (clk,temp_m4_5_23_r,temp_m4_5_23_i,temp_m4_5_31_r,temp_m4_5_31_i,temp_m4_13_23_r,temp_m4_13_23_i,temp_m4_13_31_r,temp_m4_13_31_i,temp_b4_5_23_r,temp_b4_5_23_i,temp_b4_5_31_r,temp_b4_5_31_i,temp_b4_13_23_r,temp_b4_13_23_i,temp_b4_13_31_r,temp_b4_13_31_i);
MULT MULT872 (clk,temp_b3_5_24_r,temp_b3_5_24_i,temp_b3_5_32_r,temp_b3_5_32_i,temp_b3_13_24_r,temp_b3_13_24_i,temp_b3_13_32_r,temp_b3_13_32_i,temp_m4_5_24_r,temp_m4_5_24_i,temp_m4_5_32_r,temp_m4_5_32_i,temp_m4_13_24_r,temp_m4_13_24_i,temp_m4_13_32_r,temp_m4_13_32_i,`W14_real,`W14_imag,`W8_real,`W8_imag,`W22_real,`W22_imag);
butterfly butterfly872 (clk,temp_m4_5_24_r,temp_m4_5_24_i,temp_m4_5_32_r,temp_m4_5_32_i,temp_m4_13_24_r,temp_m4_13_24_i,temp_m4_13_32_r,temp_m4_13_32_i,temp_b4_5_24_r,temp_b4_5_24_i,temp_b4_5_32_r,temp_b4_5_32_i,temp_b4_13_24_r,temp_b4_13_24_i,temp_b4_13_32_r,temp_b4_13_32_i);
MULT MULT873 (clk,temp_b3_6_17_r,temp_b3_6_17_i,temp_b3_6_25_r,temp_b3_6_25_i,temp_b3_14_17_r,temp_b3_14_17_i,temp_b3_14_25_r,temp_b3_14_25_i,temp_m4_6_17_r,temp_m4_6_17_i,temp_m4_6_25_r,temp_m4_6_25_i,temp_m4_14_17_r,temp_m4_14_17_i,temp_m4_14_25_r,temp_m4_14_25_i,`W0_real,`W0_imag,`W10_real,`W10_imag,`W10_real,`W10_imag);
butterfly butterfly873 (clk,temp_m4_6_17_r,temp_m4_6_17_i,temp_m4_6_25_r,temp_m4_6_25_i,temp_m4_14_17_r,temp_m4_14_17_i,temp_m4_14_25_r,temp_m4_14_25_i,temp_b4_6_17_r,temp_b4_6_17_i,temp_b4_6_25_r,temp_b4_6_25_i,temp_b4_14_17_r,temp_b4_14_17_i,temp_b4_14_25_r,temp_b4_14_25_i);
MULT MULT874 (clk,temp_b3_6_18_r,temp_b3_6_18_i,temp_b3_6_26_r,temp_b3_6_26_i,temp_b3_14_18_r,temp_b3_14_18_i,temp_b3_14_26_r,temp_b3_14_26_i,temp_m4_6_18_r,temp_m4_6_18_i,temp_m4_6_26_r,temp_m4_6_26_i,temp_m4_14_18_r,temp_m4_14_18_i,temp_m4_14_26_r,temp_m4_14_26_i,`W2_real,`W2_imag,`W10_real,`W10_imag,`W12_real,`W12_imag);
butterfly butterfly874 (clk,temp_m4_6_18_r,temp_m4_6_18_i,temp_m4_6_26_r,temp_m4_6_26_i,temp_m4_14_18_r,temp_m4_14_18_i,temp_m4_14_26_r,temp_m4_14_26_i,temp_b4_6_18_r,temp_b4_6_18_i,temp_b4_6_26_r,temp_b4_6_26_i,temp_b4_14_18_r,temp_b4_14_18_i,temp_b4_14_26_r,temp_b4_14_26_i);
MULT MULT875 (clk,temp_b3_6_19_r,temp_b3_6_19_i,temp_b3_6_27_r,temp_b3_6_27_i,temp_b3_14_19_r,temp_b3_14_19_i,temp_b3_14_27_r,temp_b3_14_27_i,temp_m4_6_19_r,temp_m4_6_19_i,temp_m4_6_27_r,temp_m4_6_27_i,temp_m4_14_19_r,temp_m4_14_19_i,temp_m4_14_27_r,temp_m4_14_27_i,`W4_real,`W4_imag,`W10_real,`W10_imag,`W14_real,`W14_imag);
butterfly butterfly875 (clk,temp_m4_6_19_r,temp_m4_6_19_i,temp_m4_6_27_r,temp_m4_6_27_i,temp_m4_14_19_r,temp_m4_14_19_i,temp_m4_14_27_r,temp_m4_14_27_i,temp_b4_6_19_r,temp_b4_6_19_i,temp_b4_6_27_r,temp_b4_6_27_i,temp_b4_14_19_r,temp_b4_14_19_i,temp_b4_14_27_r,temp_b4_14_27_i);
MULT MULT876 (clk,temp_b3_6_20_r,temp_b3_6_20_i,temp_b3_6_28_r,temp_b3_6_28_i,temp_b3_14_20_r,temp_b3_14_20_i,temp_b3_14_28_r,temp_b3_14_28_i,temp_m4_6_20_r,temp_m4_6_20_i,temp_m4_6_28_r,temp_m4_6_28_i,temp_m4_14_20_r,temp_m4_14_20_i,temp_m4_14_28_r,temp_m4_14_28_i,`W6_real,`W6_imag,`W10_real,`W10_imag,`W16_real,`W16_imag);
butterfly butterfly876 (clk,temp_m4_6_20_r,temp_m4_6_20_i,temp_m4_6_28_r,temp_m4_6_28_i,temp_m4_14_20_r,temp_m4_14_20_i,temp_m4_14_28_r,temp_m4_14_28_i,temp_b4_6_20_r,temp_b4_6_20_i,temp_b4_6_28_r,temp_b4_6_28_i,temp_b4_14_20_r,temp_b4_14_20_i,temp_b4_14_28_r,temp_b4_14_28_i);
MULT MULT877 (clk,temp_b3_6_21_r,temp_b3_6_21_i,temp_b3_6_29_r,temp_b3_6_29_i,temp_b3_14_21_r,temp_b3_14_21_i,temp_b3_14_29_r,temp_b3_14_29_i,temp_m4_6_21_r,temp_m4_6_21_i,temp_m4_6_29_r,temp_m4_6_29_i,temp_m4_14_21_r,temp_m4_14_21_i,temp_m4_14_29_r,temp_m4_14_29_i,`W8_real,`W8_imag,`W10_real,`W10_imag,`W18_real,`W18_imag);
butterfly butterfly877 (clk,temp_m4_6_21_r,temp_m4_6_21_i,temp_m4_6_29_r,temp_m4_6_29_i,temp_m4_14_21_r,temp_m4_14_21_i,temp_m4_14_29_r,temp_m4_14_29_i,temp_b4_6_21_r,temp_b4_6_21_i,temp_b4_6_29_r,temp_b4_6_29_i,temp_b4_14_21_r,temp_b4_14_21_i,temp_b4_14_29_r,temp_b4_14_29_i);
MULT MULT878 (clk,temp_b3_6_22_r,temp_b3_6_22_i,temp_b3_6_30_r,temp_b3_6_30_i,temp_b3_14_22_r,temp_b3_14_22_i,temp_b3_14_30_r,temp_b3_14_30_i,temp_m4_6_22_r,temp_m4_6_22_i,temp_m4_6_30_r,temp_m4_6_30_i,temp_m4_14_22_r,temp_m4_14_22_i,temp_m4_14_30_r,temp_m4_14_30_i,`W10_real,`W10_imag,`W10_real,`W10_imag,`W20_real,`W20_imag);
butterfly butterfly878 (clk,temp_m4_6_22_r,temp_m4_6_22_i,temp_m4_6_30_r,temp_m4_6_30_i,temp_m4_14_22_r,temp_m4_14_22_i,temp_m4_14_30_r,temp_m4_14_30_i,temp_b4_6_22_r,temp_b4_6_22_i,temp_b4_6_30_r,temp_b4_6_30_i,temp_b4_14_22_r,temp_b4_14_22_i,temp_b4_14_30_r,temp_b4_14_30_i);
MULT MULT879 (clk,temp_b3_6_23_r,temp_b3_6_23_i,temp_b3_6_31_r,temp_b3_6_31_i,temp_b3_14_23_r,temp_b3_14_23_i,temp_b3_14_31_r,temp_b3_14_31_i,temp_m4_6_23_r,temp_m4_6_23_i,temp_m4_6_31_r,temp_m4_6_31_i,temp_m4_14_23_r,temp_m4_14_23_i,temp_m4_14_31_r,temp_m4_14_31_i,`W12_real,`W12_imag,`W10_real,`W10_imag,`W22_real,`W22_imag);
butterfly butterfly879 (clk,temp_m4_6_23_r,temp_m4_6_23_i,temp_m4_6_31_r,temp_m4_6_31_i,temp_m4_14_23_r,temp_m4_14_23_i,temp_m4_14_31_r,temp_m4_14_31_i,temp_b4_6_23_r,temp_b4_6_23_i,temp_b4_6_31_r,temp_b4_6_31_i,temp_b4_14_23_r,temp_b4_14_23_i,temp_b4_14_31_r,temp_b4_14_31_i);
MULT MULT880 (clk,temp_b3_6_24_r,temp_b3_6_24_i,temp_b3_6_32_r,temp_b3_6_32_i,temp_b3_14_24_r,temp_b3_14_24_i,temp_b3_14_32_r,temp_b3_14_32_i,temp_m4_6_24_r,temp_m4_6_24_i,temp_m4_6_32_r,temp_m4_6_32_i,temp_m4_14_24_r,temp_m4_14_24_i,temp_m4_14_32_r,temp_m4_14_32_i,`W14_real,`W14_imag,`W10_real,`W10_imag,`W24_real,`W24_imag);
butterfly butterfly880 (clk,temp_m4_6_24_r,temp_m4_6_24_i,temp_m4_6_32_r,temp_m4_6_32_i,temp_m4_14_24_r,temp_m4_14_24_i,temp_m4_14_32_r,temp_m4_14_32_i,temp_b4_6_24_r,temp_b4_6_24_i,temp_b4_6_32_r,temp_b4_6_32_i,temp_b4_14_24_r,temp_b4_14_24_i,temp_b4_14_32_r,temp_b4_14_32_i);
MULT MULT881 (clk,temp_b3_7_17_r,temp_b3_7_17_i,temp_b3_7_25_r,temp_b3_7_25_i,temp_b3_15_17_r,temp_b3_15_17_i,temp_b3_15_25_r,temp_b3_15_25_i,temp_m4_7_17_r,temp_m4_7_17_i,temp_m4_7_25_r,temp_m4_7_25_i,temp_m4_15_17_r,temp_m4_15_17_i,temp_m4_15_25_r,temp_m4_15_25_i,`W0_real,`W0_imag,`W12_real,`W12_imag,`W12_real,`W12_imag);
butterfly butterfly881 (clk,temp_m4_7_17_r,temp_m4_7_17_i,temp_m4_7_25_r,temp_m4_7_25_i,temp_m4_15_17_r,temp_m4_15_17_i,temp_m4_15_25_r,temp_m4_15_25_i,temp_b4_7_17_r,temp_b4_7_17_i,temp_b4_7_25_r,temp_b4_7_25_i,temp_b4_15_17_r,temp_b4_15_17_i,temp_b4_15_25_r,temp_b4_15_25_i);
MULT MULT882 (clk,temp_b3_7_18_r,temp_b3_7_18_i,temp_b3_7_26_r,temp_b3_7_26_i,temp_b3_15_18_r,temp_b3_15_18_i,temp_b3_15_26_r,temp_b3_15_26_i,temp_m4_7_18_r,temp_m4_7_18_i,temp_m4_7_26_r,temp_m4_7_26_i,temp_m4_15_18_r,temp_m4_15_18_i,temp_m4_15_26_r,temp_m4_15_26_i,`W2_real,`W2_imag,`W12_real,`W12_imag,`W14_real,`W14_imag);
butterfly butterfly882 (clk,temp_m4_7_18_r,temp_m4_7_18_i,temp_m4_7_26_r,temp_m4_7_26_i,temp_m4_15_18_r,temp_m4_15_18_i,temp_m4_15_26_r,temp_m4_15_26_i,temp_b4_7_18_r,temp_b4_7_18_i,temp_b4_7_26_r,temp_b4_7_26_i,temp_b4_15_18_r,temp_b4_15_18_i,temp_b4_15_26_r,temp_b4_15_26_i);
MULT MULT883 (clk,temp_b3_7_19_r,temp_b3_7_19_i,temp_b3_7_27_r,temp_b3_7_27_i,temp_b3_15_19_r,temp_b3_15_19_i,temp_b3_15_27_r,temp_b3_15_27_i,temp_m4_7_19_r,temp_m4_7_19_i,temp_m4_7_27_r,temp_m4_7_27_i,temp_m4_15_19_r,temp_m4_15_19_i,temp_m4_15_27_r,temp_m4_15_27_i,`W4_real,`W4_imag,`W12_real,`W12_imag,`W16_real,`W16_imag);
butterfly butterfly883 (clk,temp_m4_7_19_r,temp_m4_7_19_i,temp_m4_7_27_r,temp_m4_7_27_i,temp_m4_15_19_r,temp_m4_15_19_i,temp_m4_15_27_r,temp_m4_15_27_i,temp_b4_7_19_r,temp_b4_7_19_i,temp_b4_7_27_r,temp_b4_7_27_i,temp_b4_15_19_r,temp_b4_15_19_i,temp_b4_15_27_r,temp_b4_15_27_i);
MULT MULT884 (clk,temp_b3_7_20_r,temp_b3_7_20_i,temp_b3_7_28_r,temp_b3_7_28_i,temp_b3_15_20_r,temp_b3_15_20_i,temp_b3_15_28_r,temp_b3_15_28_i,temp_m4_7_20_r,temp_m4_7_20_i,temp_m4_7_28_r,temp_m4_7_28_i,temp_m4_15_20_r,temp_m4_15_20_i,temp_m4_15_28_r,temp_m4_15_28_i,`W6_real,`W6_imag,`W12_real,`W12_imag,`W18_real,`W18_imag);
butterfly butterfly884 (clk,temp_m4_7_20_r,temp_m4_7_20_i,temp_m4_7_28_r,temp_m4_7_28_i,temp_m4_15_20_r,temp_m4_15_20_i,temp_m4_15_28_r,temp_m4_15_28_i,temp_b4_7_20_r,temp_b4_7_20_i,temp_b4_7_28_r,temp_b4_7_28_i,temp_b4_15_20_r,temp_b4_15_20_i,temp_b4_15_28_r,temp_b4_15_28_i);
MULT MULT885 (clk,temp_b3_7_21_r,temp_b3_7_21_i,temp_b3_7_29_r,temp_b3_7_29_i,temp_b3_15_21_r,temp_b3_15_21_i,temp_b3_15_29_r,temp_b3_15_29_i,temp_m4_7_21_r,temp_m4_7_21_i,temp_m4_7_29_r,temp_m4_7_29_i,temp_m4_15_21_r,temp_m4_15_21_i,temp_m4_15_29_r,temp_m4_15_29_i,`W8_real,`W8_imag,`W12_real,`W12_imag,`W20_real,`W20_imag);
butterfly butterfly885 (clk,temp_m4_7_21_r,temp_m4_7_21_i,temp_m4_7_29_r,temp_m4_7_29_i,temp_m4_15_21_r,temp_m4_15_21_i,temp_m4_15_29_r,temp_m4_15_29_i,temp_b4_7_21_r,temp_b4_7_21_i,temp_b4_7_29_r,temp_b4_7_29_i,temp_b4_15_21_r,temp_b4_15_21_i,temp_b4_15_29_r,temp_b4_15_29_i);
MULT MULT886 (clk,temp_b3_7_22_r,temp_b3_7_22_i,temp_b3_7_30_r,temp_b3_7_30_i,temp_b3_15_22_r,temp_b3_15_22_i,temp_b3_15_30_r,temp_b3_15_30_i,temp_m4_7_22_r,temp_m4_7_22_i,temp_m4_7_30_r,temp_m4_7_30_i,temp_m4_15_22_r,temp_m4_15_22_i,temp_m4_15_30_r,temp_m4_15_30_i,`W10_real,`W10_imag,`W12_real,`W12_imag,`W22_real,`W22_imag);
butterfly butterfly886 (clk,temp_m4_7_22_r,temp_m4_7_22_i,temp_m4_7_30_r,temp_m4_7_30_i,temp_m4_15_22_r,temp_m4_15_22_i,temp_m4_15_30_r,temp_m4_15_30_i,temp_b4_7_22_r,temp_b4_7_22_i,temp_b4_7_30_r,temp_b4_7_30_i,temp_b4_15_22_r,temp_b4_15_22_i,temp_b4_15_30_r,temp_b4_15_30_i);
MULT MULT887 (clk,temp_b3_7_23_r,temp_b3_7_23_i,temp_b3_7_31_r,temp_b3_7_31_i,temp_b3_15_23_r,temp_b3_15_23_i,temp_b3_15_31_r,temp_b3_15_31_i,temp_m4_7_23_r,temp_m4_7_23_i,temp_m4_7_31_r,temp_m4_7_31_i,temp_m4_15_23_r,temp_m4_15_23_i,temp_m4_15_31_r,temp_m4_15_31_i,`W12_real,`W12_imag,`W12_real,`W12_imag,`W24_real,`W24_imag);
butterfly butterfly887 (clk,temp_m4_7_23_r,temp_m4_7_23_i,temp_m4_7_31_r,temp_m4_7_31_i,temp_m4_15_23_r,temp_m4_15_23_i,temp_m4_15_31_r,temp_m4_15_31_i,temp_b4_7_23_r,temp_b4_7_23_i,temp_b4_7_31_r,temp_b4_7_31_i,temp_b4_15_23_r,temp_b4_15_23_i,temp_b4_15_31_r,temp_b4_15_31_i);
MULT MULT888 (clk,temp_b3_7_24_r,temp_b3_7_24_i,temp_b3_7_32_r,temp_b3_7_32_i,temp_b3_15_24_r,temp_b3_15_24_i,temp_b3_15_32_r,temp_b3_15_32_i,temp_m4_7_24_r,temp_m4_7_24_i,temp_m4_7_32_r,temp_m4_7_32_i,temp_m4_15_24_r,temp_m4_15_24_i,temp_m4_15_32_r,temp_m4_15_32_i,`W14_real,`W14_imag,`W12_real,`W12_imag,`W26_real,`W26_imag);
butterfly butterfly888 (clk,temp_m4_7_24_r,temp_m4_7_24_i,temp_m4_7_32_r,temp_m4_7_32_i,temp_m4_15_24_r,temp_m4_15_24_i,temp_m4_15_32_r,temp_m4_15_32_i,temp_b4_7_24_r,temp_b4_7_24_i,temp_b4_7_32_r,temp_b4_7_32_i,temp_b4_15_24_r,temp_b4_15_24_i,temp_b4_15_32_r,temp_b4_15_32_i);
MULT MULT889 (clk,temp_b3_8_17_r,temp_b3_8_17_i,temp_b3_8_25_r,temp_b3_8_25_i,temp_b3_16_17_r,temp_b3_16_17_i,temp_b3_16_25_r,temp_b3_16_25_i,temp_m4_8_17_r,temp_m4_8_17_i,temp_m4_8_25_r,temp_m4_8_25_i,temp_m4_16_17_r,temp_m4_16_17_i,temp_m4_16_25_r,temp_m4_16_25_i,`W0_real,`W0_imag,`W14_real,`W14_imag,`W14_real,`W14_imag);
butterfly butterfly889 (clk,temp_m4_8_17_r,temp_m4_8_17_i,temp_m4_8_25_r,temp_m4_8_25_i,temp_m4_16_17_r,temp_m4_16_17_i,temp_m4_16_25_r,temp_m4_16_25_i,temp_b4_8_17_r,temp_b4_8_17_i,temp_b4_8_25_r,temp_b4_8_25_i,temp_b4_16_17_r,temp_b4_16_17_i,temp_b4_16_25_r,temp_b4_16_25_i);
MULT MULT890 (clk,temp_b3_8_18_r,temp_b3_8_18_i,temp_b3_8_26_r,temp_b3_8_26_i,temp_b3_16_18_r,temp_b3_16_18_i,temp_b3_16_26_r,temp_b3_16_26_i,temp_m4_8_18_r,temp_m4_8_18_i,temp_m4_8_26_r,temp_m4_8_26_i,temp_m4_16_18_r,temp_m4_16_18_i,temp_m4_16_26_r,temp_m4_16_26_i,`W2_real,`W2_imag,`W14_real,`W14_imag,`W16_real,`W16_imag);
butterfly butterfly890 (clk,temp_m4_8_18_r,temp_m4_8_18_i,temp_m4_8_26_r,temp_m4_8_26_i,temp_m4_16_18_r,temp_m4_16_18_i,temp_m4_16_26_r,temp_m4_16_26_i,temp_b4_8_18_r,temp_b4_8_18_i,temp_b4_8_26_r,temp_b4_8_26_i,temp_b4_16_18_r,temp_b4_16_18_i,temp_b4_16_26_r,temp_b4_16_26_i);
MULT MULT891 (clk,temp_b3_8_19_r,temp_b3_8_19_i,temp_b3_8_27_r,temp_b3_8_27_i,temp_b3_16_19_r,temp_b3_16_19_i,temp_b3_16_27_r,temp_b3_16_27_i,temp_m4_8_19_r,temp_m4_8_19_i,temp_m4_8_27_r,temp_m4_8_27_i,temp_m4_16_19_r,temp_m4_16_19_i,temp_m4_16_27_r,temp_m4_16_27_i,`W4_real,`W4_imag,`W14_real,`W14_imag,`W18_real,`W18_imag);
butterfly butterfly891 (clk,temp_m4_8_19_r,temp_m4_8_19_i,temp_m4_8_27_r,temp_m4_8_27_i,temp_m4_16_19_r,temp_m4_16_19_i,temp_m4_16_27_r,temp_m4_16_27_i,temp_b4_8_19_r,temp_b4_8_19_i,temp_b4_8_27_r,temp_b4_8_27_i,temp_b4_16_19_r,temp_b4_16_19_i,temp_b4_16_27_r,temp_b4_16_27_i);
MULT MULT892 (clk,temp_b3_8_20_r,temp_b3_8_20_i,temp_b3_8_28_r,temp_b3_8_28_i,temp_b3_16_20_r,temp_b3_16_20_i,temp_b3_16_28_r,temp_b3_16_28_i,temp_m4_8_20_r,temp_m4_8_20_i,temp_m4_8_28_r,temp_m4_8_28_i,temp_m4_16_20_r,temp_m4_16_20_i,temp_m4_16_28_r,temp_m4_16_28_i,`W6_real,`W6_imag,`W14_real,`W14_imag,`W20_real,`W20_imag);
butterfly butterfly892 (clk,temp_m4_8_20_r,temp_m4_8_20_i,temp_m4_8_28_r,temp_m4_8_28_i,temp_m4_16_20_r,temp_m4_16_20_i,temp_m4_16_28_r,temp_m4_16_28_i,temp_b4_8_20_r,temp_b4_8_20_i,temp_b4_8_28_r,temp_b4_8_28_i,temp_b4_16_20_r,temp_b4_16_20_i,temp_b4_16_28_r,temp_b4_16_28_i);
MULT MULT893 (clk,temp_b3_8_21_r,temp_b3_8_21_i,temp_b3_8_29_r,temp_b3_8_29_i,temp_b3_16_21_r,temp_b3_16_21_i,temp_b3_16_29_r,temp_b3_16_29_i,temp_m4_8_21_r,temp_m4_8_21_i,temp_m4_8_29_r,temp_m4_8_29_i,temp_m4_16_21_r,temp_m4_16_21_i,temp_m4_16_29_r,temp_m4_16_29_i,`W8_real,`W8_imag,`W14_real,`W14_imag,`W22_real,`W22_imag);
butterfly butterfly893 (clk,temp_m4_8_21_r,temp_m4_8_21_i,temp_m4_8_29_r,temp_m4_8_29_i,temp_m4_16_21_r,temp_m4_16_21_i,temp_m4_16_29_r,temp_m4_16_29_i,temp_b4_8_21_r,temp_b4_8_21_i,temp_b4_8_29_r,temp_b4_8_29_i,temp_b4_16_21_r,temp_b4_16_21_i,temp_b4_16_29_r,temp_b4_16_29_i);
MULT MULT894 (clk,temp_b3_8_22_r,temp_b3_8_22_i,temp_b3_8_30_r,temp_b3_8_30_i,temp_b3_16_22_r,temp_b3_16_22_i,temp_b3_16_30_r,temp_b3_16_30_i,temp_m4_8_22_r,temp_m4_8_22_i,temp_m4_8_30_r,temp_m4_8_30_i,temp_m4_16_22_r,temp_m4_16_22_i,temp_m4_16_30_r,temp_m4_16_30_i,`W10_real,`W10_imag,`W14_real,`W14_imag,`W24_real,`W24_imag);
butterfly butterfly894 (clk,temp_m4_8_22_r,temp_m4_8_22_i,temp_m4_8_30_r,temp_m4_8_30_i,temp_m4_16_22_r,temp_m4_16_22_i,temp_m4_16_30_r,temp_m4_16_30_i,temp_b4_8_22_r,temp_b4_8_22_i,temp_b4_8_30_r,temp_b4_8_30_i,temp_b4_16_22_r,temp_b4_16_22_i,temp_b4_16_30_r,temp_b4_16_30_i);
MULT MULT895 (clk,temp_b3_8_23_r,temp_b3_8_23_i,temp_b3_8_31_r,temp_b3_8_31_i,temp_b3_16_23_r,temp_b3_16_23_i,temp_b3_16_31_r,temp_b3_16_31_i,temp_m4_8_23_r,temp_m4_8_23_i,temp_m4_8_31_r,temp_m4_8_31_i,temp_m4_16_23_r,temp_m4_16_23_i,temp_m4_16_31_r,temp_m4_16_31_i,`W12_real,`W12_imag,`W14_real,`W14_imag,`W26_real,`W26_imag);
butterfly butterfly895 (clk,temp_m4_8_23_r,temp_m4_8_23_i,temp_m4_8_31_r,temp_m4_8_31_i,temp_m4_16_23_r,temp_m4_16_23_i,temp_m4_16_31_r,temp_m4_16_31_i,temp_b4_8_23_r,temp_b4_8_23_i,temp_b4_8_31_r,temp_b4_8_31_i,temp_b4_16_23_r,temp_b4_16_23_i,temp_b4_16_31_r,temp_b4_16_31_i);
MULT MULT896 (clk,temp_b3_8_24_r,temp_b3_8_24_i,temp_b3_8_32_r,temp_b3_8_32_i,temp_b3_16_24_r,temp_b3_16_24_i,temp_b3_16_32_r,temp_b3_16_32_i,temp_m4_8_24_r,temp_m4_8_24_i,temp_m4_8_32_r,temp_m4_8_32_i,temp_m4_16_24_r,temp_m4_16_24_i,temp_m4_16_32_r,temp_m4_16_32_i,`W14_real,`W14_imag,`W14_real,`W14_imag,`W28_real,`W28_imag);
butterfly butterfly896 (clk,temp_m4_8_24_r,temp_m4_8_24_i,temp_m4_8_32_r,temp_m4_8_32_i,temp_m4_16_24_r,temp_m4_16_24_i,temp_m4_16_32_r,temp_m4_16_32_i,temp_b4_8_24_r,temp_b4_8_24_i,temp_b4_8_32_r,temp_b4_8_32_i,temp_b4_16_24_r,temp_b4_16_24_i,temp_b4_16_32_r,temp_b4_16_32_i);
MULT MULT897 (clk,temp_b3_17_1_r,temp_b3_17_1_i,temp_b3_17_9_r,temp_b3_17_9_i,temp_b3_25_1_r,temp_b3_25_1_i,temp_b3_25_9_r,temp_b3_25_9_i,temp_m4_17_1_r,temp_m4_17_1_i,temp_m4_17_9_r,temp_m4_17_9_i,temp_m4_25_1_r,temp_m4_25_1_i,temp_m4_25_9_r,temp_m4_25_9_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly897 (clk,temp_m4_17_1_r,temp_m4_17_1_i,temp_m4_17_9_r,temp_m4_17_9_i,temp_m4_25_1_r,temp_m4_25_1_i,temp_m4_25_9_r,temp_m4_25_9_i,temp_b4_17_1_r,temp_b4_17_1_i,temp_b4_17_9_r,temp_b4_17_9_i,temp_b4_25_1_r,temp_b4_25_1_i,temp_b4_25_9_r,temp_b4_25_9_i);
MULT MULT898 (clk,temp_b3_17_2_r,temp_b3_17_2_i,temp_b3_17_10_r,temp_b3_17_10_i,temp_b3_25_2_r,temp_b3_25_2_i,temp_b3_25_10_r,temp_b3_25_10_i,temp_m4_17_2_r,temp_m4_17_2_i,temp_m4_17_10_r,temp_m4_17_10_i,temp_m4_25_2_r,temp_m4_25_2_i,temp_m4_25_10_r,temp_m4_25_10_i,`W2_real,`W2_imag,`W0_real,`W0_imag,`W2_real,`W2_imag);
butterfly butterfly898 (clk,temp_m4_17_2_r,temp_m4_17_2_i,temp_m4_17_10_r,temp_m4_17_10_i,temp_m4_25_2_r,temp_m4_25_2_i,temp_m4_25_10_r,temp_m4_25_10_i,temp_b4_17_2_r,temp_b4_17_2_i,temp_b4_17_10_r,temp_b4_17_10_i,temp_b4_25_2_r,temp_b4_25_2_i,temp_b4_25_10_r,temp_b4_25_10_i);
MULT MULT899 (clk,temp_b3_17_3_r,temp_b3_17_3_i,temp_b3_17_11_r,temp_b3_17_11_i,temp_b3_25_3_r,temp_b3_25_3_i,temp_b3_25_11_r,temp_b3_25_11_i,temp_m4_17_3_r,temp_m4_17_3_i,temp_m4_17_11_r,temp_m4_17_11_i,temp_m4_25_3_r,temp_m4_25_3_i,temp_m4_25_11_r,temp_m4_25_11_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly899 (clk,temp_m4_17_3_r,temp_m4_17_3_i,temp_m4_17_11_r,temp_m4_17_11_i,temp_m4_25_3_r,temp_m4_25_3_i,temp_m4_25_11_r,temp_m4_25_11_i,temp_b4_17_3_r,temp_b4_17_3_i,temp_b4_17_11_r,temp_b4_17_11_i,temp_b4_25_3_r,temp_b4_25_3_i,temp_b4_25_11_r,temp_b4_25_11_i);
MULT MULT900 (clk,temp_b3_17_4_r,temp_b3_17_4_i,temp_b3_17_12_r,temp_b3_17_12_i,temp_b3_25_4_r,temp_b3_25_4_i,temp_b3_25_12_r,temp_b3_25_12_i,temp_m4_17_4_r,temp_m4_17_4_i,temp_m4_17_12_r,temp_m4_17_12_i,temp_m4_25_4_r,temp_m4_25_4_i,temp_m4_25_12_r,temp_m4_25_12_i,`W6_real,`W6_imag,`W0_real,`W0_imag,`W6_real,`W6_imag);
butterfly butterfly900 (clk,temp_m4_17_4_r,temp_m4_17_4_i,temp_m4_17_12_r,temp_m4_17_12_i,temp_m4_25_4_r,temp_m4_25_4_i,temp_m4_25_12_r,temp_m4_25_12_i,temp_b4_17_4_r,temp_b4_17_4_i,temp_b4_17_12_r,temp_b4_17_12_i,temp_b4_25_4_r,temp_b4_25_4_i,temp_b4_25_12_r,temp_b4_25_12_i);
MULT MULT901 (clk,temp_b3_17_5_r,temp_b3_17_5_i,temp_b3_17_13_r,temp_b3_17_13_i,temp_b3_25_5_r,temp_b3_25_5_i,temp_b3_25_13_r,temp_b3_25_13_i,temp_m4_17_5_r,temp_m4_17_5_i,temp_m4_17_13_r,temp_m4_17_13_i,temp_m4_25_5_r,temp_m4_25_5_i,temp_m4_25_13_r,temp_m4_25_13_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly901 (clk,temp_m4_17_5_r,temp_m4_17_5_i,temp_m4_17_13_r,temp_m4_17_13_i,temp_m4_25_5_r,temp_m4_25_5_i,temp_m4_25_13_r,temp_m4_25_13_i,temp_b4_17_5_r,temp_b4_17_5_i,temp_b4_17_13_r,temp_b4_17_13_i,temp_b4_25_5_r,temp_b4_25_5_i,temp_b4_25_13_r,temp_b4_25_13_i);
MULT MULT902 (clk,temp_b3_17_6_r,temp_b3_17_6_i,temp_b3_17_14_r,temp_b3_17_14_i,temp_b3_25_6_r,temp_b3_25_6_i,temp_b3_25_14_r,temp_b3_25_14_i,temp_m4_17_6_r,temp_m4_17_6_i,temp_m4_17_14_r,temp_m4_17_14_i,temp_m4_25_6_r,temp_m4_25_6_i,temp_m4_25_14_r,temp_m4_25_14_i,`W10_real,`W10_imag,`W0_real,`W0_imag,`W10_real,`W10_imag);
butterfly butterfly902 (clk,temp_m4_17_6_r,temp_m4_17_6_i,temp_m4_17_14_r,temp_m4_17_14_i,temp_m4_25_6_r,temp_m4_25_6_i,temp_m4_25_14_r,temp_m4_25_14_i,temp_b4_17_6_r,temp_b4_17_6_i,temp_b4_17_14_r,temp_b4_17_14_i,temp_b4_25_6_r,temp_b4_25_6_i,temp_b4_25_14_r,temp_b4_25_14_i);
MULT MULT903 (clk,temp_b3_17_7_r,temp_b3_17_7_i,temp_b3_17_15_r,temp_b3_17_15_i,temp_b3_25_7_r,temp_b3_25_7_i,temp_b3_25_15_r,temp_b3_25_15_i,temp_m4_17_7_r,temp_m4_17_7_i,temp_m4_17_15_r,temp_m4_17_15_i,temp_m4_25_7_r,temp_m4_25_7_i,temp_m4_25_15_r,temp_m4_25_15_i,`W12_real,`W12_imag,`W0_real,`W0_imag,`W12_real,`W12_imag);
butterfly butterfly903 (clk,temp_m4_17_7_r,temp_m4_17_7_i,temp_m4_17_15_r,temp_m4_17_15_i,temp_m4_25_7_r,temp_m4_25_7_i,temp_m4_25_15_r,temp_m4_25_15_i,temp_b4_17_7_r,temp_b4_17_7_i,temp_b4_17_15_r,temp_b4_17_15_i,temp_b4_25_7_r,temp_b4_25_7_i,temp_b4_25_15_r,temp_b4_25_15_i);
MULT MULT904 (clk,temp_b3_17_8_r,temp_b3_17_8_i,temp_b3_17_16_r,temp_b3_17_16_i,temp_b3_25_8_r,temp_b3_25_8_i,temp_b3_25_16_r,temp_b3_25_16_i,temp_m4_17_8_r,temp_m4_17_8_i,temp_m4_17_16_r,temp_m4_17_16_i,temp_m4_25_8_r,temp_m4_25_8_i,temp_m4_25_16_r,temp_m4_25_16_i,`W14_real,`W14_imag,`W0_real,`W0_imag,`W14_real,`W14_imag);
butterfly butterfly904 (clk,temp_m4_17_8_r,temp_m4_17_8_i,temp_m4_17_16_r,temp_m4_17_16_i,temp_m4_25_8_r,temp_m4_25_8_i,temp_m4_25_16_r,temp_m4_25_16_i,temp_b4_17_8_r,temp_b4_17_8_i,temp_b4_17_16_r,temp_b4_17_16_i,temp_b4_25_8_r,temp_b4_25_8_i,temp_b4_25_16_r,temp_b4_25_16_i);
MULT MULT905 (clk,temp_b3_18_1_r,temp_b3_18_1_i,temp_b3_18_9_r,temp_b3_18_9_i,temp_b3_26_1_r,temp_b3_26_1_i,temp_b3_26_9_r,temp_b3_26_9_i,temp_m4_18_1_r,temp_m4_18_1_i,temp_m4_18_9_r,temp_m4_18_9_i,temp_m4_26_1_r,temp_m4_26_1_i,temp_m4_26_9_r,temp_m4_26_9_i,`W0_real,`W0_imag,`W2_real,`W2_imag,`W2_real,`W2_imag);
butterfly butterfly905 (clk,temp_m4_18_1_r,temp_m4_18_1_i,temp_m4_18_9_r,temp_m4_18_9_i,temp_m4_26_1_r,temp_m4_26_1_i,temp_m4_26_9_r,temp_m4_26_9_i,temp_b4_18_1_r,temp_b4_18_1_i,temp_b4_18_9_r,temp_b4_18_9_i,temp_b4_26_1_r,temp_b4_26_1_i,temp_b4_26_9_r,temp_b4_26_9_i);
MULT MULT906 (clk,temp_b3_18_2_r,temp_b3_18_2_i,temp_b3_18_10_r,temp_b3_18_10_i,temp_b3_26_2_r,temp_b3_26_2_i,temp_b3_26_10_r,temp_b3_26_10_i,temp_m4_18_2_r,temp_m4_18_2_i,temp_m4_18_10_r,temp_m4_18_10_i,temp_m4_26_2_r,temp_m4_26_2_i,temp_m4_26_10_r,temp_m4_26_10_i,`W2_real,`W2_imag,`W2_real,`W2_imag,`W4_real,`W4_imag);
butterfly butterfly906 (clk,temp_m4_18_2_r,temp_m4_18_2_i,temp_m4_18_10_r,temp_m4_18_10_i,temp_m4_26_2_r,temp_m4_26_2_i,temp_m4_26_10_r,temp_m4_26_10_i,temp_b4_18_2_r,temp_b4_18_2_i,temp_b4_18_10_r,temp_b4_18_10_i,temp_b4_26_2_r,temp_b4_26_2_i,temp_b4_26_10_r,temp_b4_26_10_i);
MULT MULT907 (clk,temp_b3_18_3_r,temp_b3_18_3_i,temp_b3_18_11_r,temp_b3_18_11_i,temp_b3_26_3_r,temp_b3_26_3_i,temp_b3_26_11_r,temp_b3_26_11_i,temp_m4_18_3_r,temp_m4_18_3_i,temp_m4_18_11_r,temp_m4_18_11_i,temp_m4_26_3_r,temp_m4_26_3_i,temp_m4_26_11_r,temp_m4_26_11_i,`W4_real,`W4_imag,`W2_real,`W2_imag,`W6_real,`W6_imag);
butterfly butterfly907 (clk,temp_m4_18_3_r,temp_m4_18_3_i,temp_m4_18_11_r,temp_m4_18_11_i,temp_m4_26_3_r,temp_m4_26_3_i,temp_m4_26_11_r,temp_m4_26_11_i,temp_b4_18_3_r,temp_b4_18_3_i,temp_b4_18_11_r,temp_b4_18_11_i,temp_b4_26_3_r,temp_b4_26_3_i,temp_b4_26_11_r,temp_b4_26_11_i);
MULT MULT908 (clk,temp_b3_18_4_r,temp_b3_18_4_i,temp_b3_18_12_r,temp_b3_18_12_i,temp_b3_26_4_r,temp_b3_26_4_i,temp_b3_26_12_r,temp_b3_26_12_i,temp_m4_18_4_r,temp_m4_18_4_i,temp_m4_18_12_r,temp_m4_18_12_i,temp_m4_26_4_r,temp_m4_26_4_i,temp_m4_26_12_r,temp_m4_26_12_i,`W6_real,`W6_imag,`W2_real,`W2_imag,`W8_real,`W8_imag);
butterfly butterfly908 (clk,temp_m4_18_4_r,temp_m4_18_4_i,temp_m4_18_12_r,temp_m4_18_12_i,temp_m4_26_4_r,temp_m4_26_4_i,temp_m4_26_12_r,temp_m4_26_12_i,temp_b4_18_4_r,temp_b4_18_4_i,temp_b4_18_12_r,temp_b4_18_12_i,temp_b4_26_4_r,temp_b4_26_4_i,temp_b4_26_12_r,temp_b4_26_12_i);
MULT MULT909 (clk,temp_b3_18_5_r,temp_b3_18_5_i,temp_b3_18_13_r,temp_b3_18_13_i,temp_b3_26_5_r,temp_b3_26_5_i,temp_b3_26_13_r,temp_b3_26_13_i,temp_m4_18_5_r,temp_m4_18_5_i,temp_m4_18_13_r,temp_m4_18_13_i,temp_m4_26_5_r,temp_m4_26_5_i,temp_m4_26_13_r,temp_m4_26_13_i,`W8_real,`W8_imag,`W2_real,`W2_imag,`W10_real,`W10_imag);
butterfly butterfly909 (clk,temp_m4_18_5_r,temp_m4_18_5_i,temp_m4_18_13_r,temp_m4_18_13_i,temp_m4_26_5_r,temp_m4_26_5_i,temp_m4_26_13_r,temp_m4_26_13_i,temp_b4_18_5_r,temp_b4_18_5_i,temp_b4_18_13_r,temp_b4_18_13_i,temp_b4_26_5_r,temp_b4_26_5_i,temp_b4_26_13_r,temp_b4_26_13_i);
MULT MULT910 (clk,temp_b3_18_6_r,temp_b3_18_6_i,temp_b3_18_14_r,temp_b3_18_14_i,temp_b3_26_6_r,temp_b3_26_6_i,temp_b3_26_14_r,temp_b3_26_14_i,temp_m4_18_6_r,temp_m4_18_6_i,temp_m4_18_14_r,temp_m4_18_14_i,temp_m4_26_6_r,temp_m4_26_6_i,temp_m4_26_14_r,temp_m4_26_14_i,`W10_real,`W10_imag,`W2_real,`W2_imag,`W12_real,`W12_imag);
butterfly butterfly910 (clk,temp_m4_18_6_r,temp_m4_18_6_i,temp_m4_18_14_r,temp_m4_18_14_i,temp_m4_26_6_r,temp_m4_26_6_i,temp_m4_26_14_r,temp_m4_26_14_i,temp_b4_18_6_r,temp_b4_18_6_i,temp_b4_18_14_r,temp_b4_18_14_i,temp_b4_26_6_r,temp_b4_26_6_i,temp_b4_26_14_r,temp_b4_26_14_i);
MULT MULT911 (clk,temp_b3_18_7_r,temp_b3_18_7_i,temp_b3_18_15_r,temp_b3_18_15_i,temp_b3_26_7_r,temp_b3_26_7_i,temp_b3_26_15_r,temp_b3_26_15_i,temp_m4_18_7_r,temp_m4_18_7_i,temp_m4_18_15_r,temp_m4_18_15_i,temp_m4_26_7_r,temp_m4_26_7_i,temp_m4_26_15_r,temp_m4_26_15_i,`W12_real,`W12_imag,`W2_real,`W2_imag,`W14_real,`W14_imag);
butterfly butterfly911 (clk,temp_m4_18_7_r,temp_m4_18_7_i,temp_m4_18_15_r,temp_m4_18_15_i,temp_m4_26_7_r,temp_m4_26_7_i,temp_m4_26_15_r,temp_m4_26_15_i,temp_b4_18_7_r,temp_b4_18_7_i,temp_b4_18_15_r,temp_b4_18_15_i,temp_b4_26_7_r,temp_b4_26_7_i,temp_b4_26_15_r,temp_b4_26_15_i);
MULT MULT912 (clk,temp_b3_18_8_r,temp_b3_18_8_i,temp_b3_18_16_r,temp_b3_18_16_i,temp_b3_26_8_r,temp_b3_26_8_i,temp_b3_26_16_r,temp_b3_26_16_i,temp_m4_18_8_r,temp_m4_18_8_i,temp_m4_18_16_r,temp_m4_18_16_i,temp_m4_26_8_r,temp_m4_26_8_i,temp_m4_26_16_r,temp_m4_26_16_i,`W14_real,`W14_imag,`W2_real,`W2_imag,`W16_real,`W16_imag);
butterfly butterfly912 (clk,temp_m4_18_8_r,temp_m4_18_8_i,temp_m4_18_16_r,temp_m4_18_16_i,temp_m4_26_8_r,temp_m4_26_8_i,temp_m4_26_16_r,temp_m4_26_16_i,temp_b4_18_8_r,temp_b4_18_8_i,temp_b4_18_16_r,temp_b4_18_16_i,temp_b4_26_8_r,temp_b4_26_8_i,temp_b4_26_16_r,temp_b4_26_16_i);
MULT MULT913 (clk,temp_b3_19_1_r,temp_b3_19_1_i,temp_b3_19_9_r,temp_b3_19_9_i,temp_b3_27_1_r,temp_b3_27_1_i,temp_b3_27_9_r,temp_b3_27_9_i,temp_m4_19_1_r,temp_m4_19_1_i,temp_m4_19_9_r,temp_m4_19_9_i,temp_m4_27_1_r,temp_m4_27_1_i,temp_m4_27_9_r,temp_m4_27_9_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly913 (clk,temp_m4_19_1_r,temp_m4_19_1_i,temp_m4_19_9_r,temp_m4_19_9_i,temp_m4_27_1_r,temp_m4_27_1_i,temp_m4_27_9_r,temp_m4_27_9_i,temp_b4_19_1_r,temp_b4_19_1_i,temp_b4_19_9_r,temp_b4_19_9_i,temp_b4_27_1_r,temp_b4_27_1_i,temp_b4_27_9_r,temp_b4_27_9_i);
MULT MULT914 (clk,temp_b3_19_2_r,temp_b3_19_2_i,temp_b3_19_10_r,temp_b3_19_10_i,temp_b3_27_2_r,temp_b3_27_2_i,temp_b3_27_10_r,temp_b3_27_10_i,temp_m4_19_2_r,temp_m4_19_2_i,temp_m4_19_10_r,temp_m4_19_10_i,temp_m4_27_2_r,temp_m4_27_2_i,temp_m4_27_10_r,temp_m4_27_10_i,`W2_real,`W2_imag,`W4_real,`W4_imag,`W6_real,`W6_imag);
butterfly butterfly914 (clk,temp_m4_19_2_r,temp_m4_19_2_i,temp_m4_19_10_r,temp_m4_19_10_i,temp_m4_27_2_r,temp_m4_27_2_i,temp_m4_27_10_r,temp_m4_27_10_i,temp_b4_19_2_r,temp_b4_19_2_i,temp_b4_19_10_r,temp_b4_19_10_i,temp_b4_27_2_r,temp_b4_27_2_i,temp_b4_27_10_r,temp_b4_27_10_i);
MULT MULT915 (clk,temp_b3_19_3_r,temp_b3_19_3_i,temp_b3_19_11_r,temp_b3_19_11_i,temp_b3_27_3_r,temp_b3_27_3_i,temp_b3_27_11_r,temp_b3_27_11_i,temp_m4_19_3_r,temp_m4_19_3_i,temp_m4_19_11_r,temp_m4_19_11_i,temp_m4_27_3_r,temp_m4_27_3_i,temp_m4_27_11_r,temp_m4_27_11_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly915 (clk,temp_m4_19_3_r,temp_m4_19_3_i,temp_m4_19_11_r,temp_m4_19_11_i,temp_m4_27_3_r,temp_m4_27_3_i,temp_m4_27_11_r,temp_m4_27_11_i,temp_b4_19_3_r,temp_b4_19_3_i,temp_b4_19_11_r,temp_b4_19_11_i,temp_b4_27_3_r,temp_b4_27_3_i,temp_b4_27_11_r,temp_b4_27_11_i);
MULT MULT916 (clk,temp_b3_19_4_r,temp_b3_19_4_i,temp_b3_19_12_r,temp_b3_19_12_i,temp_b3_27_4_r,temp_b3_27_4_i,temp_b3_27_12_r,temp_b3_27_12_i,temp_m4_19_4_r,temp_m4_19_4_i,temp_m4_19_12_r,temp_m4_19_12_i,temp_m4_27_4_r,temp_m4_27_4_i,temp_m4_27_12_r,temp_m4_27_12_i,`W6_real,`W6_imag,`W4_real,`W4_imag,`W10_real,`W10_imag);
butterfly butterfly916 (clk,temp_m4_19_4_r,temp_m4_19_4_i,temp_m4_19_12_r,temp_m4_19_12_i,temp_m4_27_4_r,temp_m4_27_4_i,temp_m4_27_12_r,temp_m4_27_12_i,temp_b4_19_4_r,temp_b4_19_4_i,temp_b4_19_12_r,temp_b4_19_12_i,temp_b4_27_4_r,temp_b4_27_4_i,temp_b4_27_12_r,temp_b4_27_12_i);
MULT MULT917 (clk,temp_b3_19_5_r,temp_b3_19_5_i,temp_b3_19_13_r,temp_b3_19_13_i,temp_b3_27_5_r,temp_b3_27_5_i,temp_b3_27_13_r,temp_b3_27_13_i,temp_m4_19_5_r,temp_m4_19_5_i,temp_m4_19_13_r,temp_m4_19_13_i,temp_m4_27_5_r,temp_m4_27_5_i,temp_m4_27_13_r,temp_m4_27_13_i,`W8_real,`W8_imag,`W4_real,`W4_imag,`W12_real,`W12_imag);
butterfly butterfly917 (clk,temp_m4_19_5_r,temp_m4_19_5_i,temp_m4_19_13_r,temp_m4_19_13_i,temp_m4_27_5_r,temp_m4_27_5_i,temp_m4_27_13_r,temp_m4_27_13_i,temp_b4_19_5_r,temp_b4_19_5_i,temp_b4_19_13_r,temp_b4_19_13_i,temp_b4_27_5_r,temp_b4_27_5_i,temp_b4_27_13_r,temp_b4_27_13_i);
MULT MULT918 (clk,temp_b3_19_6_r,temp_b3_19_6_i,temp_b3_19_14_r,temp_b3_19_14_i,temp_b3_27_6_r,temp_b3_27_6_i,temp_b3_27_14_r,temp_b3_27_14_i,temp_m4_19_6_r,temp_m4_19_6_i,temp_m4_19_14_r,temp_m4_19_14_i,temp_m4_27_6_r,temp_m4_27_6_i,temp_m4_27_14_r,temp_m4_27_14_i,`W10_real,`W10_imag,`W4_real,`W4_imag,`W14_real,`W14_imag);
butterfly butterfly918 (clk,temp_m4_19_6_r,temp_m4_19_6_i,temp_m4_19_14_r,temp_m4_19_14_i,temp_m4_27_6_r,temp_m4_27_6_i,temp_m4_27_14_r,temp_m4_27_14_i,temp_b4_19_6_r,temp_b4_19_6_i,temp_b4_19_14_r,temp_b4_19_14_i,temp_b4_27_6_r,temp_b4_27_6_i,temp_b4_27_14_r,temp_b4_27_14_i);
MULT MULT919 (clk,temp_b3_19_7_r,temp_b3_19_7_i,temp_b3_19_15_r,temp_b3_19_15_i,temp_b3_27_7_r,temp_b3_27_7_i,temp_b3_27_15_r,temp_b3_27_15_i,temp_m4_19_7_r,temp_m4_19_7_i,temp_m4_19_15_r,temp_m4_19_15_i,temp_m4_27_7_r,temp_m4_27_7_i,temp_m4_27_15_r,temp_m4_27_15_i,`W12_real,`W12_imag,`W4_real,`W4_imag,`W16_real,`W16_imag);
butterfly butterfly919 (clk,temp_m4_19_7_r,temp_m4_19_7_i,temp_m4_19_15_r,temp_m4_19_15_i,temp_m4_27_7_r,temp_m4_27_7_i,temp_m4_27_15_r,temp_m4_27_15_i,temp_b4_19_7_r,temp_b4_19_7_i,temp_b4_19_15_r,temp_b4_19_15_i,temp_b4_27_7_r,temp_b4_27_7_i,temp_b4_27_15_r,temp_b4_27_15_i);
MULT MULT920 (clk,temp_b3_19_8_r,temp_b3_19_8_i,temp_b3_19_16_r,temp_b3_19_16_i,temp_b3_27_8_r,temp_b3_27_8_i,temp_b3_27_16_r,temp_b3_27_16_i,temp_m4_19_8_r,temp_m4_19_8_i,temp_m4_19_16_r,temp_m4_19_16_i,temp_m4_27_8_r,temp_m4_27_8_i,temp_m4_27_16_r,temp_m4_27_16_i,`W14_real,`W14_imag,`W4_real,`W4_imag,`W18_real,`W18_imag);
butterfly butterfly920 (clk,temp_m4_19_8_r,temp_m4_19_8_i,temp_m4_19_16_r,temp_m4_19_16_i,temp_m4_27_8_r,temp_m4_27_8_i,temp_m4_27_16_r,temp_m4_27_16_i,temp_b4_19_8_r,temp_b4_19_8_i,temp_b4_19_16_r,temp_b4_19_16_i,temp_b4_27_8_r,temp_b4_27_8_i,temp_b4_27_16_r,temp_b4_27_16_i);
MULT MULT921 (clk,temp_b3_20_1_r,temp_b3_20_1_i,temp_b3_20_9_r,temp_b3_20_9_i,temp_b3_28_1_r,temp_b3_28_1_i,temp_b3_28_9_r,temp_b3_28_9_i,temp_m4_20_1_r,temp_m4_20_1_i,temp_m4_20_9_r,temp_m4_20_9_i,temp_m4_28_1_r,temp_m4_28_1_i,temp_m4_28_9_r,temp_m4_28_9_i,`W0_real,`W0_imag,`W6_real,`W6_imag,`W6_real,`W6_imag);
butterfly butterfly921 (clk,temp_m4_20_1_r,temp_m4_20_1_i,temp_m4_20_9_r,temp_m4_20_9_i,temp_m4_28_1_r,temp_m4_28_1_i,temp_m4_28_9_r,temp_m4_28_9_i,temp_b4_20_1_r,temp_b4_20_1_i,temp_b4_20_9_r,temp_b4_20_9_i,temp_b4_28_1_r,temp_b4_28_1_i,temp_b4_28_9_r,temp_b4_28_9_i);
MULT MULT922 (clk,temp_b3_20_2_r,temp_b3_20_2_i,temp_b3_20_10_r,temp_b3_20_10_i,temp_b3_28_2_r,temp_b3_28_2_i,temp_b3_28_10_r,temp_b3_28_10_i,temp_m4_20_2_r,temp_m4_20_2_i,temp_m4_20_10_r,temp_m4_20_10_i,temp_m4_28_2_r,temp_m4_28_2_i,temp_m4_28_10_r,temp_m4_28_10_i,`W2_real,`W2_imag,`W6_real,`W6_imag,`W8_real,`W8_imag);
butterfly butterfly922 (clk,temp_m4_20_2_r,temp_m4_20_2_i,temp_m4_20_10_r,temp_m4_20_10_i,temp_m4_28_2_r,temp_m4_28_2_i,temp_m4_28_10_r,temp_m4_28_10_i,temp_b4_20_2_r,temp_b4_20_2_i,temp_b4_20_10_r,temp_b4_20_10_i,temp_b4_28_2_r,temp_b4_28_2_i,temp_b4_28_10_r,temp_b4_28_10_i);
MULT MULT923 (clk,temp_b3_20_3_r,temp_b3_20_3_i,temp_b3_20_11_r,temp_b3_20_11_i,temp_b3_28_3_r,temp_b3_28_3_i,temp_b3_28_11_r,temp_b3_28_11_i,temp_m4_20_3_r,temp_m4_20_3_i,temp_m4_20_11_r,temp_m4_20_11_i,temp_m4_28_3_r,temp_m4_28_3_i,temp_m4_28_11_r,temp_m4_28_11_i,`W4_real,`W4_imag,`W6_real,`W6_imag,`W10_real,`W10_imag);
butterfly butterfly923 (clk,temp_m4_20_3_r,temp_m4_20_3_i,temp_m4_20_11_r,temp_m4_20_11_i,temp_m4_28_3_r,temp_m4_28_3_i,temp_m4_28_11_r,temp_m4_28_11_i,temp_b4_20_3_r,temp_b4_20_3_i,temp_b4_20_11_r,temp_b4_20_11_i,temp_b4_28_3_r,temp_b4_28_3_i,temp_b4_28_11_r,temp_b4_28_11_i);
MULT MULT924 (clk,temp_b3_20_4_r,temp_b3_20_4_i,temp_b3_20_12_r,temp_b3_20_12_i,temp_b3_28_4_r,temp_b3_28_4_i,temp_b3_28_12_r,temp_b3_28_12_i,temp_m4_20_4_r,temp_m4_20_4_i,temp_m4_20_12_r,temp_m4_20_12_i,temp_m4_28_4_r,temp_m4_28_4_i,temp_m4_28_12_r,temp_m4_28_12_i,`W6_real,`W6_imag,`W6_real,`W6_imag,`W12_real,`W12_imag);
butterfly butterfly924 (clk,temp_m4_20_4_r,temp_m4_20_4_i,temp_m4_20_12_r,temp_m4_20_12_i,temp_m4_28_4_r,temp_m4_28_4_i,temp_m4_28_12_r,temp_m4_28_12_i,temp_b4_20_4_r,temp_b4_20_4_i,temp_b4_20_12_r,temp_b4_20_12_i,temp_b4_28_4_r,temp_b4_28_4_i,temp_b4_28_12_r,temp_b4_28_12_i);
MULT MULT925 (clk,temp_b3_20_5_r,temp_b3_20_5_i,temp_b3_20_13_r,temp_b3_20_13_i,temp_b3_28_5_r,temp_b3_28_5_i,temp_b3_28_13_r,temp_b3_28_13_i,temp_m4_20_5_r,temp_m4_20_5_i,temp_m4_20_13_r,temp_m4_20_13_i,temp_m4_28_5_r,temp_m4_28_5_i,temp_m4_28_13_r,temp_m4_28_13_i,`W8_real,`W8_imag,`W6_real,`W6_imag,`W14_real,`W14_imag);
butterfly butterfly925 (clk,temp_m4_20_5_r,temp_m4_20_5_i,temp_m4_20_13_r,temp_m4_20_13_i,temp_m4_28_5_r,temp_m4_28_5_i,temp_m4_28_13_r,temp_m4_28_13_i,temp_b4_20_5_r,temp_b4_20_5_i,temp_b4_20_13_r,temp_b4_20_13_i,temp_b4_28_5_r,temp_b4_28_5_i,temp_b4_28_13_r,temp_b4_28_13_i);
MULT MULT926 (clk,temp_b3_20_6_r,temp_b3_20_6_i,temp_b3_20_14_r,temp_b3_20_14_i,temp_b3_28_6_r,temp_b3_28_6_i,temp_b3_28_14_r,temp_b3_28_14_i,temp_m4_20_6_r,temp_m4_20_6_i,temp_m4_20_14_r,temp_m4_20_14_i,temp_m4_28_6_r,temp_m4_28_6_i,temp_m4_28_14_r,temp_m4_28_14_i,`W10_real,`W10_imag,`W6_real,`W6_imag,`W16_real,`W16_imag);
butterfly butterfly926 (clk,temp_m4_20_6_r,temp_m4_20_6_i,temp_m4_20_14_r,temp_m4_20_14_i,temp_m4_28_6_r,temp_m4_28_6_i,temp_m4_28_14_r,temp_m4_28_14_i,temp_b4_20_6_r,temp_b4_20_6_i,temp_b4_20_14_r,temp_b4_20_14_i,temp_b4_28_6_r,temp_b4_28_6_i,temp_b4_28_14_r,temp_b4_28_14_i);
MULT MULT927 (clk,temp_b3_20_7_r,temp_b3_20_7_i,temp_b3_20_15_r,temp_b3_20_15_i,temp_b3_28_7_r,temp_b3_28_7_i,temp_b3_28_15_r,temp_b3_28_15_i,temp_m4_20_7_r,temp_m4_20_7_i,temp_m4_20_15_r,temp_m4_20_15_i,temp_m4_28_7_r,temp_m4_28_7_i,temp_m4_28_15_r,temp_m4_28_15_i,`W12_real,`W12_imag,`W6_real,`W6_imag,`W18_real,`W18_imag);
butterfly butterfly927 (clk,temp_m4_20_7_r,temp_m4_20_7_i,temp_m4_20_15_r,temp_m4_20_15_i,temp_m4_28_7_r,temp_m4_28_7_i,temp_m4_28_15_r,temp_m4_28_15_i,temp_b4_20_7_r,temp_b4_20_7_i,temp_b4_20_15_r,temp_b4_20_15_i,temp_b4_28_7_r,temp_b4_28_7_i,temp_b4_28_15_r,temp_b4_28_15_i);
MULT MULT928 (clk,temp_b3_20_8_r,temp_b3_20_8_i,temp_b3_20_16_r,temp_b3_20_16_i,temp_b3_28_8_r,temp_b3_28_8_i,temp_b3_28_16_r,temp_b3_28_16_i,temp_m4_20_8_r,temp_m4_20_8_i,temp_m4_20_16_r,temp_m4_20_16_i,temp_m4_28_8_r,temp_m4_28_8_i,temp_m4_28_16_r,temp_m4_28_16_i,`W14_real,`W14_imag,`W6_real,`W6_imag,`W20_real,`W20_imag);
butterfly butterfly928 (clk,temp_m4_20_8_r,temp_m4_20_8_i,temp_m4_20_16_r,temp_m4_20_16_i,temp_m4_28_8_r,temp_m4_28_8_i,temp_m4_28_16_r,temp_m4_28_16_i,temp_b4_20_8_r,temp_b4_20_8_i,temp_b4_20_16_r,temp_b4_20_16_i,temp_b4_28_8_r,temp_b4_28_8_i,temp_b4_28_16_r,temp_b4_28_16_i);
MULT MULT929 (clk,temp_b3_21_1_r,temp_b3_21_1_i,temp_b3_21_9_r,temp_b3_21_9_i,temp_b3_29_1_r,temp_b3_29_1_i,temp_b3_29_9_r,temp_b3_29_9_i,temp_m4_21_1_r,temp_m4_21_1_i,temp_m4_21_9_r,temp_m4_21_9_i,temp_m4_29_1_r,temp_m4_29_1_i,temp_m4_29_9_r,temp_m4_29_9_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly929 (clk,temp_m4_21_1_r,temp_m4_21_1_i,temp_m4_21_9_r,temp_m4_21_9_i,temp_m4_29_1_r,temp_m4_29_1_i,temp_m4_29_9_r,temp_m4_29_9_i,temp_b4_21_1_r,temp_b4_21_1_i,temp_b4_21_9_r,temp_b4_21_9_i,temp_b4_29_1_r,temp_b4_29_1_i,temp_b4_29_9_r,temp_b4_29_9_i);
MULT MULT930 (clk,temp_b3_21_2_r,temp_b3_21_2_i,temp_b3_21_10_r,temp_b3_21_10_i,temp_b3_29_2_r,temp_b3_29_2_i,temp_b3_29_10_r,temp_b3_29_10_i,temp_m4_21_2_r,temp_m4_21_2_i,temp_m4_21_10_r,temp_m4_21_10_i,temp_m4_29_2_r,temp_m4_29_2_i,temp_m4_29_10_r,temp_m4_29_10_i,`W2_real,`W2_imag,`W8_real,`W8_imag,`W10_real,`W10_imag);
butterfly butterfly930 (clk,temp_m4_21_2_r,temp_m4_21_2_i,temp_m4_21_10_r,temp_m4_21_10_i,temp_m4_29_2_r,temp_m4_29_2_i,temp_m4_29_10_r,temp_m4_29_10_i,temp_b4_21_2_r,temp_b4_21_2_i,temp_b4_21_10_r,temp_b4_21_10_i,temp_b4_29_2_r,temp_b4_29_2_i,temp_b4_29_10_r,temp_b4_29_10_i);
MULT MULT931 (clk,temp_b3_21_3_r,temp_b3_21_3_i,temp_b3_21_11_r,temp_b3_21_11_i,temp_b3_29_3_r,temp_b3_29_3_i,temp_b3_29_11_r,temp_b3_29_11_i,temp_m4_21_3_r,temp_m4_21_3_i,temp_m4_21_11_r,temp_m4_21_11_i,temp_m4_29_3_r,temp_m4_29_3_i,temp_m4_29_11_r,temp_m4_29_11_i,`W4_real,`W4_imag,`W8_real,`W8_imag,`W12_real,`W12_imag);
butterfly butterfly931 (clk,temp_m4_21_3_r,temp_m4_21_3_i,temp_m4_21_11_r,temp_m4_21_11_i,temp_m4_29_3_r,temp_m4_29_3_i,temp_m4_29_11_r,temp_m4_29_11_i,temp_b4_21_3_r,temp_b4_21_3_i,temp_b4_21_11_r,temp_b4_21_11_i,temp_b4_29_3_r,temp_b4_29_3_i,temp_b4_29_11_r,temp_b4_29_11_i);
MULT MULT932 (clk,temp_b3_21_4_r,temp_b3_21_4_i,temp_b3_21_12_r,temp_b3_21_12_i,temp_b3_29_4_r,temp_b3_29_4_i,temp_b3_29_12_r,temp_b3_29_12_i,temp_m4_21_4_r,temp_m4_21_4_i,temp_m4_21_12_r,temp_m4_21_12_i,temp_m4_29_4_r,temp_m4_29_4_i,temp_m4_29_12_r,temp_m4_29_12_i,`W6_real,`W6_imag,`W8_real,`W8_imag,`W14_real,`W14_imag);
butterfly butterfly932 (clk,temp_m4_21_4_r,temp_m4_21_4_i,temp_m4_21_12_r,temp_m4_21_12_i,temp_m4_29_4_r,temp_m4_29_4_i,temp_m4_29_12_r,temp_m4_29_12_i,temp_b4_21_4_r,temp_b4_21_4_i,temp_b4_21_12_r,temp_b4_21_12_i,temp_b4_29_4_r,temp_b4_29_4_i,temp_b4_29_12_r,temp_b4_29_12_i);
MULT MULT933 (clk,temp_b3_21_5_r,temp_b3_21_5_i,temp_b3_21_13_r,temp_b3_21_13_i,temp_b3_29_5_r,temp_b3_29_5_i,temp_b3_29_13_r,temp_b3_29_13_i,temp_m4_21_5_r,temp_m4_21_5_i,temp_m4_21_13_r,temp_m4_21_13_i,temp_m4_29_5_r,temp_m4_29_5_i,temp_m4_29_13_r,temp_m4_29_13_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly933 (clk,temp_m4_21_5_r,temp_m4_21_5_i,temp_m4_21_13_r,temp_m4_21_13_i,temp_m4_29_5_r,temp_m4_29_5_i,temp_m4_29_13_r,temp_m4_29_13_i,temp_b4_21_5_r,temp_b4_21_5_i,temp_b4_21_13_r,temp_b4_21_13_i,temp_b4_29_5_r,temp_b4_29_5_i,temp_b4_29_13_r,temp_b4_29_13_i);
MULT MULT934 (clk,temp_b3_21_6_r,temp_b3_21_6_i,temp_b3_21_14_r,temp_b3_21_14_i,temp_b3_29_6_r,temp_b3_29_6_i,temp_b3_29_14_r,temp_b3_29_14_i,temp_m4_21_6_r,temp_m4_21_6_i,temp_m4_21_14_r,temp_m4_21_14_i,temp_m4_29_6_r,temp_m4_29_6_i,temp_m4_29_14_r,temp_m4_29_14_i,`W10_real,`W10_imag,`W8_real,`W8_imag,`W18_real,`W18_imag);
butterfly butterfly934 (clk,temp_m4_21_6_r,temp_m4_21_6_i,temp_m4_21_14_r,temp_m4_21_14_i,temp_m4_29_6_r,temp_m4_29_6_i,temp_m4_29_14_r,temp_m4_29_14_i,temp_b4_21_6_r,temp_b4_21_6_i,temp_b4_21_14_r,temp_b4_21_14_i,temp_b4_29_6_r,temp_b4_29_6_i,temp_b4_29_14_r,temp_b4_29_14_i);
MULT MULT935 (clk,temp_b3_21_7_r,temp_b3_21_7_i,temp_b3_21_15_r,temp_b3_21_15_i,temp_b3_29_7_r,temp_b3_29_7_i,temp_b3_29_15_r,temp_b3_29_15_i,temp_m4_21_7_r,temp_m4_21_7_i,temp_m4_21_15_r,temp_m4_21_15_i,temp_m4_29_7_r,temp_m4_29_7_i,temp_m4_29_15_r,temp_m4_29_15_i,`W12_real,`W12_imag,`W8_real,`W8_imag,`W20_real,`W20_imag);
butterfly butterfly935 (clk,temp_m4_21_7_r,temp_m4_21_7_i,temp_m4_21_15_r,temp_m4_21_15_i,temp_m4_29_7_r,temp_m4_29_7_i,temp_m4_29_15_r,temp_m4_29_15_i,temp_b4_21_7_r,temp_b4_21_7_i,temp_b4_21_15_r,temp_b4_21_15_i,temp_b4_29_7_r,temp_b4_29_7_i,temp_b4_29_15_r,temp_b4_29_15_i);
MULT MULT936 (clk,temp_b3_21_8_r,temp_b3_21_8_i,temp_b3_21_16_r,temp_b3_21_16_i,temp_b3_29_8_r,temp_b3_29_8_i,temp_b3_29_16_r,temp_b3_29_16_i,temp_m4_21_8_r,temp_m4_21_8_i,temp_m4_21_16_r,temp_m4_21_16_i,temp_m4_29_8_r,temp_m4_29_8_i,temp_m4_29_16_r,temp_m4_29_16_i,`W14_real,`W14_imag,`W8_real,`W8_imag,`W22_real,`W22_imag);
butterfly butterfly936 (clk,temp_m4_21_8_r,temp_m4_21_8_i,temp_m4_21_16_r,temp_m4_21_16_i,temp_m4_29_8_r,temp_m4_29_8_i,temp_m4_29_16_r,temp_m4_29_16_i,temp_b4_21_8_r,temp_b4_21_8_i,temp_b4_21_16_r,temp_b4_21_16_i,temp_b4_29_8_r,temp_b4_29_8_i,temp_b4_29_16_r,temp_b4_29_16_i);
MULT MULT937 (clk,temp_b3_22_1_r,temp_b3_22_1_i,temp_b3_22_9_r,temp_b3_22_9_i,temp_b3_30_1_r,temp_b3_30_1_i,temp_b3_30_9_r,temp_b3_30_9_i,temp_m4_22_1_r,temp_m4_22_1_i,temp_m4_22_9_r,temp_m4_22_9_i,temp_m4_30_1_r,temp_m4_30_1_i,temp_m4_30_9_r,temp_m4_30_9_i,`W0_real,`W0_imag,`W10_real,`W10_imag,`W10_real,`W10_imag);
butterfly butterfly937 (clk,temp_m4_22_1_r,temp_m4_22_1_i,temp_m4_22_9_r,temp_m4_22_9_i,temp_m4_30_1_r,temp_m4_30_1_i,temp_m4_30_9_r,temp_m4_30_9_i,temp_b4_22_1_r,temp_b4_22_1_i,temp_b4_22_9_r,temp_b4_22_9_i,temp_b4_30_1_r,temp_b4_30_1_i,temp_b4_30_9_r,temp_b4_30_9_i);
MULT MULT938 (clk,temp_b3_22_2_r,temp_b3_22_2_i,temp_b3_22_10_r,temp_b3_22_10_i,temp_b3_30_2_r,temp_b3_30_2_i,temp_b3_30_10_r,temp_b3_30_10_i,temp_m4_22_2_r,temp_m4_22_2_i,temp_m4_22_10_r,temp_m4_22_10_i,temp_m4_30_2_r,temp_m4_30_2_i,temp_m4_30_10_r,temp_m4_30_10_i,`W2_real,`W2_imag,`W10_real,`W10_imag,`W12_real,`W12_imag);
butterfly butterfly938 (clk,temp_m4_22_2_r,temp_m4_22_2_i,temp_m4_22_10_r,temp_m4_22_10_i,temp_m4_30_2_r,temp_m4_30_2_i,temp_m4_30_10_r,temp_m4_30_10_i,temp_b4_22_2_r,temp_b4_22_2_i,temp_b4_22_10_r,temp_b4_22_10_i,temp_b4_30_2_r,temp_b4_30_2_i,temp_b4_30_10_r,temp_b4_30_10_i);
MULT MULT939 (clk,temp_b3_22_3_r,temp_b3_22_3_i,temp_b3_22_11_r,temp_b3_22_11_i,temp_b3_30_3_r,temp_b3_30_3_i,temp_b3_30_11_r,temp_b3_30_11_i,temp_m4_22_3_r,temp_m4_22_3_i,temp_m4_22_11_r,temp_m4_22_11_i,temp_m4_30_3_r,temp_m4_30_3_i,temp_m4_30_11_r,temp_m4_30_11_i,`W4_real,`W4_imag,`W10_real,`W10_imag,`W14_real,`W14_imag);
butterfly butterfly939 (clk,temp_m4_22_3_r,temp_m4_22_3_i,temp_m4_22_11_r,temp_m4_22_11_i,temp_m4_30_3_r,temp_m4_30_3_i,temp_m4_30_11_r,temp_m4_30_11_i,temp_b4_22_3_r,temp_b4_22_3_i,temp_b4_22_11_r,temp_b4_22_11_i,temp_b4_30_3_r,temp_b4_30_3_i,temp_b4_30_11_r,temp_b4_30_11_i);
MULT MULT940 (clk,temp_b3_22_4_r,temp_b3_22_4_i,temp_b3_22_12_r,temp_b3_22_12_i,temp_b3_30_4_r,temp_b3_30_4_i,temp_b3_30_12_r,temp_b3_30_12_i,temp_m4_22_4_r,temp_m4_22_4_i,temp_m4_22_12_r,temp_m4_22_12_i,temp_m4_30_4_r,temp_m4_30_4_i,temp_m4_30_12_r,temp_m4_30_12_i,`W6_real,`W6_imag,`W10_real,`W10_imag,`W16_real,`W16_imag);
butterfly butterfly940 (clk,temp_m4_22_4_r,temp_m4_22_4_i,temp_m4_22_12_r,temp_m4_22_12_i,temp_m4_30_4_r,temp_m4_30_4_i,temp_m4_30_12_r,temp_m4_30_12_i,temp_b4_22_4_r,temp_b4_22_4_i,temp_b4_22_12_r,temp_b4_22_12_i,temp_b4_30_4_r,temp_b4_30_4_i,temp_b4_30_12_r,temp_b4_30_12_i);
MULT MULT941 (clk,temp_b3_22_5_r,temp_b3_22_5_i,temp_b3_22_13_r,temp_b3_22_13_i,temp_b3_30_5_r,temp_b3_30_5_i,temp_b3_30_13_r,temp_b3_30_13_i,temp_m4_22_5_r,temp_m4_22_5_i,temp_m4_22_13_r,temp_m4_22_13_i,temp_m4_30_5_r,temp_m4_30_5_i,temp_m4_30_13_r,temp_m4_30_13_i,`W8_real,`W8_imag,`W10_real,`W10_imag,`W18_real,`W18_imag);
butterfly butterfly941 (clk,temp_m4_22_5_r,temp_m4_22_5_i,temp_m4_22_13_r,temp_m4_22_13_i,temp_m4_30_5_r,temp_m4_30_5_i,temp_m4_30_13_r,temp_m4_30_13_i,temp_b4_22_5_r,temp_b4_22_5_i,temp_b4_22_13_r,temp_b4_22_13_i,temp_b4_30_5_r,temp_b4_30_5_i,temp_b4_30_13_r,temp_b4_30_13_i);
MULT MULT942 (clk,temp_b3_22_6_r,temp_b3_22_6_i,temp_b3_22_14_r,temp_b3_22_14_i,temp_b3_30_6_r,temp_b3_30_6_i,temp_b3_30_14_r,temp_b3_30_14_i,temp_m4_22_6_r,temp_m4_22_6_i,temp_m4_22_14_r,temp_m4_22_14_i,temp_m4_30_6_r,temp_m4_30_6_i,temp_m4_30_14_r,temp_m4_30_14_i,`W10_real,`W10_imag,`W10_real,`W10_imag,`W20_real,`W20_imag);
butterfly butterfly942 (clk,temp_m4_22_6_r,temp_m4_22_6_i,temp_m4_22_14_r,temp_m4_22_14_i,temp_m4_30_6_r,temp_m4_30_6_i,temp_m4_30_14_r,temp_m4_30_14_i,temp_b4_22_6_r,temp_b4_22_6_i,temp_b4_22_14_r,temp_b4_22_14_i,temp_b4_30_6_r,temp_b4_30_6_i,temp_b4_30_14_r,temp_b4_30_14_i);
MULT MULT943 (clk,temp_b3_22_7_r,temp_b3_22_7_i,temp_b3_22_15_r,temp_b3_22_15_i,temp_b3_30_7_r,temp_b3_30_7_i,temp_b3_30_15_r,temp_b3_30_15_i,temp_m4_22_7_r,temp_m4_22_7_i,temp_m4_22_15_r,temp_m4_22_15_i,temp_m4_30_7_r,temp_m4_30_7_i,temp_m4_30_15_r,temp_m4_30_15_i,`W12_real,`W12_imag,`W10_real,`W10_imag,`W22_real,`W22_imag);
butterfly butterfly943 (clk,temp_m4_22_7_r,temp_m4_22_7_i,temp_m4_22_15_r,temp_m4_22_15_i,temp_m4_30_7_r,temp_m4_30_7_i,temp_m4_30_15_r,temp_m4_30_15_i,temp_b4_22_7_r,temp_b4_22_7_i,temp_b4_22_15_r,temp_b4_22_15_i,temp_b4_30_7_r,temp_b4_30_7_i,temp_b4_30_15_r,temp_b4_30_15_i);
MULT MULT944 (clk,temp_b3_22_8_r,temp_b3_22_8_i,temp_b3_22_16_r,temp_b3_22_16_i,temp_b3_30_8_r,temp_b3_30_8_i,temp_b3_30_16_r,temp_b3_30_16_i,temp_m4_22_8_r,temp_m4_22_8_i,temp_m4_22_16_r,temp_m4_22_16_i,temp_m4_30_8_r,temp_m4_30_8_i,temp_m4_30_16_r,temp_m4_30_16_i,`W14_real,`W14_imag,`W10_real,`W10_imag,`W24_real,`W24_imag);
butterfly butterfly944 (clk,temp_m4_22_8_r,temp_m4_22_8_i,temp_m4_22_16_r,temp_m4_22_16_i,temp_m4_30_8_r,temp_m4_30_8_i,temp_m4_30_16_r,temp_m4_30_16_i,temp_b4_22_8_r,temp_b4_22_8_i,temp_b4_22_16_r,temp_b4_22_16_i,temp_b4_30_8_r,temp_b4_30_8_i,temp_b4_30_16_r,temp_b4_30_16_i);
MULT MULT945 (clk,temp_b3_23_1_r,temp_b3_23_1_i,temp_b3_23_9_r,temp_b3_23_9_i,temp_b3_31_1_r,temp_b3_31_1_i,temp_b3_31_9_r,temp_b3_31_9_i,temp_m4_23_1_r,temp_m4_23_1_i,temp_m4_23_9_r,temp_m4_23_9_i,temp_m4_31_1_r,temp_m4_31_1_i,temp_m4_31_9_r,temp_m4_31_9_i,`W0_real,`W0_imag,`W12_real,`W12_imag,`W12_real,`W12_imag);
butterfly butterfly945 (clk,temp_m4_23_1_r,temp_m4_23_1_i,temp_m4_23_9_r,temp_m4_23_9_i,temp_m4_31_1_r,temp_m4_31_1_i,temp_m4_31_9_r,temp_m4_31_9_i,temp_b4_23_1_r,temp_b4_23_1_i,temp_b4_23_9_r,temp_b4_23_9_i,temp_b4_31_1_r,temp_b4_31_1_i,temp_b4_31_9_r,temp_b4_31_9_i);
MULT MULT946 (clk,temp_b3_23_2_r,temp_b3_23_2_i,temp_b3_23_10_r,temp_b3_23_10_i,temp_b3_31_2_r,temp_b3_31_2_i,temp_b3_31_10_r,temp_b3_31_10_i,temp_m4_23_2_r,temp_m4_23_2_i,temp_m4_23_10_r,temp_m4_23_10_i,temp_m4_31_2_r,temp_m4_31_2_i,temp_m4_31_10_r,temp_m4_31_10_i,`W2_real,`W2_imag,`W12_real,`W12_imag,`W14_real,`W14_imag);
butterfly butterfly946 (clk,temp_m4_23_2_r,temp_m4_23_2_i,temp_m4_23_10_r,temp_m4_23_10_i,temp_m4_31_2_r,temp_m4_31_2_i,temp_m4_31_10_r,temp_m4_31_10_i,temp_b4_23_2_r,temp_b4_23_2_i,temp_b4_23_10_r,temp_b4_23_10_i,temp_b4_31_2_r,temp_b4_31_2_i,temp_b4_31_10_r,temp_b4_31_10_i);
MULT MULT947 (clk,temp_b3_23_3_r,temp_b3_23_3_i,temp_b3_23_11_r,temp_b3_23_11_i,temp_b3_31_3_r,temp_b3_31_3_i,temp_b3_31_11_r,temp_b3_31_11_i,temp_m4_23_3_r,temp_m4_23_3_i,temp_m4_23_11_r,temp_m4_23_11_i,temp_m4_31_3_r,temp_m4_31_3_i,temp_m4_31_11_r,temp_m4_31_11_i,`W4_real,`W4_imag,`W12_real,`W12_imag,`W16_real,`W16_imag);
butterfly butterfly947 (clk,temp_m4_23_3_r,temp_m4_23_3_i,temp_m4_23_11_r,temp_m4_23_11_i,temp_m4_31_3_r,temp_m4_31_3_i,temp_m4_31_11_r,temp_m4_31_11_i,temp_b4_23_3_r,temp_b4_23_3_i,temp_b4_23_11_r,temp_b4_23_11_i,temp_b4_31_3_r,temp_b4_31_3_i,temp_b4_31_11_r,temp_b4_31_11_i);
MULT MULT948 (clk,temp_b3_23_4_r,temp_b3_23_4_i,temp_b3_23_12_r,temp_b3_23_12_i,temp_b3_31_4_r,temp_b3_31_4_i,temp_b3_31_12_r,temp_b3_31_12_i,temp_m4_23_4_r,temp_m4_23_4_i,temp_m4_23_12_r,temp_m4_23_12_i,temp_m4_31_4_r,temp_m4_31_4_i,temp_m4_31_12_r,temp_m4_31_12_i,`W6_real,`W6_imag,`W12_real,`W12_imag,`W18_real,`W18_imag);
butterfly butterfly948 (clk,temp_m4_23_4_r,temp_m4_23_4_i,temp_m4_23_12_r,temp_m4_23_12_i,temp_m4_31_4_r,temp_m4_31_4_i,temp_m4_31_12_r,temp_m4_31_12_i,temp_b4_23_4_r,temp_b4_23_4_i,temp_b4_23_12_r,temp_b4_23_12_i,temp_b4_31_4_r,temp_b4_31_4_i,temp_b4_31_12_r,temp_b4_31_12_i);
MULT MULT949 (clk,temp_b3_23_5_r,temp_b3_23_5_i,temp_b3_23_13_r,temp_b3_23_13_i,temp_b3_31_5_r,temp_b3_31_5_i,temp_b3_31_13_r,temp_b3_31_13_i,temp_m4_23_5_r,temp_m4_23_5_i,temp_m4_23_13_r,temp_m4_23_13_i,temp_m4_31_5_r,temp_m4_31_5_i,temp_m4_31_13_r,temp_m4_31_13_i,`W8_real,`W8_imag,`W12_real,`W12_imag,`W20_real,`W20_imag);
butterfly butterfly949 (clk,temp_m4_23_5_r,temp_m4_23_5_i,temp_m4_23_13_r,temp_m4_23_13_i,temp_m4_31_5_r,temp_m4_31_5_i,temp_m4_31_13_r,temp_m4_31_13_i,temp_b4_23_5_r,temp_b4_23_5_i,temp_b4_23_13_r,temp_b4_23_13_i,temp_b4_31_5_r,temp_b4_31_5_i,temp_b4_31_13_r,temp_b4_31_13_i);
MULT MULT950 (clk,temp_b3_23_6_r,temp_b3_23_6_i,temp_b3_23_14_r,temp_b3_23_14_i,temp_b3_31_6_r,temp_b3_31_6_i,temp_b3_31_14_r,temp_b3_31_14_i,temp_m4_23_6_r,temp_m4_23_6_i,temp_m4_23_14_r,temp_m4_23_14_i,temp_m4_31_6_r,temp_m4_31_6_i,temp_m4_31_14_r,temp_m4_31_14_i,`W10_real,`W10_imag,`W12_real,`W12_imag,`W22_real,`W22_imag);
butterfly butterfly950 (clk,temp_m4_23_6_r,temp_m4_23_6_i,temp_m4_23_14_r,temp_m4_23_14_i,temp_m4_31_6_r,temp_m4_31_6_i,temp_m4_31_14_r,temp_m4_31_14_i,temp_b4_23_6_r,temp_b4_23_6_i,temp_b4_23_14_r,temp_b4_23_14_i,temp_b4_31_6_r,temp_b4_31_6_i,temp_b4_31_14_r,temp_b4_31_14_i);
MULT MULT951 (clk,temp_b3_23_7_r,temp_b3_23_7_i,temp_b3_23_15_r,temp_b3_23_15_i,temp_b3_31_7_r,temp_b3_31_7_i,temp_b3_31_15_r,temp_b3_31_15_i,temp_m4_23_7_r,temp_m4_23_7_i,temp_m4_23_15_r,temp_m4_23_15_i,temp_m4_31_7_r,temp_m4_31_7_i,temp_m4_31_15_r,temp_m4_31_15_i,`W12_real,`W12_imag,`W12_real,`W12_imag,`W24_real,`W24_imag);
butterfly butterfly951 (clk,temp_m4_23_7_r,temp_m4_23_7_i,temp_m4_23_15_r,temp_m4_23_15_i,temp_m4_31_7_r,temp_m4_31_7_i,temp_m4_31_15_r,temp_m4_31_15_i,temp_b4_23_7_r,temp_b4_23_7_i,temp_b4_23_15_r,temp_b4_23_15_i,temp_b4_31_7_r,temp_b4_31_7_i,temp_b4_31_15_r,temp_b4_31_15_i);
MULT MULT952 (clk,temp_b3_23_8_r,temp_b3_23_8_i,temp_b3_23_16_r,temp_b3_23_16_i,temp_b3_31_8_r,temp_b3_31_8_i,temp_b3_31_16_r,temp_b3_31_16_i,temp_m4_23_8_r,temp_m4_23_8_i,temp_m4_23_16_r,temp_m4_23_16_i,temp_m4_31_8_r,temp_m4_31_8_i,temp_m4_31_16_r,temp_m4_31_16_i,`W14_real,`W14_imag,`W12_real,`W12_imag,`W26_real,`W26_imag);
butterfly butterfly952 (clk,temp_m4_23_8_r,temp_m4_23_8_i,temp_m4_23_16_r,temp_m4_23_16_i,temp_m4_31_8_r,temp_m4_31_8_i,temp_m4_31_16_r,temp_m4_31_16_i,temp_b4_23_8_r,temp_b4_23_8_i,temp_b4_23_16_r,temp_b4_23_16_i,temp_b4_31_8_r,temp_b4_31_8_i,temp_b4_31_16_r,temp_b4_31_16_i);
MULT MULT953 (clk,temp_b3_24_1_r,temp_b3_24_1_i,temp_b3_24_9_r,temp_b3_24_9_i,temp_b3_32_1_r,temp_b3_32_1_i,temp_b3_32_9_r,temp_b3_32_9_i,temp_m4_24_1_r,temp_m4_24_1_i,temp_m4_24_9_r,temp_m4_24_9_i,temp_m4_32_1_r,temp_m4_32_1_i,temp_m4_32_9_r,temp_m4_32_9_i,`W0_real,`W0_imag,`W14_real,`W14_imag,`W14_real,`W14_imag);
butterfly butterfly953 (clk,temp_m4_24_1_r,temp_m4_24_1_i,temp_m4_24_9_r,temp_m4_24_9_i,temp_m4_32_1_r,temp_m4_32_1_i,temp_m4_32_9_r,temp_m4_32_9_i,temp_b4_24_1_r,temp_b4_24_1_i,temp_b4_24_9_r,temp_b4_24_9_i,temp_b4_32_1_r,temp_b4_32_1_i,temp_b4_32_9_r,temp_b4_32_9_i);
MULT MULT954 (clk,temp_b3_24_2_r,temp_b3_24_2_i,temp_b3_24_10_r,temp_b3_24_10_i,temp_b3_32_2_r,temp_b3_32_2_i,temp_b3_32_10_r,temp_b3_32_10_i,temp_m4_24_2_r,temp_m4_24_2_i,temp_m4_24_10_r,temp_m4_24_10_i,temp_m4_32_2_r,temp_m4_32_2_i,temp_m4_32_10_r,temp_m4_32_10_i,`W2_real,`W2_imag,`W14_real,`W14_imag,`W16_real,`W16_imag);
butterfly butterfly954 (clk,temp_m4_24_2_r,temp_m4_24_2_i,temp_m4_24_10_r,temp_m4_24_10_i,temp_m4_32_2_r,temp_m4_32_2_i,temp_m4_32_10_r,temp_m4_32_10_i,temp_b4_24_2_r,temp_b4_24_2_i,temp_b4_24_10_r,temp_b4_24_10_i,temp_b4_32_2_r,temp_b4_32_2_i,temp_b4_32_10_r,temp_b4_32_10_i);
MULT MULT955 (clk,temp_b3_24_3_r,temp_b3_24_3_i,temp_b3_24_11_r,temp_b3_24_11_i,temp_b3_32_3_r,temp_b3_32_3_i,temp_b3_32_11_r,temp_b3_32_11_i,temp_m4_24_3_r,temp_m4_24_3_i,temp_m4_24_11_r,temp_m4_24_11_i,temp_m4_32_3_r,temp_m4_32_3_i,temp_m4_32_11_r,temp_m4_32_11_i,`W4_real,`W4_imag,`W14_real,`W14_imag,`W18_real,`W18_imag);
butterfly butterfly955 (clk,temp_m4_24_3_r,temp_m4_24_3_i,temp_m4_24_11_r,temp_m4_24_11_i,temp_m4_32_3_r,temp_m4_32_3_i,temp_m4_32_11_r,temp_m4_32_11_i,temp_b4_24_3_r,temp_b4_24_3_i,temp_b4_24_11_r,temp_b4_24_11_i,temp_b4_32_3_r,temp_b4_32_3_i,temp_b4_32_11_r,temp_b4_32_11_i);
MULT MULT956 (clk,temp_b3_24_4_r,temp_b3_24_4_i,temp_b3_24_12_r,temp_b3_24_12_i,temp_b3_32_4_r,temp_b3_32_4_i,temp_b3_32_12_r,temp_b3_32_12_i,temp_m4_24_4_r,temp_m4_24_4_i,temp_m4_24_12_r,temp_m4_24_12_i,temp_m4_32_4_r,temp_m4_32_4_i,temp_m4_32_12_r,temp_m4_32_12_i,`W6_real,`W6_imag,`W14_real,`W14_imag,`W20_real,`W20_imag);
butterfly butterfly956 (clk,temp_m4_24_4_r,temp_m4_24_4_i,temp_m4_24_12_r,temp_m4_24_12_i,temp_m4_32_4_r,temp_m4_32_4_i,temp_m4_32_12_r,temp_m4_32_12_i,temp_b4_24_4_r,temp_b4_24_4_i,temp_b4_24_12_r,temp_b4_24_12_i,temp_b4_32_4_r,temp_b4_32_4_i,temp_b4_32_12_r,temp_b4_32_12_i);
MULT MULT957 (clk,temp_b3_24_5_r,temp_b3_24_5_i,temp_b3_24_13_r,temp_b3_24_13_i,temp_b3_32_5_r,temp_b3_32_5_i,temp_b3_32_13_r,temp_b3_32_13_i,temp_m4_24_5_r,temp_m4_24_5_i,temp_m4_24_13_r,temp_m4_24_13_i,temp_m4_32_5_r,temp_m4_32_5_i,temp_m4_32_13_r,temp_m4_32_13_i,`W8_real,`W8_imag,`W14_real,`W14_imag,`W22_real,`W22_imag);
butterfly butterfly957 (clk,temp_m4_24_5_r,temp_m4_24_5_i,temp_m4_24_13_r,temp_m4_24_13_i,temp_m4_32_5_r,temp_m4_32_5_i,temp_m4_32_13_r,temp_m4_32_13_i,temp_b4_24_5_r,temp_b4_24_5_i,temp_b4_24_13_r,temp_b4_24_13_i,temp_b4_32_5_r,temp_b4_32_5_i,temp_b4_32_13_r,temp_b4_32_13_i);
MULT MULT958 (clk,temp_b3_24_6_r,temp_b3_24_6_i,temp_b3_24_14_r,temp_b3_24_14_i,temp_b3_32_6_r,temp_b3_32_6_i,temp_b3_32_14_r,temp_b3_32_14_i,temp_m4_24_6_r,temp_m4_24_6_i,temp_m4_24_14_r,temp_m4_24_14_i,temp_m4_32_6_r,temp_m4_32_6_i,temp_m4_32_14_r,temp_m4_32_14_i,`W10_real,`W10_imag,`W14_real,`W14_imag,`W24_real,`W24_imag);
butterfly butterfly958 (clk,temp_m4_24_6_r,temp_m4_24_6_i,temp_m4_24_14_r,temp_m4_24_14_i,temp_m4_32_6_r,temp_m4_32_6_i,temp_m4_32_14_r,temp_m4_32_14_i,temp_b4_24_6_r,temp_b4_24_6_i,temp_b4_24_14_r,temp_b4_24_14_i,temp_b4_32_6_r,temp_b4_32_6_i,temp_b4_32_14_r,temp_b4_32_14_i);
MULT MULT959 (clk,temp_b3_24_7_r,temp_b3_24_7_i,temp_b3_24_15_r,temp_b3_24_15_i,temp_b3_32_7_r,temp_b3_32_7_i,temp_b3_32_15_r,temp_b3_32_15_i,temp_m4_24_7_r,temp_m4_24_7_i,temp_m4_24_15_r,temp_m4_24_15_i,temp_m4_32_7_r,temp_m4_32_7_i,temp_m4_32_15_r,temp_m4_32_15_i,`W12_real,`W12_imag,`W14_real,`W14_imag,`W26_real,`W26_imag);
butterfly butterfly959 (clk,temp_m4_24_7_r,temp_m4_24_7_i,temp_m4_24_15_r,temp_m4_24_15_i,temp_m4_32_7_r,temp_m4_32_7_i,temp_m4_32_15_r,temp_m4_32_15_i,temp_b4_24_7_r,temp_b4_24_7_i,temp_b4_24_15_r,temp_b4_24_15_i,temp_b4_32_7_r,temp_b4_32_7_i,temp_b4_32_15_r,temp_b4_32_15_i);
MULT MULT960 (clk,temp_b3_24_8_r,temp_b3_24_8_i,temp_b3_24_16_r,temp_b3_24_16_i,temp_b3_32_8_r,temp_b3_32_8_i,temp_b3_32_16_r,temp_b3_32_16_i,temp_m4_24_8_r,temp_m4_24_8_i,temp_m4_24_16_r,temp_m4_24_16_i,temp_m4_32_8_r,temp_m4_32_8_i,temp_m4_32_16_r,temp_m4_32_16_i,`W14_real,`W14_imag,`W14_real,`W14_imag,`W28_real,`W28_imag);
butterfly butterfly960 (clk,temp_m4_24_8_r,temp_m4_24_8_i,temp_m4_24_16_r,temp_m4_24_16_i,temp_m4_32_8_r,temp_m4_32_8_i,temp_m4_32_16_r,temp_m4_32_16_i,temp_b4_24_8_r,temp_b4_24_8_i,temp_b4_24_16_r,temp_b4_24_16_i,temp_b4_32_8_r,temp_b4_32_8_i,temp_b4_32_16_r,temp_b4_32_16_i);
MULT MULT961 (clk,temp_b3_17_17_r,temp_b3_17_17_i,temp_b3_17_25_r,temp_b3_17_25_i,temp_b3_25_17_r,temp_b3_25_17_i,temp_b3_25_25_r,temp_b3_25_25_i,temp_m4_17_17_r,temp_m4_17_17_i,temp_m4_17_25_r,temp_m4_17_25_i,temp_m4_25_17_r,temp_m4_25_17_i,temp_m4_25_25_r,temp_m4_25_25_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly961 (clk,temp_m4_17_17_r,temp_m4_17_17_i,temp_m4_17_25_r,temp_m4_17_25_i,temp_m4_25_17_r,temp_m4_25_17_i,temp_m4_25_25_r,temp_m4_25_25_i,temp_b4_17_17_r,temp_b4_17_17_i,temp_b4_17_25_r,temp_b4_17_25_i,temp_b4_25_17_r,temp_b4_25_17_i,temp_b4_25_25_r,temp_b4_25_25_i);
MULT MULT962 (clk,temp_b3_17_18_r,temp_b3_17_18_i,temp_b3_17_26_r,temp_b3_17_26_i,temp_b3_25_18_r,temp_b3_25_18_i,temp_b3_25_26_r,temp_b3_25_26_i,temp_m4_17_18_r,temp_m4_17_18_i,temp_m4_17_26_r,temp_m4_17_26_i,temp_m4_25_18_r,temp_m4_25_18_i,temp_m4_25_26_r,temp_m4_25_26_i,`W2_real,`W2_imag,`W0_real,`W0_imag,`W2_real,`W2_imag);
butterfly butterfly962 (clk,temp_m4_17_18_r,temp_m4_17_18_i,temp_m4_17_26_r,temp_m4_17_26_i,temp_m4_25_18_r,temp_m4_25_18_i,temp_m4_25_26_r,temp_m4_25_26_i,temp_b4_17_18_r,temp_b4_17_18_i,temp_b4_17_26_r,temp_b4_17_26_i,temp_b4_25_18_r,temp_b4_25_18_i,temp_b4_25_26_r,temp_b4_25_26_i);
MULT MULT963 (clk,temp_b3_17_19_r,temp_b3_17_19_i,temp_b3_17_27_r,temp_b3_17_27_i,temp_b3_25_19_r,temp_b3_25_19_i,temp_b3_25_27_r,temp_b3_25_27_i,temp_m4_17_19_r,temp_m4_17_19_i,temp_m4_17_27_r,temp_m4_17_27_i,temp_m4_25_19_r,temp_m4_25_19_i,temp_m4_25_27_r,temp_m4_25_27_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly963 (clk,temp_m4_17_19_r,temp_m4_17_19_i,temp_m4_17_27_r,temp_m4_17_27_i,temp_m4_25_19_r,temp_m4_25_19_i,temp_m4_25_27_r,temp_m4_25_27_i,temp_b4_17_19_r,temp_b4_17_19_i,temp_b4_17_27_r,temp_b4_17_27_i,temp_b4_25_19_r,temp_b4_25_19_i,temp_b4_25_27_r,temp_b4_25_27_i);
MULT MULT964 (clk,temp_b3_17_20_r,temp_b3_17_20_i,temp_b3_17_28_r,temp_b3_17_28_i,temp_b3_25_20_r,temp_b3_25_20_i,temp_b3_25_28_r,temp_b3_25_28_i,temp_m4_17_20_r,temp_m4_17_20_i,temp_m4_17_28_r,temp_m4_17_28_i,temp_m4_25_20_r,temp_m4_25_20_i,temp_m4_25_28_r,temp_m4_25_28_i,`W6_real,`W6_imag,`W0_real,`W0_imag,`W6_real,`W6_imag);
butterfly butterfly964 (clk,temp_m4_17_20_r,temp_m4_17_20_i,temp_m4_17_28_r,temp_m4_17_28_i,temp_m4_25_20_r,temp_m4_25_20_i,temp_m4_25_28_r,temp_m4_25_28_i,temp_b4_17_20_r,temp_b4_17_20_i,temp_b4_17_28_r,temp_b4_17_28_i,temp_b4_25_20_r,temp_b4_25_20_i,temp_b4_25_28_r,temp_b4_25_28_i);
MULT MULT965 (clk,temp_b3_17_21_r,temp_b3_17_21_i,temp_b3_17_29_r,temp_b3_17_29_i,temp_b3_25_21_r,temp_b3_25_21_i,temp_b3_25_29_r,temp_b3_25_29_i,temp_m4_17_21_r,temp_m4_17_21_i,temp_m4_17_29_r,temp_m4_17_29_i,temp_m4_25_21_r,temp_m4_25_21_i,temp_m4_25_29_r,temp_m4_25_29_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly965 (clk,temp_m4_17_21_r,temp_m4_17_21_i,temp_m4_17_29_r,temp_m4_17_29_i,temp_m4_25_21_r,temp_m4_25_21_i,temp_m4_25_29_r,temp_m4_25_29_i,temp_b4_17_21_r,temp_b4_17_21_i,temp_b4_17_29_r,temp_b4_17_29_i,temp_b4_25_21_r,temp_b4_25_21_i,temp_b4_25_29_r,temp_b4_25_29_i);
MULT MULT966 (clk,temp_b3_17_22_r,temp_b3_17_22_i,temp_b3_17_30_r,temp_b3_17_30_i,temp_b3_25_22_r,temp_b3_25_22_i,temp_b3_25_30_r,temp_b3_25_30_i,temp_m4_17_22_r,temp_m4_17_22_i,temp_m4_17_30_r,temp_m4_17_30_i,temp_m4_25_22_r,temp_m4_25_22_i,temp_m4_25_30_r,temp_m4_25_30_i,`W10_real,`W10_imag,`W0_real,`W0_imag,`W10_real,`W10_imag);
butterfly butterfly966 (clk,temp_m4_17_22_r,temp_m4_17_22_i,temp_m4_17_30_r,temp_m4_17_30_i,temp_m4_25_22_r,temp_m4_25_22_i,temp_m4_25_30_r,temp_m4_25_30_i,temp_b4_17_22_r,temp_b4_17_22_i,temp_b4_17_30_r,temp_b4_17_30_i,temp_b4_25_22_r,temp_b4_25_22_i,temp_b4_25_30_r,temp_b4_25_30_i);
MULT MULT967 (clk,temp_b3_17_23_r,temp_b3_17_23_i,temp_b3_17_31_r,temp_b3_17_31_i,temp_b3_25_23_r,temp_b3_25_23_i,temp_b3_25_31_r,temp_b3_25_31_i,temp_m4_17_23_r,temp_m4_17_23_i,temp_m4_17_31_r,temp_m4_17_31_i,temp_m4_25_23_r,temp_m4_25_23_i,temp_m4_25_31_r,temp_m4_25_31_i,`W12_real,`W12_imag,`W0_real,`W0_imag,`W12_real,`W12_imag);
butterfly butterfly967 (clk,temp_m4_17_23_r,temp_m4_17_23_i,temp_m4_17_31_r,temp_m4_17_31_i,temp_m4_25_23_r,temp_m4_25_23_i,temp_m4_25_31_r,temp_m4_25_31_i,temp_b4_17_23_r,temp_b4_17_23_i,temp_b4_17_31_r,temp_b4_17_31_i,temp_b4_25_23_r,temp_b4_25_23_i,temp_b4_25_31_r,temp_b4_25_31_i);
MULT MULT968 (clk,temp_b3_17_24_r,temp_b3_17_24_i,temp_b3_17_32_r,temp_b3_17_32_i,temp_b3_25_24_r,temp_b3_25_24_i,temp_b3_25_32_r,temp_b3_25_32_i,temp_m4_17_24_r,temp_m4_17_24_i,temp_m4_17_32_r,temp_m4_17_32_i,temp_m4_25_24_r,temp_m4_25_24_i,temp_m4_25_32_r,temp_m4_25_32_i,`W14_real,`W14_imag,`W0_real,`W0_imag,`W14_real,`W14_imag);
butterfly butterfly968 (clk,temp_m4_17_24_r,temp_m4_17_24_i,temp_m4_17_32_r,temp_m4_17_32_i,temp_m4_25_24_r,temp_m4_25_24_i,temp_m4_25_32_r,temp_m4_25_32_i,temp_b4_17_24_r,temp_b4_17_24_i,temp_b4_17_32_r,temp_b4_17_32_i,temp_b4_25_24_r,temp_b4_25_24_i,temp_b4_25_32_r,temp_b4_25_32_i);
MULT MULT969 (clk,temp_b3_18_17_r,temp_b3_18_17_i,temp_b3_18_25_r,temp_b3_18_25_i,temp_b3_26_17_r,temp_b3_26_17_i,temp_b3_26_25_r,temp_b3_26_25_i,temp_m4_18_17_r,temp_m4_18_17_i,temp_m4_18_25_r,temp_m4_18_25_i,temp_m4_26_17_r,temp_m4_26_17_i,temp_m4_26_25_r,temp_m4_26_25_i,`W0_real,`W0_imag,`W2_real,`W2_imag,`W2_real,`W2_imag);
butterfly butterfly969 (clk,temp_m4_18_17_r,temp_m4_18_17_i,temp_m4_18_25_r,temp_m4_18_25_i,temp_m4_26_17_r,temp_m4_26_17_i,temp_m4_26_25_r,temp_m4_26_25_i,temp_b4_18_17_r,temp_b4_18_17_i,temp_b4_18_25_r,temp_b4_18_25_i,temp_b4_26_17_r,temp_b4_26_17_i,temp_b4_26_25_r,temp_b4_26_25_i);
MULT MULT970 (clk,temp_b3_18_18_r,temp_b3_18_18_i,temp_b3_18_26_r,temp_b3_18_26_i,temp_b3_26_18_r,temp_b3_26_18_i,temp_b3_26_26_r,temp_b3_26_26_i,temp_m4_18_18_r,temp_m4_18_18_i,temp_m4_18_26_r,temp_m4_18_26_i,temp_m4_26_18_r,temp_m4_26_18_i,temp_m4_26_26_r,temp_m4_26_26_i,`W2_real,`W2_imag,`W2_real,`W2_imag,`W4_real,`W4_imag);
butterfly butterfly970 (clk,temp_m4_18_18_r,temp_m4_18_18_i,temp_m4_18_26_r,temp_m4_18_26_i,temp_m4_26_18_r,temp_m4_26_18_i,temp_m4_26_26_r,temp_m4_26_26_i,temp_b4_18_18_r,temp_b4_18_18_i,temp_b4_18_26_r,temp_b4_18_26_i,temp_b4_26_18_r,temp_b4_26_18_i,temp_b4_26_26_r,temp_b4_26_26_i);
MULT MULT971 (clk,temp_b3_18_19_r,temp_b3_18_19_i,temp_b3_18_27_r,temp_b3_18_27_i,temp_b3_26_19_r,temp_b3_26_19_i,temp_b3_26_27_r,temp_b3_26_27_i,temp_m4_18_19_r,temp_m4_18_19_i,temp_m4_18_27_r,temp_m4_18_27_i,temp_m4_26_19_r,temp_m4_26_19_i,temp_m4_26_27_r,temp_m4_26_27_i,`W4_real,`W4_imag,`W2_real,`W2_imag,`W6_real,`W6_imag);
butterfly butterfly971 (clk,temp_m4_18_19_r,temp_m4_18_19_i,temp_m4_18_27_r,temp_m4_18_27_i,temp_m4_26_19_r,temp_m4_26_19_i,temp_m4_26_27_r,temp_m4_26_27_i,temp_b4_18_19_r,temp_b4_18_19_i,temp_b4_18_27_r,temp_b4_18_27_i,temp_b4_26_19_r,temp_b4_26_19_i,temp_b4_26_27_r,temp_b4_26_27_i);
MULT MULT972 (clk,temp_b3_18_20_r,temp_b3_18_20_i,temp_b3_18_28_r,temp_b3_18_28_i,temp_b3_26_20_r,temp_b3_26_20_i,temp_b3_26_28_r,temp_b3_26_28_i,temp_m4_18_20_r,temp_m4_18_20_i,temp_m4_18_28_r,temp_m4_18_28_i,temp_m4_26_20_r,temp_m4_26_20_i,temp_m4_26_28_r,temp_m4_26_28_i,`W6_real,`W6_imag,`W2_real,`W2_imag,`W8_real,`W8_imag);
butterfly butterfly972 (clk,temp_m4_18_20_r,temp_m4_18_20_i,temp_m4_18_28_r,temp_m4_18_28_i,temp_m4_26_20_r,temp_m4_26_20_i,temp_m4_26_28_r,temp_m4_26_28_i,temp_b4_18_20_r,temp_b4_18_20_i,temp_b4_18_28_r,temp_b4_18_28_i,temp_b4_26_20_r,temp_b4_26_20_i,temp_b4_26_28_r,temp_b4_26_28_i);
MULT MULT973 (clk,temp_b3_18_21_r,temp_b3_18_21_i,temp_b3_18_29_r,temp_b3_18_29_i,temp_b3_26_21_r,temp_b3_26_21_i,temp_b3_26_29_r,temp_b3_26_29_i,temp_m4_18_21_r,temp_m4_18_21_i,temp_m4_18_29_r,temp_m4_18_29_i,temp_m4_26_21_r,temp_m4_26_21_i,temp_m4_26_29_r,temp_m4_26_29_i,`W8_real,`W8_imag,`W2_real,`W2_imag,`W10_real,`W10_imag);
butterfly butterfly973 (clk,temp_m4_18_21_r,temp_m4_18_21_i,temp_m4_18_29_r,temp_m4_18_29_i,temp_m4_26_21_r,temp_m4_26_21_i,temp_m4_26_29_r,temp_m4_26_29_i,temp_b4_18_21_r,temp_b4_18_21_i,temp_b4_18_29_r,temp_b4_18_29_i,temp_b4_26_21_r,temp_b4_26_21_i,temp_b4_26_29_r,temp_b4_26_29_i);
MULT MULT974 (clk,temp_b3_18_22_r,temp_b3_18_22_i,temp_b3_18_30_r,temp_b3_18_30_i,temp_b3_26_22_r,temp_b3_26_22_i,temp_b3_26_30_r,temp_b3_26_30_i,temp_m4_18_22_r,temp_m4_18_22_i,temp_m4_18_30_r,temp_m4_18_30_i,temp_m4_26_22_r,temp_m4_26_22_i,temp_m4_26_30_r,temp_m4_26_30_i,`W10_real,`W10_imag,`W2_real,`W2_imag,`W12_real,`W12_imag);
butterfly butterfly974 (clk,temp_m4_18_22_r,temp_m4_18_22_i,temp_m4_18_30_r,temp_m4_18_30_i,temp_m4_26_22_r,temp_m4_26_22_i,temp_m4_26_30_r,temp_m4_26_30_i,temp_b4_18_22_r,temp_b4_18_22_i,temp_b4_18_30_r,temp_b4_18_30_i,temp_b4_26_22_r,temp_b4_26_22_i,temp_b4_26_30_r,temp_b4_26_30_i);
MULT MULT975 (clk,temp_b3_18_23_r,temp_b3_18_23_i,temp_b3_18_31_r,temp_b3_18_31_i,temp_b3_26_23_r,temp_b3_26_23_i,temp_b3_26_31_r,temp_b3_26_31_i,temp_m4_18_23_r,temp_m4_18_23_i,temp_m4_18_31_r,temp_m4_18_31_i,temp_m4_26_23_r,temp_m4_26_23_i,temp_m4_26_31_r,temp_m4_26_31_i,`W12_real,`W12_imag,`W2_real,`W2_imag,`W14_real,`W14_imag);
butterfly butterfly975 (clk,temp_m4_18_23_r,temp_m4_18_23_i,temp_m4_18_31_r,temp_m4_18_31_i,temp_m4_26_23_r,temp_m4_26_23_i,temp_m4_26_31_r,temp_m4_26_31_i,temp_b4_18_23_r,temp_b4_18_23_i,temp_b4_18_31_r,temp_b4_18_31_i,temp_b4_26_23_r,temp_b4_26_23_i,temp_b4_26_31_r,temp_b4_26_31_i);
MULT MULT976 (clk,temp_b3_18_24_r,temp_b3_18_24_i,temp_b3_18_32_r,temp_b3_18_32_i,temp_b3_26_24_r,temp_b3_26_24_i,temp_b3_26_32_r,temp_b3_26_32_i,temp_m4_18_24_r,temp_m4_18_24_i,temp_m4_18_32_r,temp_m4_18_32_i,temp_m4_26_24_r,temp_m4_26_24_i,temp_m4_26_32_r,temp_m4_26_32_i,`W14_real,`W14_imag,`W2_real,`W2_imag,`W16_real,`W16_imag);
butterfly butterfly976 (clk,temp_m4_18_24_r,temp_m4_18_24_i,temp_m4_18_32_r,temp_m4_18_32_i,temp_m4_26_24_r,temp_m4_26_24_i,temp_m4_26_32_r,temp_m4_26_32_i,temp_b4_18_24_r,temp_b4_18_24_i,temp_b4_18_32_r,temp_b4_18_32_i,temp_b4_26_24_r,temp_b4_26_24_i,temp_b4_26_32_r,temp_b4_26_32_i);
MULT MULT977 (clk,temp_b3_19_17_r,temp_b3_19_17_i,temp_b3_19_25_r,temp_b3_19_25_i,temp_b3_27_17_r,temp_b3_27_17_i,temp_b3_27_25_r,temp_b3_27_25_i,temp_m4_19_17_r,temp_m4_19_17_i,temp_m4_19_25_r,temp_m4_19_25_i,temp_m4_27_17_r,temp_m4_27_17_i,temp_m4_27_25_r,temp_m4_27_25_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly977 (clk,temp_m4_19_17_r,temp_m4_19_17_i,temp_m4_19_25_r,temp_m4_19_25_i,temp_m4_27_17_r,temp_m4_27_17_i,temp_m4_27_25_r,temp_m4_27_25_i,temp_b4_19_17_r,temp_b4_19_17_i,temp_b4_19_25_r,temp_b4_19_25_i,temp_b4_27_17_r,temp_b4_27_17_i,temp_b4_27_25_r,temp_b4_27_25_i);
MULT MULT978 (clk,temp_b3_19_18_r,temp_b3_19_18_i,temp_b3_19_26_r,temp_b3_19_26_i,temp_b3_27_18_r,temp_b3_27_18_i,temp_b3_27_26_r,temp_b3_27_26_i,temp_m4_19_18_r,temp_m4_19_18_i,temp_m4_19_26_r,temp_m4_19_26_i,temp_m4_27_18_r,temp_m4_27_18_i,temp_m4_27_26_r,temp_m4_27_26_i,`W2_real,`W2_imag,`W4_real,`W4_imag,`W6_real,`W6_imag);
butterfly butterfly978 (clk,temp_m4_19_18_r,temp_m4_19_18_i,temp_m4_19_26_r,temp_m4_19_26_i,temp_m4_27_18_r,temp_m4_27_18_i,temp_m4_27_26_r,temp_m4_27_26_i,temp_b4_19_18_r,temp_b4_19_18_i,temp_b4_19_26_r,temp_b4_19_26_i,temp_b4_27_18_r,temp_b4_27_18_i,temp_b4_27_26_r,temp_b4_27_26_i);
MULT MULT979 (clk,temp_b3_19_19_r,temp_b3_19_19_i,temp_b3_19_27_r,temp_b3_19_27_i,temp_b3_27_19_r,temp_b3_27_19_i,temp_b3_27_27_r,temp_b3_27_27_i,temp_m4_19_19_r,temp_m4_19_19_i,temp_m4_19_27_r,temp_m4_19_27_i,temp_m4_27_19_r,temp_m4_27_19_i,temp_m4_27_27_r,temp_m4_27_27_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly979 (clk,temp_m4_19_19_r,temp_m4_19_19_i,temp_m4_19_27_r,temp_m4_19_27_i,temp_m4_27_19_r,temp_m4_27_19_i,temp_m4_27_27_r,temp_m4_27_27_i,temp_b4_19_19_r,temp_b4_19_19_i,temp_b4_19_27_r,temp_b4_19_27_i,temp_b4_27_19_r,temp_b4_27_19_i,temp_b4_27_27_r,temp_b4_27_27_i);
MULT MULT980 (clk,temp_b3_19_20_r,temp_b3_19_20_i,temp_b3_19_28_r,temp_b3_19_28_i,temp_b3_27_20_r,temp_b3_27_20_i,temp_b3_27_28_r,temp_b3_27_28_i,temp_m4_19_20_r,temp_m4_19_20_i,temp_m4_19_28_r,temp_m4_19_28_i,temp_m4_27_20_r,temp_m4_27_20_i,temp_m4_27_28_r,temp_m4_27_28_i,`W6_real,`W6_imag,`W4_real,`W4_imag,`W10_real,`W10_imag);
butterfly butterfly980 (clk,temp_m4_19_20_r,temp_m4_19_20_i,temp_m4_19_28_r,temp_m4_19_28_i,temp_m4_27_20_r,temp_m4_27_20_i,temp_m4_27_28_r,temp_m4_27_28_i,temp_b4_19_20_r,temp_b4_19_20_i,temp_b4_19_28_r,temp_b4_19_28_i,temp_b4_27_20_r,temp_b4_27_20_i,temp_b4_27_28_r,temp_b4_27_28_i);
MULT MULT981 (clk,temp_b3_19_21_r,temp_b3_19_21_i,temp_b3_19_29_r,temp_b3_19_29_i,temp_b3_27_21_r,temp_b3_27_21_i,temp_b3_27_29_r,temp_b3_27_29_i,temp_m4_19_21_r,temp_m4_19_21_i,temp_m4_19_29_r,temp_m4_19_29_i,temp_m4_27_21_r,temp_m4_27_21_i,temp_m4_27_29_r,temp_m4_27_29_i,`W8_real,`W8_imag,`W4_real,`W4_imag,`W12_real,`W12_imag);
butterfly butterfly981 (clk,temp_m4_19_21_r,temp_m4_19_21_i,temp_m4_19_29_r,temp_m4_19_29_i,temp_m4_27_21_r,temp_m4_27_21_i,temp_m4_27_29_r,temp_m4_27_29_i,temp_b4_19_21_r,temp_b4_19_21_i,temp_b4_19_29_r,temp_b4_19_29_i,temp_b4_27_21_r,temp_b4_27_21_i,temp_b4_27_29_r,temp_b4_27_29_i);
MULT MULT982 (clk,temp_b3_19_22_r,temp_b3_19_22_i,temp_b3_19_30_r,temp_b3_19_30_i,temp_b3_27_22_r,temp_b3_27_22_i,temp_b3_27_30_r,temp_b3_27_30_i,temp_m4_19_22_r,temp_m4_19_22_i,temp_m4_19_30_r,temp_m4_19_30_i,temp_m4_27_22_r,temp_m4_27_22_i,temp_m4_27_30_r,temp_m4_27_30_i,`W10_real,`W10_imag,`W4_real,`W4_imag,`W14_real,`W14_imag);
butterfly butterfly982 (clk,temp_m4_19_22_r,temp_m4_19_22_i,temp_m4_19_30_r,temp_m4_19_30_i,temp_m4_27_22_r,temp_m4_27_22_i,temp_m4_27_30_r,temp_m4_27_30_i,temp_b4_19_22_r,temp_b4_19_22_i,temp_b4_19_30_r,temp_b4_19_30_i,temp_b4_27_22_r,temp_b4_27_22_i,temp_b4_27_30_r,temp_b4_27_30_i);
MULT MULT983 (clk,temp_b3_19_23_r,temp_b3_19_23_i,temp_b3_19_31_r,temp_b3_19_31_i,temp_b3_27_23_r,temp_b3_27_23_i,temp_b3_27_31_r,temp_b3_27_31_i,temp_m4_19_23_r,temp_m4_19_23_i,temp_m4_19_31_r,temp_m4_19_31_i,temp_m4_27_23_r,temp_m4_27_23_i,temp_m4_27_31_r,temp_m4_27_31_i,`W12_real,`W12_imag,`W4_real,`W4_imag,`W16_real,`W16_imag);
butterfly butterfly983 (clk,temp_m4_19_23_r,temp_m4_19_23_i,temp_m4_19_31_r,temp_m4_19_31_i,temp_m4_27_23_r,temp_m4_27_23_i,temp_m4_27_31_r,temp_m4_27_31_i,temp_b4_19_23_r,temp_b4_19_23_i,temp_b4_19_31_r,temp_b4_19_31_i,temp_b4_27_23_r,temp_b4_27_23_i,temp_b4_27_31_r,temp_b4_27_31_i);
MULT MULT984 (clk,temp_b3_19_24_r,temp_b3_19_24_i,temp_b3_19_32_r,temp_b3_19_32_i,temp_b3_27_24_r,temp_b3_27_24_i,temp_b3_27_32_r,temp_b3_27_32_i,temp_m4_19_24_r,temp_m4_19_24_i,temp_m4_19_32_r,temp_m4_19_32_i,temp_m4_27_24_r,temp_m4_27_24_i,temp_m4_27_32_r,temp_m4_27_32_i,`W14_real,`W14_imag,`W4_real,`W4_imag,`W18_real,`W18_imag);
butterfly butterfly984 (clk,temp_m4_19_24_r,temp_m4_19_24_i,temp_m4_19_32_r,temp_m4_19_32_i,temp_m4_27_24_r,temp_m4_27_24_i,temp_m4_27_32_r,temp_m4_27_32_i,temp_b4_19_24_r,temp_b4_19_24_i,temp_b4_19_32_r,temp_b4_19_32_i,temp_b4_27_24_r,temp_b4_27_24_i,temp_b4_27_32_r,temp_b4_27_32_i);
MULT MULT985 (clk,temp_b3_20_17_r,temp_b3_20_17_i,temp_b3_20_25_r,temp_b3_20_25_i,temp_b3_28_17_r,temp_b3_28_17_i,temp_b3_28_25_r,temp_b3_28_25_i,temp_m4_20_17_r,temp_m4_20_17_i,temp_m4_20_25_r,temp_m4_20_25_i,temp_m4_28_17_r,temp_m4_28_17_i,temp_m4_28_25_r,temp_m4_28_25_i,`W0_real,`W0_imag,`W6_real,`W6_imag,`W6_real,`W6_imag);
butterfly butterfly985 (clk,temp_m4_20_17_r,temp_m4_20_17_i,temp_m4_20_25_r,temp_m4_20_25_i,temp_m4_28_17_r,temp_m4_28_17_i,temp_m4_28_25_r,temp_m4_28_25_i,temp_b4_20_17_r,temp_b4_20_17_i,temp_b4_20_25_r,temp_b4_20_25_i,temp_b4_28_17_r,temp_b4_28_17_i,temp_b4_28_25_r,temp_b4_28_25_i);
MULT MULT986 (clk,temp_b3_20_18_r,temp_b3_20_18_i,temp_b3_20_26_r,temp_b3_20_26_i,temp_b3_28_18_r,temp_b3_28_18_i,temp_b3_28_26_r,temp_b3_28_26_i,temp_m4_20_18_r,temp_m4_20_18_i,temp_m4_20_26_r,temp_m4_20_26_i,temp_m4_28_18_r,temp_m4_28_18_i,temp_m4_28_26_r,temp_m4_28_26_i,`W2_real,`W2_imag,`W6_real,`W6_imag,`W8_real,`W8_imag);
butterfly butterfly986 (clk,temp_m4_20_18_r,temp_m4_20_18_i,temp_m4_20_26_r,temp_m4_20_26_i,temp_m4_28_18_r,temp_m4_28_18_i,temp_m4_28_26_r,temp_m4_28_26_i,temp_b4_20_18_r,temp_b4_20_18_i,temp_b4_20_26_r,temp_b4_20_26_i,temp_b4_28_18_r,temp_b4_28_18_i,temp_b4_28_26_r,temp_b4_28_26_i);
MULT MULT987 (clk,temp_b3_20_19_r,temp_b3_20_19_i,temp_b3_20_27_r,temp_b3_20_27_i,temp_b3_28_19_r,temp_b3_28_19_i,temp_b3_28_27_r,temp_b3_28_27_i,temp_m4_20_19_r,temp_m4_20_19_i,temp_m4_20_27_r,temp_m4_20_27_i,temp_m4_28_19_r,temp_m4_28_19_i,temp_m4_28_27_r,temp_m4_28_27_i,`W4_real,`W4_imag,`W6_real,`W6_imag,`W10_real,`W10_imag);
butterfly butterfly987 (clk,temp_m4_20_19_r,temp_m4_20_19_i,temp_m4_20_27_r,temp_m4_20_27_i,temp_m4_28_19_r,temp_m4_28_19_i,temp_m4_28_27_r,temp_m4_28_27_i,temp_b4_20_19_r,temp_b4_20_19_i,temp_b4_20_27_r,temp_b4_20_27_i,temp_b4_28_19_r,temp_b4_28_19_i,temp_b4_28_27_r,temp_b4_28_27_i);
MULT MULT988 (clk,temp_b3_20_20_r,temp_b3_20_20_i,temp_b3_20_28_r,temp_b3_20_28_i,temp_b3_28_20_r,temp_b3_28_20_i,temp_b3_28_28_r,temp_b3_28_28_i,temp_m4_20_20_r,temp_m4_20_20_i,temp_m4_20_28_r,temp_m4_20_28_i,temp_m4_28_20_r,temp_m4_28_20_i,temp_m4_28_28_r,temp_m4_28_28_i,`W6_real,`W6_imag,`W6_real,`W6_imag,`W12_real,`W12_imag);
butterfly butterfly988 (clk,temp_m4_20_20_r,temp_m4_20_20_i,temp_m4_20_28_r,temp_m4_20_28_i,temp_m4_28_20_r,temp_m4_28_20_i,temp_m4_28_28_r,temp_m4_28_28_i,temp_b4_20_20_r,temp_b4_20_20_i,temp_b4_20_28_r,temp_b4_20_28_i,temp_b4_28_20_r,temp_b4_28_20_i,temp_b4_28_28_r,temp_b4_28_28_i);
MULT MULT989 (clk,temp_b3_20_21_r,temp_b3_20_21_i,temp_b3_20_29_r,temp_b3_20_29_i,temp_b3_28_21_r,temp_b3_28_21_i,temp_b3_28_29_r,temp_b3_28_29_i,temp_m4_20_21_r,temp_m4_20_21_i,temp_m4_20_29_r,temp_m4_20_29_i,temp_m4_28_21_r,temp_m4_28_21_i,temp_m4_28_29_r,temp_m4_28_29_i,`W8_real,`W8_imag,`W6_real,`W6_imag,`W14_real,`W14_imag);
butterfly butterfly989 (clk,temp_m4_20_21_r,temp_m4_20_21_i,temp_m4_20_29_r,temp_m4_20_29_i,temp_m4_28_21_r,temp_m4_28_21_i,temp_m4_28_29_r,temp_m4_28_29_i,temp_b4_20_21_r,temp_b4_20_21_i,temp_b4_20_29_r,temp_b4_20_29_i,temp_b4_28_21_r,temp_b4_28_21_i,temp_b4_28_29_r,temp_b4_28_29_i);
MULT MULT990 (clk,temp_b3_20_22_r,temp_b3_20_22_i,temp_b3_20_30_r,temp_b3_20_30_i,temp_b3_28_22_r,temp_b3_28_22_i,temp_b3_28_30_r,temp_b3_28_30_i,temp_m4_20_22_r,temp_m4_20_22_i,temp_m4_20_30_r,temp_m4_20_30_i,temp_m4_28_22_r,temp_m4_28_22_i,temp_m4_28_30_r,temp_m4_28_30_i,`W10_real,`W10_imag,`W6_real,`W6_imag,`W16_real,`W16_imag);
butterfly butterfly990 (clk,temp_m4_20_22_r,temp_m4_20_22_i,temp_m4_20_30_r,temp_m4_20_30_i,temp_m4_28_22_r,temp_m4_28_22_i,temp_m4_28_30_r,temp_m4_28_30_i,temp_b4_20_22_r,temp_b4_20_22_i,temp_b4_20_30_r,temp_b4_20_30_i,temp_b4_28_22_r,temp_b4_28_22_i,temp_b4_28_30_r,temp_b4_28_30_i);
MULT MULT991 (clk,temp_b3_20_23_r,temp_b3_20_23_i,temp_b3_20_31_r,temp_b3_20_31_i,temp_b3_28_23_r,temp_b3_28_23_i,temp_b3_28_31_r,temp_b3_28_31_i,temp_m4_20_23_r,temp_m4_20_23_i,temp_m4_20_31_r,temp_m4_20_31_i,temp_m4_28_23_r,temp_m4_28_23_i,temp_m4_28_31_r,temp_m4_28_31_i,`W12_real,`W12_imag,`W6_real,`W6_imag,`W18_real,`W18_imag);
butterfly butterfly991 (clk,temp_m4_20_23_r,temp_m4_20_23_i,temp_m4_20_31_r,temp_m4_20_31_i,temp_m4_28_23_r,temp_m4_28_23_i,temp_m4_28_31_r,temp_m4_28_31_i,temp_b4_20_23_r,temp_b4_20_23_i,temp_b4_20_31_r,temp_b4_20_31_i,temp_b4_28_23_r,temp_b4_28_23_i,temp_b4_28_31_r,temp_b4_28_31_i);
MULT MULT992 (clk,temp_b3_20_24_r,temp_b3_20_24_i,temp_b3_20_32_r,temp_b3_20_32_i,temp_b3_28_24_r,temp_b3_28_24_i,temp_b3_28_32_r,temp_b3_28_32_i,temp_m4_20_24_r,temp_m4_20_24_i,temp_m4_20_32_r,temp_m4_20_32_i,temp_m4_28_24_r,temp_m4_28_24_i,temp_m4_28_32_r,temp_m4_28_32_i,`W14_real,`W14_imag,`W6_real,`W6_imag,`W20_real,`W20_imag);
butterfly butterfly992 (clk,temp_m4_20_24_r,temp_m4_20_24_i,temp_m4_20_32_r,temp_m4_20_32_i,temp_m4_28_24_r,temp_m4_28_24_i,temp_m4_28_32_r,temp_m4_28_32_i,temp_b4_20_24_r,temp_b4_20_24_i,temp_b4_20_32_r,temp_b4_20_32_i,temp_b4_28_24_r,temp_b4_28_24_i,temp_b4_28_32_r,temp_b4_28_32_i);
MULT MULT993 (clk,temp_b3_21_17_r,temp_b3_21_17_i,temp_b3_21_25_r,temp_b3_21_25_i,temp_b3_29_17_r,temp_b3_29_17_i,temp_b3_29_25_r,temp_b3_29_25_i,temp_m4_21_17_r,temp_m4_21_17_i,temp_m4_21_25_r,temp_m4_21_25_i,temp_m4_29_17_r,temp_m4_29_17_i,temp_m4_29_25_r,temp_m4_29_25_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly993 (clk,temp_m4_21_17_r,temp_m4_21_17_i,temp_m4_21_25_r,temp_m4_21_25_i,temp_m4_29_17_r,temp_m4_29_17_i,temp_m4_29_25_r,temp_m4_29_25_i,temp_b4_21_17_r,temp_b4_21_17_i,temp_b4_21_25_r,temp_b4_21_25_i,temp_b4_29_17_r,temp_b4_29_17_i,temp_b4_29_25_r,temp_b4_29_25_i);
MULT MULT994 (clk,temp_b3_21_18_r,temp_b3_21_18_i,temp_b3_21_26_r,temp_b3_21_26_i,temp_b3_29_18_r,temp_b3_29_18_i,temp_b3_29_26_r,temp_b3_29_26_i,temp_m4_21_18_r,temp_m4_21_18_i,temp_m4_21_26_r,temp_m4_21_26_i,temp_m4_29_18_r,temp_m4_29_18_i,temp_m4_29_26_r,temp_m4_29_26_i,`W2_real,`W2_imag,`W8_real,`W8_imag,`W10_real,`W10_imag);
butterfly butterfly994 (clk,temp_m4_21_18_r,temp_m4_21_18_i,temp_m4_21_26_r,temp_m4_21_26_i,temp_m4_29_18_r,temp_m4_29_18_i,temp_m4_29_26_r,temp_m4_29_26_i,temp_b4_21_18_r,temp_b4_21_18_i,temp_b4_21_26_r,temp_b4_21_26_i,temp_b4_29_18_r,temp_b4_29_18_i,temp_b4_29_26_r,temp_b4_29_26_i);
MULT MULT995 (clk,temp_b3_21_19_r,temp_b3_21_19_i,temp_b3_21_27_r,temp_b3_21_27_i,temp_b3_29_19_r,temp_b3_29_19_i,temp_b3_29_27_r,temp_b3_29_27_i,temp_m4_21_19_r,temp_m4_21_19_i,temp_m4_21_27_r,temp_m4_21_27_i,temp_m4_29_19_r,temp_m4_29_19_i,temp_m4_29_27_r,temp_m4_29_27_i,`W4_real,`W4_imag,`W8_real,`W8_imag,`W12_real,`W12_imag);
butterfly butterfly995 (clk,temp_m4_21_19_r,temp_m4_21_19_i,temp_m4_21_27_r,temp_m4_21_27_i,temp_m4_29_19_r,temp_m4_29_19_i,temp_m4_29_27_r,temp_m4_29_27_i,temp_b4_21_19_r,temp_b4_21_19_i,temp_b4_21_27_r,temp_b4_21_27_i,temp_b4_29_19_r,temp_b4_29_19_i,temp_b4_29_27_r,temp_b4_29_27_i);
MULT MULT996 (clk,temp_b3_21_20_r,temp_b3_21_20_i,temp_b3_21_28_r,temp_b3_21_28_i,temp_b3_29_20_r,temp_b3_29_20_i,temp_b3_29_28_r,temp_b3_29_28_i,temp_m4_21_20_r,temp_m4_21_20_i,temp_m4_21_28_r,temp_m4_21_28_i,temp_m4_29_20_r,temp_m4_29_20_i,temp_m4_29_28_r,temp_m4_29_28_i,`W6_real,`W6_imag,`W8_real,`W8_imag,`W14_real,`W14_imag);
butterfly butterfly996 (clk,temp_m4_21_20_r,temp_m4_21_20_i,temp_m4_21_28_r,temp_m4_21_28_i,temp_m4_29_20_r,temp_m4_29_20_i,temp_m4_29_28_r,temp_m4_29_28_i,temp_b4_21_20_r,temp_b4_21_20_i,temp_b4_21_28_r,temp_b4_21_28_i,temp_b4_29_20_r,temp_b4_29_20_i,temp_b4_29_28_r,temp_b4_29_28_i);
MULT MULT997 (clk,temp_b3_21_21_r,temp_b3_21_21_i,temp_b3_21_29_r,temp_b3_21_29_i,temp_b3_29_21_r,temp_b3_29_21_i,temp_b3_29_29_r,temp_b3_29_29_i,temp_m4_21_21_r,temp_m4_21_21_i,temp_m4_21_29_r,temp_m4_21_29_i,temp_m4_29_21_r,temp_m4_29_21_i,temp_m4_29_29_r,temp_m4_29_29_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly997 (clk,temp_m4_21_21_r,temp_m4_21_21_i,temp_m4_21_29_r,temp_m4_21_29_i,temp_m4_29_21_r,temp_m4_29_21_i,temp_m4_29_29_r,temp_m4_29_29_i,temp_b4_21_21_r,temp_b4_21_21_i,temp_b4_21_29_r,temp_b4_21_29_i,temp_b4_29_21_r,temp_b4_29_21_i,temp_b4_29_29_r,temp_b4_29_29_i);
MULT MULT998 (clk,temp_b3_21_22_r,temp_b3_21_22_i,temp_b3_21_30_r,temp_b3_21_30_i,temp_b3_29_22_r,temp_b3_29_22_i,temp_b3_29_30_r,temp_b3_29_30_i,temp_m4_21_22_r,temp_m4_21_22_i,temp_m4_21_30_r,temp_m4_21_30_i,temp_m4_29_22_r,temp_m4_29_22_i,temp_m4_29_30_r,temp_m4_29_30_i,`W10_real,`W10_imag,`W8_real,`W8_imag,`W18_real,`W18_imag);
butterfly butterfly998 (clk,temp_m4_21_22_r,temp_m4_21_22_i,temp_m4_21_30_r,temp_m4_21_30_i,temp_m4_29_22_r,temp_m4_29_22_i,temp_m4_29_30_r,temp_m4_29_30_i,temp_b4_21_22_r,temp_b4_21_22_i,temp_b4_21_30_r,temp_b4_21_30_i,temp_b4_29_22_r,temp_b4_29_22_i,temp_b4_29_30_r,temp_b4_29_30_i);
MULT MULT999 (clk,temp_b3_21_23_r,temp_b3_21_23_i,temp_b3_21_31_r,temp_b3_21_31_i,temp_b3_29_23_r,temp_b3_29_23_i,temp_b3_29_31_r,temp_b3_29_31_i,temp_m4_21_23_r,temp_m4_21_23_i,temp_m4_21_31_r,temp_m4_21_31_i,temp_m4_29_23_r,temp_m4_29_23_i,temp_m4_29_31_r,temp_m4_29_31_i,`W12_real,`W12_imag,`W8_real,`W8_imag,`W20_real,`W20_imag);
butterfly butterfly999 (clk,temp_m4_21_23_r,temp_m4_21_23_i,temp_m4_21_31_r,temp_m4_21_31_i,temp_m4_29_23_r,temp_m4_29_23_i,temp_m4_29_31_r,temp_m4_29_31_i,temp_b4_21_23_r,temp_b4_21_23_i,temp_b4_21_31_r,temp_b4_21_31_i,temp_b4_29_23_r,temp_b4_29_23_i,temp_b4_29_31_r,temp_b4_29_31_i);
MULT MULT1000 (clk,temp_b3_21_24_r,temp_b3_21_24_i,temp_b3_21_32_r,temp_b3_21_32_i,temp_b3_29_24_r,temp_b3_29_24_i,temp_b3_29_32_r,temp_b3_29_32_i,temp_m4_21_24_r,temp_m4_21_24_i,temp_m4_21_32_r,temp_m4_21_32_i,temp_m4_29_24_r,temp_m4_29_24_i,temp_m4_29_32_r,temp_m4_29_32_i,`W14_real,`W14_imag,`W8_real,`W8_imag,`W22_real,`W22_imag);
butterfly butterfly1000 (clk,temp_m4_21_24_r,temp_m4_21_24_i,temp_m4_21_32_r,temp_m4_21_32_i,temp_m4_29_24_r,temp_m4_29_24_i,temp_m4_29_32_r,temp_m4_29_32_i,temp_b4_21_24_r,temp_b4_21_24_i,temp_b4_21_32_r,temp_b4_21_32_i,temp_b4_29_24_r,temp_b4_29_24_i,temp_b4_29_32_r,temp_b4_29_32_i);
MULT MULT1001 (clk,temp_b3_22_17_r,temp_b3_22_17_i,temp_b3_22_25_r,temp_b3_22_25_i,temp_b3_30_17_r,temp_b3_30_17_i,temp_b3_30_25_r,temp_b3_30_25_i,temp_m4_22_17_r,temp_m4_22_17_i,temp_m4_22_25_r,temp_m4_22_25_i,temp_m4_30_17_r,temp_m4_30_17_i,temp_m4_30_25_r,temp_m4_30_25_i,`W0_real,`W0_imag,`W10_real,`W10_imag,`W10_real,`W10_imag);
butterfly butterfly1001 (clk,temp_m4_22_17_r,temp_m4_22_17_i,temp_m4_22_25_r,temp_m4_22_25_i,temp_m4_30_17_r,temp_m4_30_17_i,temp_m4_30_25_r,temp_m4_30_25_i,temp_b4_22_17_r,temp_b4_22_17_i,temp_b4_22_25_r,temp_b4_22_25_i,temp_b4_30_17_r,temp_b4_30_17_i,temp_b4_30_25_r,temp_b4_30_25_i);
MULT MULT1002 (clk,temp_b3_22_18_r,temp_b3_22_18_i,temp_b3_22_26_r,temp_b3_22_26_i,temp_b3_30_18_r,temp_b3_30_18_i,temp_b3_30_26_r,temp_b3_30_26_i,temp_m4_22_18_r,temp_m4_22_18_i,temp_m4_22_26_r,temp_m4_22_26_i,temp_m4_30_18_r,temp_m4_30_18_i,temp_m4_30_26_r,temp_m4_30_26_i,`W2_real,`W2_imag,`W10_real,`W10_imag,`W12_real,`W12_imag);
butterfly butterfly1002 (clk,temp_m4_22_18_r,temp_m4_22_18_i,temp_m4_22_26_r,temp_m4_22_26_i,temp_m4_30_18_r,temp_m4_30_18_i,temp_m4_30_26_r,temp_m4_30_26_i,temp_b4_22_18_r,temp_b4_22_18_i,temp_b4_22_26_r,temp_b4_22_26_i,temp_b4_30_18_r,temp_b4_30_18_i,temp_b4_30_26_r,temp_b4_30_26_i);
MULT MULT1003 (clk,temp_b3_22_19_r,temp_b3_22_19_i,temp_b3_22_27_r,temp_b3_22_27_i,temp_b3_30_19_r,temp_b3_30_19_i,temp_b3_30_27_r,temp_b3_30_27_i,temp_m4_22_19_r,temp_m4_22_19_i,temp_m4_22_27_r,temp_m4_22_27_i,temp_m4_30_19_r,temp_m4_30_19_i,temp_m4_30_27_r,temp_m4_30_27_i,`W4_real,`W4_imag,`W10_real,`W10_imag,`W14_real,`W14_imag);
butterfly butterfly1003 (clk,temp_m4_22_19_r,temp_m4_22_19_i,temp_m4_22_27_r,temp_m4_22_27_i,temp_m4_30_19_r,temp_m4_30_19_i,temp_m4_30_27_r,temp_m4_30_27_i,temp_b4_22_19_r,temp_b4_22_19_i,temp_b4_22_27_r,temp_b4_22_27_i,temp_b4_30_19_r,temp_b4_30_19_i,temp_b4_30_27_r,temp_b4_30_27_i);
MULT MULT1004 (clk,temp_b3_22_20_r,temp_b3_22_20_i,temp_b3_22_28_r,temp_b3_22_28_i,temp_b3_30_20_r,temp_b3_30_20_i,temp_b3_30_28_r,temp_b3_30_28_i,temp_m4_22_20_r,temp_m4_22_20_i,temp_m4_22_28_r,temp_m4_22_28_i,temp_m4_30_20_r,temp_m4_30_20_i,temp_m4_30_28_r,temp_m4_30_28_i,`W6_real,`W6_imag,`W10_real,`W10_imag,`W16_real,`W16_imag);
butterfly butterfly1004 (clk,temp_m4_22_20_r,temp_m4_22_20_i,temp_m4_22_28_r,temp_m4_22_28_i,temp_m4_30_20_r,temp_m4_30_20_i,temp_m4_30_28_r,temp_m4_30_28_i,temp_b4_22_20_r,temp_b4_22_20_i,temp_b4_22_28_r,temp_b4_22_28_i,temp_b4_30_20_r,temp_b4_30_20_i,temp_b4_30_28_r,temp_b4_30_28_i);
MULT MULT1005 (clk,temp_b3_22_21_r,temp_b3_22_21_i,temp_b3_22_29_r,temp_b3_22_29_i,temp_b3_30_21_r,temp_b3_30_21_i,temp_b3_30_29_r,temp_b3_30_29_i,temp_m4_22_21_r,temp_m4_22_21_i,temp_m4_22_29_r,temp_m4_22_29_i,temp_m4_30_21_r,temp_m4_30_21_i,temp_m4_30_29_r,temp_m4_30_29_i,`W8_real,`W8_imag,`W10_real,`W10_imag,`W18_real,`W18_imag);
butterfly butterfly1005 (clk,temp_m4_22_21_r,temp_m4_22_21_i,temp_m4_22_29_r,temp_m4_22_29_i,temp_m4_30_21_r,temp_m4_30_21_i,temp_m4_30_29_r,temp_m4_30_29_i,temp_b4_22_21_r,temp_b4_22_21_i,temp_b4_22_29_r,temp_b4_22_29_i,temp_b4_30_21_r,temp_b4_30_21_i,temp_b4_30_29_r,temp_b4_30_29_i);
MULT MULT1006 (clk,temp_b3_22_22_r,temp_b3_22_22_i,temp_b3_22_30_r,temp_b3_22_30_i,temp_b3_30_22_r,temp_b3_30_22_i,temp_b3_30_30_r,temp_b3_30_30_i,temp_m4_22_22_r,temp_m4_22_22_i,temp_m4_22_30_r,temp_m4_22_30_i,temp_m4_30_22_r,temp_m4_30_22_i,temp_m4_30_30_r,temp_m4_30_30_i,`W10_real,`W10_imag,`W10_real,`W10_imag,`W20_real,`W20_imag);
butterfly butterfly1006 (clk,temp_m4_22_22_r,temp_m4_22_22_i,temp_m4_22_30_r,temp_m4_22_30_i,temp_m4_30_22_r,temp_m4_30_22_i,temp_m4_30_30_r,temp_m4_30_30_i,temp_b4_22_22_r,temp_b4_22_22_i,temp_b4_22_30_r,temp_b4_22_30_i,temp_b4_30_22_r,temp_b4_30_22_i,temp_b4_30_30_r,temp_b4_30_30_i);
MULT MULT1007 (clk,temp_b3_22_23_r,temp_b3_22_23_i,temp_b3_22_31_r,temp_b3_22_31_i,temp_b3_30_23_r,temp_b3_30_23_i,temp_b3_30_31_r,temp_b3_30_31_i,temp_m4_22_23_r,temp_m4_22_23_i,temp_m4_22_31_r,temp_m4_22_31_i,temp_m4_30_23_r,temp_m4_30_23_i,temp_m4_30_31_r,temp_m4_30_31_i,`W12_real,`W12_imag,`W10_real,`W10_imag,`W22_real,`W22_imag);
butterfly butterfly1007 (clk,temp_m4_22_23_r,temp_m4_22_23_i,temp_m4_22_31_r,temp_m4_22_31_i,temp_m4_30_23_r,temp_m4_30_23_i,temp_m4_30_31_r,temp_m4_30_31_i,temp_b4_22_23_r,temp_b4_22_23_i,temp_b4_22_31_r,temp_b4_22_31_i,temp_b4_30_23_r,temp_b4_30_23_i,temp_b4_30_31_r,temp_b4_30_31_i);
MULT MULT1008 (clk,temp_b3_22_24_r,temp_b3_22_24_i,temp_b3_22_32_r,temp_b3_22_32_i,temp_b3_30_24_r,temp_b3_30_24_i,temp_b3_30_32_r,temp_b3_30_32_i,temp_m4_22_24_r,temp_m4_22_24_i,temp_m4_22_32_r,temp_m4_22_32_i,temp_m4_30_24_r,temp_m4_30_24_i,temp_m4_30_32_r,temp_m4_30_32_i,`W14_real,`W14_imag,`W10_real,`W10_imag,`W24_real,`W24_imag);
butterfly butterfly1008 (clk,temp_m4_22_24_r,temp_m4_22_24_i,temp_m4_22_32_r,temp_m4_22_32_i,temp_m4_30_24_r,temp_m4_30_24_i,temp_m4_30_32_r,temp_m4_30_32_i,temp_b4_22_24_r,temp_b4_22_24_i,temp_b4_22_32_r,temp_b4_22_32_i,temp_b4_30_24_r,temp_b4_30_24_i,temp_b4_30_32_r,temp_b4_30_32_i);
MULT MULT1009 (clk,temp_b3_23_17_r,temp_b3_23_17_i,temp_b3_23_25_r,temp_b3_23_25_i,temp_b3_31_17_r,temp_b3_31_17_i,temp_b3_31_25_r,temp_b3_31_25_i,temp_m4_23_17_r,temp_m4_23_17_i,temp_m4_23_25_r,temp_m4_23_25_i,temp_m4_31_17_r,temp_m4_31_17_i,temp_m4_31_25_r,temp_m4_31_25_i,`W0_real,`W0_imag,`W12_real,`W12_imag,`W12_real,`W12_imag);
butterfly butterfly1009 (clk,temp_m4_23_17_r,temp_m4_23_17_i,temp_m4_23_25_r,temp_m4_23_25_i,temp_m4_31_17_r,temp_m4_31_17_i,temp_m4_31_25_r,temp_m4_31_25_i,temp_b4_23_17_r,temp_b4_23_17_i,temp_b4_23_25_r,temp_b4_23_25_i,temp_b4_31_17_r,temp_b4_31_17_i,temp_b4_31_25_r,temp_b4_31_25_i);
MULT MULT1010 (clk,temp_b3_23_18_r,temp_b3_23_18_i,temp_b3_23_26_r,temp_b3_23_26_i,temp_b3_31_18_r,temp_b3_31_18_i,temp_b3_31_26_r,temp_b3_31_26_i,temp_m4_23_18_r,temp_m4_23_18_i,temp_m4_23_26_r,temp_m4_23_26_i,temp_m4_31_18_r,temp_m4_31_18_i,temp_m4_31_26_r,temp_m4_31_26_i,`W2_real,`W2_imag,`W12_real,`W12_imag,`W14_real,`W14_imag);
butterfly butterfly1010 (clk,temp_m4_23_18_r,temp_m4_23_18_i,temp_m4_23_26_r,temp_m4_23_26_i,temp_m4_31_18_r,temp_m4_31_18_i,temp_m4_31_26_r,temp_m4_31_26_i,temp_b4_23_18_r,temp_b4_23_18_i,temp_b4_23_26_r,temp_b4_23_26_i,temp_b4_31_18_r,temp_b4_31_18_i,temp_b4_31_26_r,temp_b4_31_26_i);
MULT MULT1011 (clk,temp_b3_23_19_r,temp_b3_23_19_i,temp_b3_23_27_r,temp_b3_23_27_i,temp_b3_31_19_r,temp_b3_31_19_i,temp_b3_31_27_r,temp_b3_31_27_i,temp_m4_23_19_r,temp_m4_23_19_i,temp_m4_23_27_r,temp_m4_23_27_i,temp_m4_31_19_r,temp_m4_31_19_i,temp_m4_31_27_r,temp_m4_31_27_i,`W4_real,`W4_imag,`W12_real,`W12_imag,`W16_real,`W16_imag);
butterfly butterfly1011 (clk,temp_m4_23_19_r,temp_m4_23_19_i,temp_m4_23_27_r,temp_m4_23_27_i,temp_m4_31_19_r,temp_m4_31_19_i,temp_m4_31_27_r,temp_m4_31_27_i,temp_b4_23_19_r,temp_b4_23_19_i,temp_b4_23_27_r,temp_b4_23_27_i,temp_b4_31_19_r,temp_b4_31_19_i,temp_b4_31_27_r,temp_b4_31_27_i);
MULT MULT1012 (clk,temp_b3_23_20_r,temp_b3_23_20_i,temp_b3_23_28_r,temp_b3_23_28_i,temp_b3_31_20_r,temp_b3_31_20_i,temp_b3_31_28_r,temp_b3_31_28_i,temp_m4_23_20_r,temp_m4_23_20_i,temp_m4_23_28_r,temp_m4_23_28_i,temp_m4_31_20_r,temp_m4_31_20_i,temp_m4_31_28_r,temp_m4_31_28_i,`W6_real,`W6_imag,`W12_real,`W12_imag,`W18_real,`W18_imag);
butterfly butterfly1012 (clk,temp_m4_23_20_r,temp_m4_23_20_i,temp_m4_23_28_r,temp_m4_23_28_i,temp_m4_31_20_r,temp_m4_31_20_i,temp_m4_31_28_r,temp_m4_31_28_i,temp_b4_23_20_r,temp_b4_23_20_i,temp_b4_23_28_r,temp_b4_23_28_i,temp_b4_31_20_r,temp_b4_31_20_i,temp_b4_31_28_r,temp_b4_31_28_i);
MULT MULT1013 (clk,temp_b3_23_21_r,temp_b3_23_21_i,temp_b3_23_29_r,temp_b3_23_29_i,temp_b3_31_21_r,temp_b3_31_21_i,temp_b3_31_29_r,temp_b3_31_29_i,temp_m4_23_21_r,temp_m4_23_21_i,temp_m4_23_29_r,temp_m4_23_29_i,temp_m4_31_21_r,temp_m4_31_21_i,temp_m4_31_29_r,temp_m4_31_29_i,`W8_real,`W8_imag,`W12_real,`W12_imag,`W20_real,`W20_imag);
butterfly butterfly1013 (clk,temp_m4_23_21_r,temp_m4_23_21_i,temp_m4_23_29_r,temp_m4_23_29_i,temp_m4_31_21_r,temp_m4_31_21_i,temp_m4_31_29_r,temp_m4_31_29_i,temp_b4_23_21_r,temp_b4_23_21_i,temp_b4_23_29_r,temp_b4_23_29_i,temp_b4_31_21_r,temp_b4_31_21_i,temp_b4_31_29_r,temp_b4_31_29_i);
MULT MULT1014 (clk,temp_b3_23_22_r,temp_b3_23_22_i,temp_b3_23_30_r,temp_b3_23_30_i,temp_b3_31_22_r,temp_b3_31_22_i,temp_b3_31_30_r,temp_b3_31_30_i,temp_m4_23_22_r,temp_m4_23_22_i,temp_m4_23_30_r,temp_m4_23_30_i,temp_m4_31_22_r,temp_m4_31_22_i,temp_m4_31_30_r,temp_m4_31_30_i,`W10_real,`W10_imag,`W12_real,`W12_imag,`W22_real,`W22_imag);
butterfly butterfly1014 (clk,temp_m4_23_22_r,temp_m4_23_22_i,temp_m4_23_30_r,temp_m4_23_30_i,temp_m4_31_22_r,temp_m4_31_22_i,temp_m4_31_30_r,temp_m4_31_30_i,temp_b4_23_22_r,temp_b4_23_22_i,temp_b4_23_30_r,temp_b4_23_30_i,temp_b4_31_22_r,temp_b4_31_22_i,temp_b4_31_30_r,temp_b4_31_30_i);
MULT MULT1015 (clk,temp_b3_23_23_r,temp_b3_23_23_i,temp_b3_23_31_r,temp_b3_23_31_i,temp_b3_31_23_r,temp_b3_31_23_i,temp_b3_31_31_r,temp_b3_31_31_i,temp_m4_23_23_r,temp_m4_23_23_i,temp_m4_23_31_r,temp_m4_23_31_i,temp_m4_31_23_r,temp_m4_31_23_i,temp_m4_31_31_r,temp_m4_31_31_i,`W12_real,`W12_imag,`W12_real,`W12_imag,`W24_real,`W24_imag);
butterfly butterfly1015 (clk,temp_m4_23_23_r,temp_m4_23_23_i,temp_m4_23_31_r,temp_m4_23_31_i,temp_m4_31_23_r,temp_m4_31_23_i,temp_m4_31_31_r,temp_m4_31_31_i,temp_b4_23_23_r,temp_b4_23_23_i,temp_b4_23_31_r,temp_b4_23_31_i,temp_b4_31_23_r,temp_b4_31_23_i,temp_b4_31_31_r,temp_b4_31_31_i);
MULT MULT1016 (clk,temp_b3_23_24_r,temp_b3_23_24_i,temp_b3_23_32_r,temp_b3_23_32_i,temp_b3_31_24_r,temp_b3_31_24_i,temp_b3_31_32_r,temp_b3_31_32_i,temp_m4_23_24_r,temp_m4_23_24_i,temp_m4_23_32_r,temp_m4_23_32_i,temp_m4_31_24_r,temp_m4_31_24_i,temp_m4_31_32_r,temp_m4_31_32_i,`W14_real,`W14_imag,`W12_real,`W12_imag,`W26_real,`W26_imag);
butterfly butterfly1016 (clk,temp_m4_23_24_r,temp_m4_23_24_i,temp_m4_23_32_r,temp_m4_23_32_i,temp_m4_31_24_r,temp_m4_31_24_i,temp_m4_31_32_r,temp_m4_31_32_i,temp_b4_23_24_r,temp_b4_23_24_i,temp_b4_23_32_r,temp_b4_23_32_i,temp_b4_31_24_r,temp_b4_31_24_i,temp_b4_31_32_r,temp_b4_31_32_i);
MULT MULT1017 (clk,temp_b3_24_17_r,temp_b3_24_17_i,temp_b3_24_25_r,temp_b3_24_25_i,temp_b3_32_17_r,temp_b3_32_17_i,temp_b3_32_25_r,temp_b3_32_25_i,temp_m4_24_17_r,temp_m4_24_17_i,temp_m4_24_25_r,temp_m4_24_25_i,temp_m4_32_17_r,temp_m4_32_17_i,temp_m4_32_25_r,temp_m4_32_25_i,`W0_real,`W0_imag,`W14_real,`W14_imag,`W14_real,`W14_imag);
butterfly butterfly1017 (clk,temp_m4_24_17_r,temp_m4_24_17_i,temp_m4_24_25_r,temp_m4_24_25_i,temp_m4_32_17_r,temp_m4_32_17_i,temp_m4_32_25_r,temp_m4_32_25_i,temp_b4_24_17_r,temp_b4_24_17_i,temp_b4_24_25_r,temp_b4_24_25_i,temp_b4_32_17_r,temp_b4_32_17_i,temp_b4_32_25_r,temp_b4_32_25_i);
MULT MULT1018 (clk,temp_b3_24_18_r,temp_b3_24_18_i,temp_b3_24_26_r,temp_b3_24_26_i,temp_b3_32_18_r,temp_b3_32_18_i,temp_b3_32_26_r,temp_b3_32_26_i,temp_m4_24_18_r,temp_m4_24_18_i,temp_m4_24_26_r,temp_m4_24_26_i,temp_m4_32_18_r,temp_m4_32_18_i,temp_m4_32_26_r,temp_m4_32_26_i,`W2_real,`W2_imag,`W14_real,`W14_imag,`W16_real,`W16_imag);
butterfly butterfly1018 (clk,temp_m4_24_18_r,temp_m4_24_18_i,temp_m4_24_26_r,temp_m4_24_26_i,temp_m4_32_18_r,temp_m4_32_18_i,temp_m4_32_26_r,temp_m4_32_26_i,temp_b4_24_18_r,temp_b4_24_18_i,temp_b4_24_26_r,temp_b4_24_26_i,temp_b4_32_18_r,temp_b4_32_18_i,temp_b4_32_26_r,temp_b4_32_26_i);
MULT MULT1019 (clk,temp_b3_24_19_r,temp_b3_24_19_i,temp_b3_24_27_r,temp_b3_24_27_i,temp_b3_32_19_r,temp_b3_32_19_i,temp_b3_32_27_r,temp_b3_32_27_i,temp_m4_24_19_r,temp_m4_24_19_i,temp_m4_24_27_r,temp_m4_24_27_i,temp_m4_32_19_r,temp_m4_32_19_i,temp_m4_32_27_r,temp_m4_32_27_i,`W4_real,`W4_imag,`W14_real,`W14_imag,`W18_real,`W18_imag);
butterfly butterfly1019 (clk,temp_m4_24_19_r,temp_m4_24_19_i,temp_m4_24_27_r,temp_m4_24_27_i,temp_m4_32_19_r,temp_m4_32_19_i,temp_m4_32_27_r,temp_m4_32_27_i,temp_b4_24_19_r,temp_b4_24_19_i,temp_b4_24_27_r,temp_b4_24_27_i,temp_b4_32_19_r,temp_b4_32_19_i,temp_b4_32_27_r,temp_b4_32_27_i);
MULT MULT1020 (clk,temp_b3_24_20_r,temp_b3_24_20_i,temp_b3_24_28_r,temp_b3_24_28_i,temp_b3_32_20_r,temp_b3_32_20_i,temp_b3_32_28_r,temp_b3_32_28_i,temp_m4_24_20_r,temp_m4_24_20_i,temp_m4_24_28_r,temp_m4_24_28_i,temp_m4_32_20_r,temp_m4_32_20_i,temp_m4_32_28_r,temp_m4_32_28_i,`W6_real,`W6_imag,`W14_real,`W14_imag,`W20_real,`W20_imag);
butterfly butterfly1020 (clk,temp_m4_24_20_r,temp_m4_24_20_i,temp_m4_24_28_r,temp_m4_24_28_i,temp_m4_32_20_r,temp_m4_32_20_i,temp_m4_32_28_r,temp_m4_32_28_i,temp_b4_24_20_r,temp_b4_24_20_i,temp_b4_24_28_r,temp_b4_24_28_i,temp_b4_32_20_r,temp_b4_32_20_i,temp_b4_32_28_r,temp_b4_32_28_i);
MULT MULT1021 (clk,temp_b3_24_21_r,temp_b3_24_21_i,temp_b3_24_29_r,temp_b3_24_29_i,temp_b3_32_21_r,temp_b3_32_21_i,temp_b3_32_29_r,temp_b3_32_29_i,temp_m4_24_21_r,temp_m4_24_21_i,temp_m4_24_29_r,temp_m4_24_29_i,temp_m4_32_21_r,temp_m4_32_21_i,temp_m4_32_29_r,temp_m4_32_29_i,`W8_real,`W8_imag,`W14_real,`W14_imag,`W22_real,`W22_imag);
butterfly butterfly1021 (clk,temp_m4_24_21_r,temp_m4_24_21_i,temp_m4_24_29_r,temp_m4_24_29_i,temp_m4_32_21_r,temp_m4_32_21_i,temp_m4_32_29_r,temp_m4_32_29_i,temp_b4_24_21_r,temp_b4_24_21_i,temp_b4_24_29_r,temp_b4_24_29_i,temp_b4_32_21_r,temp_b4_32_21_i,temp_b4_32_29_r,temp_b4_32_29_i);
MULT MULT1022 (clk,temp_b3_24_22_r,temp_b3_24_22_i,temp_b3_24_30_r,temp_b3_24_30_i,temp_b3_32_22_r,temp_b3_32_22_i,temp_b3_32_30_r,temp_b3_32_30_i,temp_m4_24_22_r,temp_m4_24_22_i,temp_m4_24_30_r,temp_m4_24_30_i,temp_m4_32_22_r,temp_m4_32_22_i,temp_m4_32_30_r,temp_m4_32_30_i,`W10_real,`W10_imag,`W14_real,`W14_imag,`W24_real,`W24_imag);
butterfly butterfly1022 (clk,temp_m4_24_22_r,temp_m4_24_22_i,temp_m4_24_30_r,temp_m4_24_30_i,temp_m4_32_22_r,temp_m4_32_22_i,temp_m4_32_30_r,temp_m4_32_30_i,temp_b4_24_22_r,temp_b4_24_22_i,temp_b4_24_30_r,temp_b4_24_30_i,temp_b4_32_22_r,temp_b4_32_22_i,temp_b4_32_30_r,temp_b4_32_30_i);
MULT MULT1023 (clk,temp_b3_24_23_r,temp_b3_24_23_i,temp_b3_24_31_r,temp_b3_24_31_i,temp_b3_32_23_r,temp_b3_32_23_i,temp_b3_32_31_r,temp_b3_32_31_i,temp_m4_24_23_r,temp_m4_24_23_i,temp_m4_24_31_r,temp_m4_24_31_i,temp_m4_32_23_r,temp_m4_32_23_i,temp_m4_32_31_r,temp_m4_32_31_i,`W12_real,`W12_imag,`W14_real,`W14_imag,`W26_real,`W26_imag);
butterfly butterfly1023 (clk,temp_m4_24_23_r,temp_m4_24_23_i,temp_m4_24_31_r,temp_m4_24_31_i,temp_m4_32_23_r,temp_m4_32_23_i,temp_m4_32_31_r,temp_m4_32_31_i,temp_b4_24_23_r,temp_b4_24_23_i,temp_b4_24_31_r,temp_b4_24_31_i,temp_b4_32_23_r,temp_b4_32_23_i,temp_b4_32_31_r,temp_b4_32_31_i);
MULT MULT1024 (clk,temp_b3_24_24_r,temp_b3_24_24_i,temp_b3_24_32_r,temp_b3_24_32_i,temp_b3_32_24_r,temp_b3_32_24_i,temp_b3_32_32_r,temp_b3_32_32_i,temp_m4_24_24_r,temp_m4_24_24_i,temp_m4_24_32_r,temp_m4_24_32_i,temp_m4_32_24_r,temp_m4_32_24_i,temp_m4_32_32_r,temp_m4_32_32_i,`W14_real,`W14_imag,`W14_real,`W14_imag,`W28_real,`W28_imag);
butterfly butterfly1024 (clk,temp_m4_24_24_r,temp_m4_24_24_i,temp_m4_24_32_r,temp_m4_24_32_i,temp_m4_32_24_r,temp_m4_32_24_i,temp_m4_32_32_r,temp_m4_32_32_i,temp_b4_24_24_r,temp_b4_24_24_i,temp_b4_24_32_r,temp_b4_24_32_i,temp_b4_32_24_r,temp_b4_32_24_i,temp_b4_32_32_r,temp_b4_32_32_i);
MULT MULT1025 (clk,temp_b4_1_1_r,temp_b4_1_1_i,temp_b4_1_17_r,temp_b4_1_17_i,temp_b4_17_1_r,temp_b4_17_1_i,temp_b4_17_17_r,temp_b4_17_17_i,temp_m5_1_1_r,temp_m5_1_1_i,temp_m5_1_17_r,temp_m5_1_17_i,temp_m5_17_1_r,temp_m5_17_1_i,temp_m5_17_17_r,temp_m5_17_17_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly1025 (clk,temp_m5_1_1_r,temp_m5_1_1_i,temp_m5_1_17_r,temp_m5_1_17_i,temp_m5_17_1_r,temp_m5_17_1_i,temp_m5_17_17_r,temp_m5_17_17_i,temp_b5_1_1_r,temp_b5_1_1_i,temp_b5_1_17_r,temp_b5_1_17_i,temp_b5_17_1_r,temp_b5_17_1_i,temp_b5_17_17_r,temp_b5_17_17_i);
MULT MULT1026 (clk,temp_b4_1_2_r,temp_b4_1_2_i,temp_b4_1_18_r,temp_b4_1_18_i,temp_b4_17_2_r,temp_b4_17_2_i,temp_b4_17_18_r,temp_b4_17_18_i,temp_m5_1_2_r,temp_m5_1_2_i,temp_m5_1_18_r,temp_m5_1_18_i,temp_m5_17_2_r,temp_m5_17_2_i,temp_m5_17_18_r,temp_m5_17_18_i,`W1_real,`W1_imag,`W0_real,`W0_imag,`W1_real,`W1_imag);
butterfly butterfly1026 (clk,temp_m5_1_2_r,temp_m5_1_2_i,temp_m5_1_18_r,temp_m5_1_18_i,temp_m5_17_2_r,temp_m5_17_2_i,temp_m5_17_18_r,temp_m5_17_18_i,temp_b5_1_2_r,temp_b5_1_2_i,temp_b5_1_18_r,temp_b5_1_18_i,temp_b5_17_2_r,temp_b5_17_2_i,temp_b5_17_18_r,temp_b5_17_18_i);
MULT MULT1027 (clk,temp_b4_1_3_r,temp_b4_1_3_i,temp_b4_1_19_r,temp_b4_1_19_i,temp_b4_17_3_r,temp_b4_17_3_i,temp_b4_17_19_r,temp_b4_17_19_i,temp_m5_1_3_r,temp_m5_1_3_i,temp_m5_1_19_r,temp_m5_1_19_i,temp_m5_17_3_r,temp_m5_17_3_i,temp_m5_17_19_r,temp_m5_17_19_i,`W2_real,`W2_imag,`W0_real,`W0_imag,`W2_real,`W2_imag);
butterfly butterfly1027 (clk,temp_m5_1_3_r,temp_m5_1_3_i,temp_m5_1_19_r,temp_m5_1_19_i,temp_m5_17_3_r,temp_m5_17_3_i,temp_m5_17_19_r,temp_m5_17_19_i,temp_b5_1_3_r,temp_b5_1_3_i,temp_b5_1_19_r,temp_b5_1_19_i,temp_b5_17_3_r,temp_b5_17_3_i,temp_b5_17_19_r,temp_b5_17_19_i);
MULT MULT1028 (clk,temp_b4_1_4_r,temp_b4_1_4_i,temp_b4_1_20_r,temp_b4_1_20_i,temp_b4_17_4_r,temp_b4_17_4_i,temp_b4_17_20_r,temp_b4_17_20_i,temp_m5_1_4_r,temp_m5_1_4_i,temp_m5_1_20_r,temp_m5_1_20_i,temp_m5_17_4_r,temp_m5_17_4_i,temp_m5_17_20_r,temp_m5_17_20_i,`W3_real,`W3_imag,`W0_real,`W0_imag,`W3_real,`W3_imag);
butterfly butterfly1028 (clk,temp_m5_1_4_r,temp_m5_1_4_i,temp_m5_1_20_r,temp_m5_1_20_i,temp_m5_17_4_r,temp_m5_17_4_i,temp_m5_17_20_r,temp_m5_17_20_i,temp_b5_1_4_r,temp_b5_1_4_i,temp_b5_1_20_r,temp_b5_1_20_i,temp_b5_17_4_r,temp_b5_17_4_i,temp_b5_17_20_r,temp_b5_17_20_i);
MULT MULT1029 (clk,temp_b4_1_5_r,temp_b4_1_5_i,temp_b4_1_21_r,temp_b4_1_21_i,temp_b4_17_5_r,temp_b4_17_5_i,temp_b4_17_21_r,temp_b4_17_21_i,temp_m5_1_5_r,temp_m5_1_5_i,temp_m5_1_21_r,temp_m5_1_21_i,temp_m5_17_5_r,temp_m5_17_5_i,temp_m5_17_21_r,temp_m5_17_21_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly1029 (clk,temp_m5_1_5_r,temp_m5_1_5_i,temp_m5_1_21_r,temp_m5_1_21_i,temp_m5_17_5_r,temp_m5_17_5_i,temp_m5_17_21_r,temp_m5_17_21_i,temp_b5_1_5_r,temp_b5_1_5_i,temp_b5_1_21_r,temp_b5_1_21_i,temp_b5_17_5_r,temp_b5_17_5_i,temp_b5_17_21_r,temp_b5_17_21_i);
MULT MULT1030 (clk,temp_b4_1_6_r,temp_b4_1_6_i,temp_b4_1_22_r,temp_b4_1_22_i,temp_b4_17_6_r,temp_b4_17_6_i,temp_b4_17_22_r,temp_b4_17_22_i,temp_m5_1_6_r,temp_m5_1_6_i,temp_m5_1_22_r,temp_m5_1_22_i,temp_m5_17_6_r,temp_m5_17_6_i,temp_m5_17_22_r,temp_m5_17_22_i,`W5_real,`W5_imag,`W0_real,`W0_imag,`W5_real,`W5_imag);
butterfly butterfly1030 (clk,temp_m5_1_6_r,temp_m5_1_6_i,temp_m5_1_22_r,temp_m5_1_22_i,temp_m5_17_6_r,temp_m5_17_6_i,temp_m5_17_22_r,temp_m5_17_22_i,temp_b5_1_6_r,temp_b5_1_6_i,temp_b5_1_22_r,temp_b5_1_22_i,temp_b5_17_6_r,temp_b5_17_6_i,temp_b5_17_22_r,temp_b5_17_22_i);
MULT MULT1031 (clk,temp_b4_1_7_r,temp_b4_1_7_i,temp_b4_1_23_r,temp_b4_1_23_i,temp_b4_17_7_r,temp_b4_17_7_i,temp_b4_17_23_r,temp_b4_17_23_i,temp_m5_1_7_r,temp_m5_1_7_i,temp_m5_1_23_r,temp_m5_1_23_i,temp_m5_17_7_r,temp_m5_17_7_i,temp_m5_17_23_r,temp_m5_17_23_i,`W6_real,`W6_imag,`W0_real,`W0_imag,`W6_real,`W6_imag);
butterfly butterfly1031 (clk,temp_m5_1_7_r,temp_m5_1_7_i,temp_m5_1_23_r,temp_m5_1_23_i,temp_m5_17_7_r,temp_m5_17_7_i,temp_m5_17_23_r,temp_m5_17_23_i,temp_b5_1_7_r,temp_b5_1_7_i,temp_b5_1_23_r,temp_b5_1_23_i,temp_b5_17_7_r,temp_b5_17_7_i,temp_b5_17_23_r,temp_b5_17_23_i);
MULT MULT1032 (clk,temp_b4_1_8_r,temp_b4_1_8_i,temp_b4_1_24_r,temp_b4_1_24_i,temp_b4_17_8_r,temp_b4_17_8_i,temp_b4_17_24_r,temp_b4_17_24_i,temp_m5_1_8_r,temp_m5_1_8_i,temp_m5_1_24_r,temp_m5_1_24_i,temp_m5_17_8_r,temp_m5_17_8_i,temp_m5_17_24_r,temp_m5_17_24_i,`W7_real,`W7_imag,`W0_real,`W0_imag,`W7_real,`W7_imag);
butterfly butterfly1032 (clk,temp_m5_1_8_r,temp_m5_1_8_i,temp_m5_1_24_r,temp_m5_1_24_i,temp_m5_17_8_r,temp_m5_17_8_i,temp_m5_17_24_r,temp_m5_17_24_i,temp_b5_1_8_r,temp_b5_1_8_i,temp_b5_1_24_r,temp_b5_1_24_i,temp_b5_17_8_r,temp_b5_17_8_i,temp_b5_17_24_r,temp_b5_17_24_i);
MULT MULT1033 (clk,temp_b4_1_9_r,temp_b4_1_9_i,temp_b4_1_25_r,temp_b4_1_25_i,temp_b4_17_9_r,temp_b4_17_9_i,temp_b4_17_25_r,temp_b4_17_25_i,temp_m5_1_9_r,temp_m5_1_9_i,temp_m5_1_25_r,temp_m5_1_25_i,temp_m5_17_9_r,temp_m5_17_9_i,temp_m5_17_25_r,temp_m5_17_25_i,`W8_real,`W8_imag,`W0_real,`W0_imag,`W8_real,`W8_imag);
butterfly butterfly1033 (clk,temp_m5_1_9_r,temp_m5_1_9_i,temp_m5_1_25_r,temp_m5_1_25_i,temp_m5_17_9_r,temp_m5_17_9_i,temp_m5_17_25_r,temp_m5_17_25_i,temp_b5_1_9_r,temp_b5_1_9_i,temp_b5_1_25_r,temp_b5_1_25_i,temp_b5_17_9_r,temp_b5_17_9_i,temp_b5_17_25_r,temp_b5_17_25_i);
MULT MULT1034 (clk,temp_b4_1_10_r,temp_b4_1_10_i,temp_b4_1_26_r,temp_b4_1_26_i,temp_b4_17_10_r,temp_b4_17_10_i,temp_b4_17_26_r,temp_b4_17_26_i,temp_m5_1_10_r,temp_m5_1_10_i,temp_m5_1_26_r,temp_m5_1_26_i,temp_m5_17_10_r,temp_m5_17_10_i,temp_m5_17_26_r,temp_m5_17_26_i,`W9_real,`W9_imag,`W0_real,`W0_imag,`W9_real,`W9_imag);
butterfly butterfly1034 (clk,temp_m5_1_10_r,temp_m5_1_10_i,temp_m5_1_26_r,temp_m5_1_26_i,temp_m5_17_10_r,temp_m5_17_10_i,temp_m5_17_26_r,temp_m5_17_26_i,temp_b5_1_10_r,temp_b5_1_10_i,temp_b5_1_26_r,temp_b5_1_26_i,temp_b5_17_10_r,temp_b5_17_10_i,temp_b5_17_26_r,temp_b5_17_26_i);
MULT MULT1035 (clk,temp_b4_1_11_r,temp_b4_1_11_i,temp_b4_1_27_r,temp_b4_1_27_i,temp_b4_17_11_r,temp_b4_17_11_i,temp_b4_17_27_r,temp_b4_17_27_i,temp_m5_1_11_r,temp_m5_1_11_i,temp_m5_1_27_r,temp_m5_1_27_i,temp_m5_17_11_r,temp_m5_17_11_i,temp_m5_17_27_r,temp_m5_17_27_i,`W10_real,`W10_imag,`W0_real,`W0_imag,`W10_real,`W10_imag);
butterfly butterfly1035 (clk,temp_m5_1_11_r,temp_m5_1_11_i,temp_m5_1_27_r,temp_m5_1_27_i,temp_m5_17_11_r,temp_m5_17_11_i,temp_m5_17_27_r,temp_m5_17_27_i,temp_b5_1_11_r,temp_b5_1_11_i,temp_b5_1_27_r,temp_b5_1_27_i,temp_b5_17_11_r,temp_b5_17_11_i,temp_b5_17_27_r,temp_b5_17_27_i);
MULT MULT1036 (clk,temp_b4_1_12_r,temp_b4_1_12_i,temp_b4_1_28_r,temp_b4_1_28_i,temp_b4_17_12_r,temp_b4_17_12_i,temp_b4_17_28_r,temp_b4_17_28_i,temp_m5_1_12_r,temp_m5_1_12_i,temp_m5_1_28_r,temp_m5_1_28_i,temp_m5_17_12_r,temp_m5_17_12_i,temp_m5_17_28_r,temp_m5_17_28_i,`W11_real,`W11_imag,`W0_real,`W0_imag,`W11_real,`W11_imag);
butterfly butterfly1036 (clk,temp_m5_1_12_r,temp_m5_1_12_i,temp_m5_1_28_r,temp_m5_1_28_i,temp_m5_17_12_r,temp_m5_17_12_i,temp_m5_17_28_r,temp_m5_17_28_i,temp_b5_1_12_r,temp_b5_1_12_i,temp_b5_1_28_r,temp_b5_1_28_i,temp_b5_17_12_r,temp_b5_17_12_i,temp_b5_17_28_r,temp_b5_17_28_i);
MULT MULT1037 (clk,temp_b4_1_13_r,temp_b4_1_13_i,temp_b4_1_29_r,temp_b4_1_29_i,temp_b4_17_13_r,temp_b4_17_13_i,temp_b4_17_29_r,temp_b4_17_29_i,temp_m5_1_13_r,temp_m5_1_13_i,temp_m5_1_29_r,temp_m5_1_29_i,temp_m5_17_13_r,temp_m5_17_13_i,temp_m5_17_29_r,temp_m5_17_29_i,`W12_real,`W12_imag,`W0_real,`W0_imag,`W12_real,`W12_imag);
butterfly butterfly1037 (clk,temp_m5_1_13_r,temp_m5_1_13_i,temp_m5_1_29_r,temp_m5_1_29_i,temp_m5_17_13_r,temp_m5_17_13_i,temp_m5_17_29_r,temp_m5_17_29_i,temp_b5_1_13_r,temp_b5_1_13_i,temp_b5_1_29_r,temp_b5_1_29_i,temp_b5_17_13_r,temp_b5_17_13_i,temp_b5_17_29_r,temp_b5_17_29_i);
MULT MULT1038 (clk,temp_b4_1_14_r,temp_b4_1_14_i,temp_b4_1_30_r,temp_b4_1_30_i,temp_b4_17_14_r,temp_b4_17_14_i,temp_b4_17_30_r,temp_b4_17_30_i,temp_m5_1_14_r,temp_m5_1_14_i,temp_m5_1_30_r,temp_m5_1_30_i,temp_m5_17_14_r,temp_m5_17_14_i,temp_m5_17_30_r,temp_m5_17_30_i,`W13_real,`W13_imag,`W0_real,`W0_imag,`W13_real,`W13_imag);
butterfly butterfly1038 (clk,temp_m5_1_14_r,temp_m5_1_14_i,temp_m5_1_30_r,temp_m5_1_30_i,temp_m5_17_14_r,temp_m5_17_14_i,temp_m5_17_30_r,temp_m5_17_30_i,temp_b5_1_14_r,temp_b5_1_14_i,temp_b5_1_30_r,temp_b5_1_30_i,temp_b5_17_14_r,temp_b5_17_14_i,temp_b5_17_30_r,temp_b5_17_30_i);
MULT MULT1039 (clk,temp_b4_1_15_r,temp_b4_1_15_i,temp_b4_1_31_r,temp_b4_1_31_i,temp_b4_17_15_r,temp_b4_17_15_i,temp_b4_17_31_r,temp_b4_17_31_i,temp_m5_1_15_r,temp_m5_1_15_i,temp_m5_1_31_r,temp_m5_1_31_i,temp_m5_17_15_r,temp_m5_17_15_i,temp_m5_17_31_r,temp_m5_17_31_i,`W14_real,`W14_imag,`W0_real,`W0_imag,`W14_real,`W14_imag);
butterfly butterfly1039 (clk,temp_m5_1_15_r,temp_m5_1_15_i,temp_m5_1_31_r,temp_m5_1_31_i,temp_m5_17_15_r,temp_m5_17_15_i,temp_m5_17_31_r,temp_m5_17_31_i,temp_b5_1_15_r,temp_b5_1_15_i,temp_b5_1_31_r,temp_b5_1_31_i,temp_b5_17_15_r,temp_b5_17_15_i,temp_b5_17_31_r,temp_b5_17_31_i);
MULT MULT1040 (clk,temp_b4_1_16_r,temp_b4_1_16_i,temp_b4_1_32_r,temp_b4_1_32_i,temp_b4_17_16_r,temp_b4_17_16_i,temp_b4_17_32_r,temp_b4_17_32_i,temp_m5_1_16_r,temp_m5_1_16_i,temp_m5_1_32_r,temp_m5_1_32_i,temp_m5_17_16_r,temp_m5_17_16_i,temp_m5_17_32_r,temp_m5_17_32_i,`W15_real,`W15_imag,`W0_real,`W0_imag,`W15_real,`W15_imag);
butterfly butterfly1040 (clk,temp_m5_1_16_r,temp_m5_1_16_i,temp_m5_1_32_r,temp_m5_1_32_i,temp_m5_17_16_r,temp_m5_17_16_i,temp_m5_17_32_r,temp_m5_17_32_i,temp_b5_1_16_r,temp_b5_1_16_i,temp_b5_1_32_r,temp_b5_1_32_i,temp_b5_17_16_r,temp_b5_17_16_i,temp_b5_17_32_r,temp_b5_17_32_i);
MULT MULT1041 (clk,temp_b4_2_1_r,temp_b4_2_1_i,temp_b4_2_17_r,temp_b4_2_17_i,temp_b4_18_1_r,temp_b4_18_1_i,temp_b4_18_17_r,temp_b4_18_17_i,temp_m5_2_1_r,temp_m5_2_1_i,temp_m5_2_17_r,temp_m5_2_17_i,temp_m5_18_1_r,temp_m5_18_1_i,temp_m5_18_17_r,temp_m5_18_17_i,`W0_real,`W0_imag,`W1_real,`W1_imag,`W1_real,`W1_imag);
butterfly butterfly1041 (clk,temp_m5_2_1_r,temp_m5_2_1_i,temp_m5_2_17_r,temp_m5_2_17_i,temp_m5_18_1_r,temp_m5_18_1_i,temp_m5_18_17_r,temp_m5_18_17_i,temp_b5_2_1_r,temp_b5_2_1_i,temp_b5_2_17_r,temp_b5_2_17_i,temp_b5_18_1_r,temp_b5_18_1_i,temp_b5_18_17_r,temp_b5_18_17_i);
MULT MULT1042 (clk,temp_b4_2_2_r,temp_b4_2_2_i,temp_b4_2_18_r,temp_b4_2_18_i,temp_b4_18_2_r,temp_b4_18_2_i,temp_b4_18_18_r,temp_b4_18_18_i,temp_m5_2_2_r,temp_m5_2_2_i,temp_m5_2_18_r,temp_m5_2_18_i,temp_m5_18_2_r,temp_m5_18_2_i,temp_m5_18_18_r,temp_m5_18_18_i,`W1_real,`W1_imag,`W1_real,`W1_imag,`W2_real,`W2_imag);
butterfly butterfly1042 (clk,temp_m5_2_2_r,temp_m5_2_2_i,temp_m5_2_18_r,temp_m5_2_18_i,temp_m5_18_2_r,temp_m5_18_2_i,temp_m5_18_18_r,temp_m5_18_18_i,temp_b5_2_2_r,temp_b5_2_2_i,temp_b5_2_18_r,temp_b5_2_18_i,temp_b5_18_2_r,temp_b5_18_2_i,temp_b5_18_18_r,temp_b5_18_18_i);
MULT MULT1043 (clk,temp_b4_2_3_r,temp_b4_2_3_i,temp_b4_2_19_r,temp_b4_2_19_i,temp_b4_18_3_r,temp_b4_18_3_i,temp_b4_18_19_r,temp_b4_18_19_i,temp_m5_2_3_r,temp_m5_2_3_i,temp_m5_2_19_r,temp_m5_2_19_i,temp_m5_18_3_r,temp_m5_18_3_i,temp_m5_18_19_r,temp_m5_18_19_i,`W2_real,`W2_imag,`W1_real,`W1_imag,`W3_real,`W3_imag);
butterfly butterfly1043 (clk,temp_m5_2_3_r,temp_m5_2_3_i,temp_m5_2_19_r,temp_m5_2_19_i,temp_m5_18_3_r,temp_m5_18_3_i,temp_m5_18_19_r,temp_m5_18_19_i,temp_b5_2_3_r,temp_b5_2_3_i,temp_b5_2_19_r,temp_b5_2_19_i,temp_b5_18_3_r,temp_b5_18_3_i,temp_b5_18_19_r,temp_b5_18_19_i);
MULT MULT1044 (clk,temp_b4_2_4_r,temp_b4_2_4_i,temp_b4_2_20_r,temp_b4_2_20_i,temp_b4_18_4_r,temp_b4_18_4_i,temp_b4_18_20_r,temp_b4_18_20_i,temp_m5_2_4_r,temp_m5_2_4_i,temp_m5_2_20_r,temp_m5_2_20_i,temp_m5_18_4_r,temp_m5_18_4_i,temp_m5_18_20_r,temp_m5_18_20_i,`W3_real,`W3_imag,`W1_real,`W1_imag,`W4_real,`W4_imag);
butterfly butterfly1044 (clk,temp_m5_2_4_r,temp_m5_2_4_i,temp_m5_2_20_r,temp_m5_2_20_i,temp_m5_18_4_r,temp_m5_18_4_i,temp_m5_18_20_r,temp_m5_18_20_i,temp_b5_2_4_r,temp_b5_2_4_i,temp_b5_2_20_r,temp_b5_2_20_i,temp_b5_18_4_r,temp_b5_18_4_i,temp_b5_18_20_r,temp_b5_18_20_i);
MULT MULT1045 (clk,temp_b4_2_5_r,temp_b4_2_5_i,temp_b4_2_21_r,temp_b4_2_21_i,temp_b4_18_5_r,temp_b4_18_5_i,temp_b4_18_21_r,temp_b4_18_21_i,temp_m5_2_5_r,temp_m5_2_5_i,temp_m5_2_21_r,temp_m5_2_21_i,temp_m5_18_5_r,temp_m5_18_5_i,temp_m5_18_21_r,temp_m5_18_21_i,`W4_real,`W4_imag,`W1_real,`W1_imag,`W5_real,`W5_imag);
butterfly butterfly1045 (clk,temp_m5_2_5_r,temp_m5_2_5_i,temp_m5_2_21_r,temp_m5_2_21_i,temp_m5_18_5_r,temp_m5_18_5_i,temp_m5_18_21_r,temp_m5_18_21_i,temp_b5_2_5_r,temp_b5_2_5_i,temp_b5_2_21_r,temp_b5_2_21_i,temp_b5_18_5_r,temp_b5_18_5_i,temp_b5_18_21_r,temp_b5_18_21_i);
MULT MULT1046 (clk,temp_b4_2_6_r,temp_b4_2_6_i,temp_b4_2_22_r,temp_b4_2_22_i,temp_b4_18_6_r,temp_b4_18_6_i,temp_b4_18_22_r,temp_b4_18_22_i,temp_m5_2_6_r,temp_m5_2_6_i,temp_m5_2_22_r,temp_m5_2_22_i,temp_m5_18_6_r,temp_m5_18_6_i,temp_m5_18_22_r,temp_m5_18_22_i,`W5_real,`W5_imag,`W1_real,`W1_imag,`W6_real,`W6_imag);
butterfly butterfly1046 (clk,temp_m5_2_6_r,temp_m5_2_6_i,temp_m5_2_22_r,temp_m5_2_22_i,temp_m5_18_6_r,temp_m5_18_6_i,temp_m5_18_22_r,temp_m5_18_22_i,temp_b5_2_6_r,temp_b5_2_6_i,temp_b5_2_22_r,temp_b5_2_22_i,temp_b5_18_6_r,temp_b5_18_6_i,temp_b5_18_22_r,temp_b5_18_22_i);
MULT MULT1047 (clk,temp_b4_2_7_r,temp_b4_2_7_i,temp_b4_2_23_r,temp_b4_2_23_i,temp_b4_18_7_r,temp_b4_18_7_i,temp_b4_18_23_r,temp_b4_18_23_i,temp_m5_2_7_r,temp_m5_2_7_i,temp_m5_2_23_r,temp_m5_2_23_i,temp_m5_18_7_r,temp_m5_18_7_i,temp_m5_18_23_r,temp_m5_18_23_i,`W6_real,`W6_imag,`W1_real,`W1_imag,`W7_real,`W7_imag);
butterfly butterfly1047 (clk,temp_m5_2_7_r,temp_m5_2_7_i,temp_m5_2_23_r,temp_m5_2_23_i,temp_m5_18_7_r,temp_m5_18_7_i,temp_m5_18_23_r,temp_m5_18_23_i,temp_b5_2_7_r,temp_b5_2_7_i,temp_b5_2_23_r,temp_b5_2_23_i,temp_b5_18_7_r,temp_b5_18_7_i,temp_b5_18_23_r,temp_b5_18_23_i);
MULT MULT1048 (clk,temp_b4_2_8_r,temp_b4_2_8_i,temp_b4_2_24_r,temp_b4_2_24_i,temp_b4_18_8_r,temp_b4_18_8_i,temp_b4_18_24_r,temp_b4_18_24_i,temp_m5_2_8_r,temp_m5_2_8_i,temp_m5_2_24_r,temp_m5_2_24_i,temp_m5_18_8_r,temp_m5_18_8_i,temp_m5_18_24_r,temp_m5_18_24_i,`W7_real,`W7_imag,`W1_real,`W1_imag,`W8_real,`W8_imag);
butterfly butterfly1048 (clk,temp_m5_2_8_r,temp_m5_2_8_i,temp_m5_2_24_r,temp_m5_2_24_i,temp_m5_18_8_r,temp_m5_18_8_i,temp_m5_18_24_r,temp_m5_18_24_i,temp_b5_2_8_r,temp_b5_2_8_i,temp_b5_2_24_r,temp_b5_2_24_i,temp_b5_18_8_r,temp_b5_18_8_i,temp_b5_18_24_r,temp_b5_18_24_i);
MULT MULT1049 (clk,temp_b4_2_9_r,temp_b4_2_9_i,temp_b4_2_25_r,temp_b4_2_25_i,temp_b4_18_9_r,temp_b4_18_9_i,temp_b4_18_25_r,temp_b4_18_25_i,temp_m5_2_9_r,temp_m5_2_9_i,temp_m5_2_25_r,temp_m5_2_25_i,temp_m5_18_9_r,temp_m5_18_9_i,temp_m5_18_25_r,temp_m5_18_25_i,`W8_real,`W8_imag,`W1_real,`W1_imag,`W9_real,`W9_imag);
butterfly butterfly1049 (clk,temp_m5_2_9_r,temp_m5_2_9_i,temp_m5_2_25_r,temp_m5_2_25_i,temp_m5_18_9_r,temp_m5_18_9_i,temp_m5_18_25_r,temp_m5_18_25_i,temp_b5_2_9_r,temp_b5_2_9_i,temp_b5_2_25_r,temp_b5_2_25_i,temp_b5_18_9_r,temp_b5_18_9_i,temp_b5_18_25_r,temp_b5_18_25_i);
MULT MULT1050 (clk,temp_b4_2_10_r,temp_b4_2_10_i,temp_b4_2_26_r,temp_b4_2_26_i,temp_b4_18_10_r,temp_b4_18_10_i,temp_b4_18_26_r,temp_b4_18_26_i,temp_m5_2_10_r,temp_m5_2_10_i,temp_m5_2_26_r,temp_m5_2_26_i,temp_m5_18_10_r,temp_m5_18_10_i,temp_m5_18_26_r,temp_m5_18_26_i,`W9_real,`W9_imag,`W1_real,`W1_imag,`W10_real,`W10_imag);
butterfly butterfly1050 (clk,temp_m5_2_10_r,temp_m5_2_10_i,temp_m5_2_26_r,temp_m5_2_26_i,temp_m5_18_10_r,temp_m5_18_10_i,temp_m5_18_26_r,temp_m5_18_26_i,temp_b5_2_10_r,temp_b5_2_10_i,temp_b5_2_26_r,temp_b5_2_26_i,temp_b5_18_10_r,temp_b5_18_10_i,temp_b5_18_26_r,temp_b5_18_26_i);
MULT MULT1051 (clk,temp_b4_2_11_r,temp_b4_2_11_i,temp_b4_2_27_r,temp_b4_2_27_i,temp_b4_18_11_r,temp_b4_18_11_i,temp_b4_18_27_r,temp_b4_18_27_i,temp_m5_2_11_r,temp_m5_2_11_i,temp_m5_2_27_r,temp_m5_2_27_i,temp_m5_18_11_r,temp_m5_18_11_i,temp_m5_18_27_r,temp_m5_18_27_i,`W10_real,`W10_imag,`W1_real,`W1_imag,`W11_real,`W11_imag);
butterfly butterfly1051 (clk,temp_m5_2_11_r,temp_m5_2_11_i,temp_m5_2_27_r,temp_m5_2_27_i,temp_m5_18_11_r,temp_m5_18_11_i,temp_m5_18_27_r,temp_m5_18_27_i,temp_b5_2_11_r,temp_b5_2_11_i,temp_b5_2_27_r,temp_b5_2_27_i,temp_b5_18_11_r,temp_b5_18_11_i,temp_b5_18_27_r,temp_b5_18_27_i);
MULT MULT1052 (clk,temp_b4_2_12_r,temp_b4_2_12_i,temp_b4_2_28_r,temp_b4_2_28_i,temp_b4_18_12_r,temp_b4_18_12_i,temp_b4_18_28_r,temp_b4_18_28_i,temp_m5_2_12_r,temp_m5_2_12_i,temp_m5_2_28_r,temp_m5_2_28_i,temp_m5_18_12_r,temp_m5_18_12_i,temp_m5_18_28_r,temp_m5_18_28_i,`W11_real,`W11_imag,`W1_real,`W1_imag,`W12_real,`W12_imag);
butterfly butterfly1052 (clk,temp_m5_2_12_r,temp_m5_2_12_i,temp_m5_2_28_r,temp_m5_2_28_i,temp_m5_18_12_r,temp_m5_18_12_i,temp_m5_18_28_r,temp_m5_18_28_i,temp_b5_2_12_r,temp_b5_2_12_i,temp_b5_2_28_r,temp_b5_2_28_i,temp_b5_18_12_r,temp_b5_18_12_i,temp_b5_18_28_r,temp_b5_18_28_i);
MULT MULT1053 (clk,temp_b4_2_13_r,temp_b4_2_13_i,temp_b4_2_29_r,temp_b4_2_29_i,temp_b4_18_13_r,temp_b4_18_13_i,temp_b4_18_29_r,temp_b4_18_29_i,temp_m5_2_13_r,temp_m5_2_13_i,temp_m5_2_29_r,temp_m5_2_29_i,temp_m5_18_13_r,temp_m5_18_13_i,temp_m5_18_29_r,temp_m5_18_29_i,`W12_real,`W12_imag,`W1_real,`W1_imag,`W13_real,`W13_imag);
butterfly butterfly1053 (clk,temp_m5_2_13_r,temp_m5_2_13_i,temp_m5_2_29_r,temp_m5_2_29_i,temp_m5_18_13_r,temp_m5_18_13_i,temp_m5_18_29_r,temp_m5_18_29_i,temp_b5_2_13_r,temp_b5_2_13_i,temp_b5_2_29_r,temp_b5_2_29_i,temp_b5_18_13_r,temp_b5_18_13_i,temp_b5_18_29_r,temp_b5_18_29_i);
MULT MULT1054 (clk,temp_b4_2_14_r,temp_b4_2_14_i,temp_b4_2_30_r,temp_b4_2_30_i,temp_b4_18_14_r,temp_b4_18_14_i,temp_b4_18_30_r,temp_b4_18_30_i,temp_m5_2_14_r,temp_m5_2_14_i,temp_m5_2_30_r,temp_m5_2_30_i,temp_m5_18_14_r,temp_m5_18_14_i,temp_m5_18_30_r,temp_m5_18_30_i,`W13_real,`W13_imag,`W1_real,`W1_imag,`W14_real,`W14_imag);
butterfly butterfly1054 (clk,temp_m5_2_14_r,temp_m5_2_14_i,temp_m5_2_30_r,temp_m5_2_30_i,temp_m5_18_14_r,temp_m5_18_14_i,temp_m5_18_30_r,temp_m5_18_30_i,temp_b5_2_14_r,temp_b5_2_14_i,temp_b5_2_30_r,temp_b5_2_30_i,temp_b5_18_14_r,temp_b5_18_14_i,temp_b5_18_30_r,temp_b5_18_30_i);
MULT MULT1055 (clk,temp_b4_2_15_r,temp_b4_2_15_i,temp_b4_2_31_r,temp_b4_2_31_i,temp_b4_18_15_r,temp_b4_18_15_i,temp_b4_18_31_r,temp_b4_18_31_i,temp_m5_2_15_r,temp_m5_2_15_i,temp_m5_2_31_r,temp_m5_2_31_i,temp_m5_18_15_r,temp_m5_18_15_i,temp_m5_18_31_r,temp_m5_18_31_i,`W14_real,`W14_imag,`W1_real,`W1_imag,`W15_real,`W15_imag);
butterfly butterfly1055 (clk,temp_m5_2_15_r,temp_m5_2_15_i,temp_m5_2_31_r,temp_m5_2_31_i,temp_m5_18_15_r,temp_m5_18_15_i,temp_m5_18_31_r,temp_m5_18_31_i,temp_b5_2_15_r,temp_b5_2_15_i,temp_b5_2_31_r,temp_b5_2_31_i,temp_b5_18_15_r,temp_b5_18_15_i,temp_b5_18_31_r,temp_b5_18_31_i);
MULT MULT1056 (clk,temp_b4_2_16_r,temp_b4_2_16_i,temp_b4_2_32_r,temp_b4_2_32_i,temp_b4_18_16_r,temp_b4_18_16_i,temp_b4_18_32_r,temp_b4_18_32_i,temp_m5_2_16_r,temp_m5_2_16_i,temp_m5_2_32_r,temp_m5_2_32_i,temp_m5_18_16_r,temp_m5_18_16_i,temp_m5_18_32_r,temp_m5_18_32_i,`W15_real,`W15_imag,`W1_real,`W1_imag,`W16_real,`W16_imag);
butterfly butterfly1056 (clk,temp_m5_2_16_r,temp_m5_2_16_i,temp_m5_2_32_r,temp_m5_2_32_i,temp_m5_18_16_r,temp_m5_18_16_i,temp_m5_18_32_r,temp_m5_18_32_i,temp_b5_2_16_r,temp_b5_2_16_i,temp_b5_2_32_r,temp_b5_2_32_i,temp_b5_18_16_r,temp_b5_18_16_i,temp_b5_18_32_r,temp_b5_18_32_i);
MULT MULT1057 (clk,temp_b4_3_1_r,temp_b4_3_1_i,temp_b4_3_17_r,temp_b4_3_17_i,temp_b4_19_1_r,temp_b4_19_1_i,temp_b4_19_17_r,temp_b4_19_17_i,temp_m5_3_1_r,temp_m5_3_1_i,temp_m5_3_17_r,temp_m5_3_17_i,temp_m5_19_1_r,temp_m5_19_1_i,temp_m5_19_17_r,temp_m5_19_17_i,`W0_real,`W0_imag,`W2_real,`W2_imag,`W2_real,`W2_imag);
butterfly butterfly1057 (clk,temp_m5_3_1_r,temp_m5_3_1_i,temp_m5_3_17_r,temp_m5_3_17_i,temp_m5_19_1_r,temp_m5_19_1_i,temp_m5_19_17_r,temp_m5_19_17_i,temp_b5_3_1_r,temp_b5_3_1_i,temp_b5_3_17_r,temp_b5_3_17_i,temp_b5_19_1_r,temp_b5_19_1_i,temp_b5_19_17_r,temp_b5_19_17_i);
MULT MULT1058 (clk,temp_b4_3_2_r,temp_b4_3_2_i,temp_b4_3_18_r,temp_b4_3_18_i,temp_b4_19_2_r,temp_b4_19_2_i,temp_b4_19_18_r,temp_b4_19_18_i,temp_m5_3_2_r,temp_m5_3_2_i,temp_m5_3_18_r,temp_m5_3_18_i,temp_m5_19_2_r,temp_m5_19_2_i,temp_m5_19_18_r,temp_m5_19_18_i,`W1_real,`W1_imag,`W2_real,`W2_imag,`W3_real,`W3_imag);
butterfly butterfly1058 (clk,temp_m5_3_2_r,temp_m5_3_2_i,temp_m5_3_18_r,temp_m5_3_18_i,temp_m5_19_2_r,temp_m5_19_2_i,temp_m5_19_18_r,temp_m5_19_18_i,temp_b5_3_2_r,temp_b5_3_2_i,temp_b5_3_18_r,temp_b5_3_18_i,temp_b5_19_2_r,temp_b5_19_2_i,temp_b5_19_18_r,temp_b5_19_18_i);
MULT MULT1059 (clk,temp_b4_3_3_r,temp_b4_3_3_i,temp_b4_3_19_r,temp_b4_3_19_i,temp_b4_19_3_r,temp_b4_19_3_i,temp_b4_19_19_r,temp_b4_19_19_i,temp_m5_3_3_r,temp_m5_3_3_i,temp_m5_3_19_r,temp_m5_3_19_i,temp_m5_19_3_r,temp_m5_19_3_i,temp_m5_19_19_r,temp_m5_19_19_i,`W2_real,`W2_imag,`W2_real,`W2_imag,`W4_real,`W4_imag);
butterfly butterfly1059 (clk,temp_m5_3_3_r,temp_m5_3_3_i,temp_m5_3_19_r,temp_m5_3_19_i,temp_m5_19_3_r,temp_m5_19_3_i,temp_m5_19_19_r,temp_m5_19_19_i,temp_b5_3_3_r,temp_b5_3_3_i,temp_b5_3_19_r,temp_b5_3_19_i,temp_b5_19_3_r,temp_b5_19_3_i,temp_b5_19_19_r,temp_b5_19_19_i);
MULT MULT1060 (clk,temp_b4_3_4_r,temp_b4_3_4_i,temp_b4_3_20_r,temp_b4_3_20_i,temp_b4_19_4_r,temp_b4_19_4_i,temp_b4_19_20_r,temp_b4_19_20_i,temp_m5_3_4_r,temp_m5_3_4_i,temp_m5_3_20_r,temp_m5_3_20_i,temp_m5_19_4_r,temp_m5_19_4_i,temp_m5_19_20_r,temp_m5_19_20_i,`W3_real,`W3_imag,`W2_real,`W2_imag,`W5_real,`W5_imag);
butterfly butterfly1060 (clk,temp_m5_3_4_r,temp_m5_3_4_i,temp_m5_3_20_r,temp_m5_3_20_i,temp_m5_19_4_r,temp_m5_19_4_i,temp_m5_19_20_r,temp_m5_19_20_i,temp_b5_3_4_r,temp_b5_3_4_i,temp_b5_3_20_r,temp_b5_3_20_i,temp_b5_19_4_r,temp_b5_19_4_i,temp_b5_19_20_r,temp_b5_19_20_i);
MULT MULT1061 (clk,temp_b4_3_5_r,temp_b4_3_5_i,temp_b4_3_21_r,temp_b4_3_21_i,temp_b4_19_5_r,temp_b4_19_5_i,temp_b4_19_21_r,temp_b4_19_21_i,temp_m5_3_5_r,temp_m5_3_5_i,temp_m5_3_21_r,temp_m5_3_21_i,temp_m5_19_5_r,temp_m5_19_5_i,temp_m5_19_21_r,temp_m5_19_21_i,`W4_real,`W4_imag,`W2_real,`W2_imag,`W6_real,`W6_imag);
butterfly butterfly1061 (clk,temp_m5_3_5_r,temp_m5_3_5_i,temp_m5_3_21_r,temp_m5_3_21_i,temp_m5_19_5_r,temp_m5_19_5_i,temp_m5_19_21_r,temp_m5_19_21_i,temp_b5_3_5_r,temp_b5_3_5_i,temp_b5_3_21_r,temp_b5_3_21_i,temp_b5_19_5_r,temp_b5_19_5_i,temp_b5_19_21_r,temp_b5_19_21_i);
MULT MULT1062 (clk,temp_b4_3_6_r,temp_b4_3_6_i,temp_b4_3_22_r,temp_b4_3_22_i,temp_b4_19_6_r,temp_b4_19_6_i,temp_b4_19_22_r,temp_b4_19_22_i,temp_m5_3_6_r,temp_m5_3_6_i,temp_m5_3_22_r,temp_m5_3_22_i,temp_m5_19_6_r,temp_m5_19_6_i,temp_m5_19_22_r,temp_m5_19_22_i,`W5_real,`W5_imag,`W2_real,`W2_imag,`W7_real,`W7_imag);
butterfly butterfly1062 (clk,temp_m5_3_6_r,temp_m5_3_6_i,temp_m5_3_22_r,temp_m5_3_22_i,temp_m5_19_6_r,temp_m5_19_6_i,temp_m5_19_22_r,temp_m5_19_22_i,temp_b5_3_6_r,temp_b5_3_6_i,temp_b5_3_22_r,temp_b5_3_22_i,temp_b5_19_6_r,temp_b5_19_6_i,temp_b5_19_22_r,temp_b5_19_22_i);
MULT MULT1063 (clk,temp_b4_3_7_r,temp_b4_3_7_i,temp_b4_3_23_r,temp_b4_3_23_i,temp_b4_19_7_r,temp_b4_19_7_i,temp_b4_19_23_r,temp_b4_19_23_i,temp_m5_3_7_r,temp_m5_3_7_i,temp_m5_3_23_r,temp_m5_3_23_i,temp_m5_19_7_r,temp_m5_19_7_i,temp_m5_19_23_r,temp_m5_19_23_i,`W6_real,`W6_imag,`W2_real,`W2_imag,`W8_real,`W8_imag);
butterfly butterfly1063 (clk,temp_m5_3_7_r,temp_m5_3_7_i,temp_m5_3_23_r,temp_m5_3_23_i,temp_m5_19_7_r,temp_m5_19_7_i,temp_m5_19_23_r,temp_m5_19_23_i,temp_b5_3_7_r,temp_b5_3_7_i,temp_b5_3_23_r,temp_b5_3_23_i,temp_b5_19_7_r,temp_b5_19_7_i,temp_b5_19_23_r,temp_b5_19_23_i);
MULT MULT1064 (clk,temp_b4_3_8_r,temp_b4_3_8_i,temp_b4_3_24_r,temp_b4_3_24_i,temp_b4_19_8_r,temp_b4_19_8_i,temp_b4_19_24_r,temp_b4_19_24_i,temp_m5_3_8_r,temp_m5_3_8_i,temp_m5_3_24_r,temp_m5_3_24_i,temp_m5_19_8_r,temp_m5_19_8_i,temp_m5_19_24_r,temp_m5_19_24_i,`W7_real,`W7_imag,`W2_real,`W2_imag,`W9_real,`W9_imag);
butterfly butterfly1064 (clk,temp_m5_3_8_r,temp_m5_3_8_i,temp_m5_3_24_r,temp_m5_3_24_i,temp_m5_19_8_r,temp_m5_19_8_i,temp_m5_19_24_r,temp_m5_19_24_i,temp_b5_3_8_r,temp_b5_3_8_i,temp_b5_3_24_r,temp_b5_3_24_i,temp_b5_19_8_r,temp_b5_19_8_i,temp_b5_19_24_r,temp_b5_19_24_i);
MULT MULT1065 (clk,temp_b4_3_9_r,temp_b4_3_9_i,temp_b4_3_25_r,temp_b4_3_25_i,temp_b4_19_9_r,temp_b4_19_9_i,temp_b4_19_25_r,temp_b4_19_25_i,temp_m5_3_9_r,temp_m5_3_9_i,temp_m5_3_25_r,temp_m5_3_25_i,temp_m5_19_9_r,temp_m5_19_9_i,temp_m5_19_25_r,temp_m5_19_25_i,`W8_real,`W8_imag,`W2_real,`W2_imag,`W10_real,`W10_imag);
butterfly butterfly1065 (clk,temp_m5_3_9_r,temp_m5_3_9_i,temp_m5_3_25_r,temp_m5_3_25_i,temp_m5_19_9_r,temp_m5_19_9_i,temp_m5_19_25_r,temp_m5_19_25_i,temp_b5_3_9_r,temp_b5_3_9_i,temp_b5_3_25_r,temp_b5_3_25_i,temp_b5_19_9_r,temp_b5_19_9_i,temp_b5_19_25_r,temp_b5_19_25_i);
MULT MULT1066 (clk,temp_b4_3_10_r,temp_b4_3_10_i,temp_b4_3_26_r,temp_b4_3_26_i,temp_b4_19_10_r,temp_b4_19_10_i,temp_b4_19_26_r,temp_b4_19_26_i,temp_m5_3_10_r,temp_m5_3_10_i,temp_m5_3_26_r,temp_m5_3_26_i,temp_m5_19_10_r,temp_m5_19_10_i,temp_m5_19_26_r,temp_m5_19_26_i,`W9_real,`W9_imag,`W2_real,`W2_imag,`W11_real,`W11_imag);
butterfly butterfly1066 (clk,temp_m5_3_10_r,temp_m5_3_10_i,temp_m5_3_26_r,temp_m5_3_26_i,temp_m5_19_10_r,temp_m5_19_10_i,temp_m5_19_26_r,temp_m5_19_26_i,temp_b5_3_10_r,temp_b5_3_10_i,temp_b5_3_26_r,temp_b5_3_26_i,temp_b5_19_10_r,temp_b5_19_10_i,temp_b5_19_26_r,temp_b5_19_26_i);
MULT MULT1067 (clk,temp_b4_3_11_r,temp_b4_3_11_i,temp_b4_3_27_r,temp_b4_3_27_i,temp_b4_19_11_r,temp_b4_19_11_i,temp_b4_19_27_r,temp_b4_19_27_i,temp_m5_3_11_r,temp_m5_3_11_i,temp_m5_3_27_r,temp_m5_3_27_i,temp_m5_19_11_r,temp_m5_19_11_i,temp_m5_19_27_r,temp_m5_19_27_i,`W10_real,`W10_imag,`W2_real,`W2_imag,`W12_real,`W12_imag);
butterfly butterfly1067 (clk,temp_m5_3_11_r,temp_m5_3_11_i,temp_m5_3_27_r,temp_m5_3_27_i,temp_m5_19_11_r,temp_m5_19_11_i,temp_m5_19_27_r,temp_m5_19_27_i,temp_b5_3_11_r,temp_b5_3_11_i,temp_b5_3_27_r,temp_b5_3_27_i,temp_b5_19_11_r,temp_b5_19_11_i,temp_b5_19_27_r,temp_b5_19_27_i);
MULT MULT1068 (clk,temp_b4_3_12_r,temp_b4_3_12_i,temp_b4_3_28_r,temp_b4_3_28_i,temp_b4_19_12_r,temp_b4_19_12_i,temp_b4_19_28_r,temp_b4_19_28_i,temp_m5_3_12_r,temp_m5_3_12_i,temp_m5_3_28_r,temp_m5_3_28_i,temp_m5_19_12_r,temp_m5_19_12_i,temp_m5_19_28_r,temp_m5_19_28_i,`W11_real,`W11_imag,`W2_real,`W2_imag,`W13_real,`W13_imag);
butterfly butterfly1068 (clk,temp_m5_3_12_r,temp_m5_3_12_i,temp_m5_3_28_r,temp_m5_3_28_i,temp_m5_19_12_r,temp_m5_19_12_i,temp_m5_19_28_r,temp_m5_19_28_i,temp_b5_3_12_r,temp_b5_3_12_i,temp_b5_3_28_r,temp_b5_3_28_i,temp_b5_19_12_r,temp_b5_19_12_i,temp_b5_19_28_r,temp_b5_19_28_i);
MULT MULT1069 (clk,temp_b4_3_13_r,temp_b4_3_13_i,temp_b4_3_29_r,temp_b4_3_29_i,temp_b4_19_13_r,temp_b4_19_13_i,temp_b4_19_29_r,temp_b4_19_29_i,temp_m5_3_13_r,temp_m5_3_13_i,temp_m5_3_29_r,temp_m5_3_29_i,temp_m5_19_13_r,temp_m5_19_13_i,temp_m5_19_29_r,temp_m5_19_29_i,`W12_real,`W12_imag,`W2_real,`W2_imag,`W14_real,`W14_imag);
butterfly butterfly1069 (clk,temp_m5_3_13_r,temp_m5_3_13_i,temp_m5_3_29_r,temp_m5_3_29_i,temp_m5_19_13_r,temp_m5_19_13_i,temp_m5_19_29_r,temp_m5_19_29_i,temp_b5_3_13_r,temp_b5_3_13_i,temp_b5_3_29_r,temp_b5_3_29_i,temp_b5_19_13_r,temp_b5_19_13_i,temp_b5_19_29_r,temp_b5_19_29_i);
MULT MULT1070 (clk,temp_b4_3_14_r,temp_b4_3_14_i,temp_b4_3_30_r,temp_b4_3_30_i,temp_b4_19_14_r,temp_b4_19_14_i,temp_b4_19_30_r,temp_b4_19_30_i,temp_m5_3_14_r,temp_m5_3_14_i,temp_m5_3_30_r,temp_m5_3_30_i,temp_m5_19_14_r,temp_m5_19_14_i,temp_m5_19_30_r,temp_m5_19_30_i,`W13_real,`W13_imag,`W2_real,`W2_imag,`W15_real,`W15_imag);
butterfly butterfly1070 (clk,temp_m5_3_14_r,temp_m5_3_14_i,temp_m5_3_30_r,temp_m5_3_30_i,temp_m5_19_14_r,temp_m5_19_14_i,temp_m5_19_30_r,temp_m5_19_30_i,temp_b5_3_14_r,temp_b5_3_14_i,temp_b5_3_30_r,temp_b5_3_30_i,temp_b5_19_14_r,temp_b5_19_14_i,temp_b5_19_30_r,temp_b5_19_30_i);
MULT MULT1071 (clk,temp_b4_3_15_r,temp_b4_3_15_i,temp_b4_3_31_r,temp_b4_3_31_i,temp_b4_19_15_r,temp_b4_19_15_i,temp_b4_19_31_r,temp_b4_19_31_i,temp_m5_3_15_r,temp_m5_3_15_i,temp_m5_3_31_r,temp_m5_3_31_i,temp_m5_19_15_r,temp_m5_19_15_i,temp_m5_19_31_r,temp_m5_19_31_i,`W14_real,`W14_imag,`W2_real,`W2_imag,`W16_real,`W16_imag);
butterfly butterfly1071 (clk,temp_m5_3_15_r,temp_m5_3_15_i,temp_m5_3_31_r,temp_m5_3_31_i,temp_m5_19_15_r,temp_m5_19_15_i,temp_m5_19_31_r,temp_m5_19_31_i,temp_b5_3_15_r,temp_b5_3_15_i,temp_b5_3_31_r,temp_b5_3_31_i,temp_b5_19_15_r,temp_b5_19_15_i,temp_b5_19_31_r,temp_b5_19_31_i);
MULT MULT1072 (clk,temp_b4_3_16_r,temp_b4_3_16_i,temp_b4_3_32_r,temp_b4_3_32_i,temp_b4_19_16_r,temp_b4_19_16_i,temp_b4_19_32_r,temp_b4_19_32_i,temp_m5_3_16_r,temp_m5_3_16_i,temp_m5_3_32_r,temp_m5_3_32_i,temp_m5_19_16_r,temp_m5_19_16_i,temp_m5_19_32_r,temp_m5_19_32_i,`W15_real,`W15_imag,`W2_real,`W2_imag,`W17_real,`W17_imag);
butterfly butterfly1072 (clk,temp_m5_3_16_r,temp_m5_3_16_i,temp_m5_3_32_r,temp_m5_3_32_i,temp_m5_19_16_r,temp_m5_19_16_i,temp_m5_19_32_r,temp_m5_19_32_i,temp_b5_3_16_r,temp_b5_3_16_i,temp_b5_3_32_r,temp_b5_3_32_i,temp_b5_19_16_r,temp_b5_19_16_i,temp_b5_19_32_r,temp_b5_19_32_i);
MULT MULT1073 (clk,temp_b4_4_1_r,temp_b4_4_1_i,temp_b4_4_17_r,temp_b4_4_17_i,temp_b4_20_1_r,temp_b4_20_1_i,temp_b4_20_17_r,temp_b4_20_17_i,temp_m5_4_1_r,temp_m5_4_1_i,temp_m5_4_17_r,temp_m5_4_17_i,temp_m5_20_1_r,temp_m5_20_1_i,temp_m5_20_17_r,temp_m5_20_17_i,`W0_real,`W0_imag,`W3_real,`W3_imag,`W3_real,`W3_imag);
butterfly butterfly1073 (clk,temp_m5_4_1_r,temp_m5_4_1_i,temp_m5_4_17_r,temp_m5_4_17_i,temp_m5_20_1_r,temp_m5_20_1_i,temp_m5_20_17_r,temp_m5_20_17_i,temp_b5_4_1_r,temp_b5_4_1_i,temp_b5_4_17_r,temp_b5_4_17_i,temp_b5_20_1_r,temp_b5_20_1_i,temp_b5_20_17_r,temp_b5_20_17_i);
MULT MULT1074 (clk,temp_b4_4_2_r,temp_b4_4_2_i,temp_b4_4_18_r,temp_b4_4_18_i,temp_b4_20_2_r,temp_b4_20_2_i,temp_b4_20_18_r,temp_b4_20_18_i,temp_m5_4_2_r,temp_m5_4_2_i,temp_m5_4_18_r,temp_m5_4_18_i,temp_m5_20_2_r,temp_m5_20_2_i,temp_m5_20_18_r,temp_m5_20_18_i,`W1_real,`W1_imag,`W3_real,`W3_imag,`W4_real,`W4_imag);
butterfly butterfly1074 (clk,temp_m5_4_2_r,temp_m5_4_2_i,temp_m5_4_18_r,temp_m5_4_18_i,temp_m5_20_2_r,temp_m5_20_2_i,temp_m5_20_18_r,temp_m5_20_18_i,temp_b5_4_2_r,temp_b5_4_2_i,temp_b5_4_18_r,temp_b5_4_18_i,temp_b5_20_2_r,temp_b5_20_2_i,temp_b5_20_18_r,temp_b5_20_18_i);
MULT MULT1075 (clk,temp_b4_4_3_r,temp_b4_4_3_i,temp_b4_4_19_r,temp_b4_4_19_i,temp_b4_20_3_r,temp_b4_20_3_i,temp_b4_20_19_r,temp_b4_20_19_i,temp_m5_4_3_r,temp_m5_4_3_i,temp_m5_4_19_r,temp_m5_4_19_i,temp_m5_20_3_r,temp_m5_20_3_i,temp_m5_20_19_r,temp_m5_20_19_i,`W2_real,`W2_imag,`W3_real,`W3_imag,`W5_real,`W5_imag);
butterfly butterfly1075 (clk,temp_m5_4_3_r,temp_m5_4_3_i,temp_m5_4_19_r,temp_m5_4_19_i,temp_m5_20_3_r,temp_m5_20_3_i,temp_m5_20_19_r,temp_m5_20_19_i,temp_b5_4_3_r,temp_b5_4_3_i,temp_b5_4_19_r,temp_b5_4_19_i,temp_b5_20_3_r,temp_b5_20_3_i,temp_b5_20_19_r,temp_b5_20_19_i);
MULT MULT1076 (clk,temp_b4_4_4_r,temp_b4_4_4_i,temp_b4_4_20_r,temp_b4_4_20_i,temp_b4_20_4_r,temp_b4_20_4_i,temp_b4_20_20_r,temp_b4_20_20_i,temp_m5_4_4_r,temp_m5_4_4_i,temp_m5_4_20_r,temp_m5_4_20_i,temp_m5_20_4_r,temp_m5_20_4_i,temp_m5_20_20_r,temp_m5_20_20_i,`W3_real,`W3_imag,`W3_real,`W3_imag,`W6_real,`W6_imag);
butterfly butterfly1076 (clk,temp_m5_4_4_r,temp_m5_4_4_i,temp_m5_4_20_r,temp_m5_4_20_i,temp_m5_20_4_r,temp_m5_20_4_i,temp_m5_20_20_r,temp_m5_20_20_i,temp_b5_4_4_r,temp_b5_4_4_i,temp_b5_4_20_r,temp_b5_4_20_i,temp_b5_20_4_r,temp_b5_20_4_i,temp_b5_20_20_r,temp_b5_20_20_i);
MULT MULT1077 (clk,temp_b4_4_5_r,temp_b4_4_5_i,temp_b4_4_21_r,temp_b4_4_21_i,temp_b4_20_5_r,temp_b4_20_5_i,temp_b4_20_21_r,temp_b4_20_21_i,temp_m5_4_5_r,temp_m5_4_5_i,temp_m5_4_21_r,temp_m5_4_21_i,temp_m5_20_5_r,temp_m5_20_5_i,temp_m5_20_21_r,temp_m5_20_21_i,`W4_real,`W4_imag,`W3_real,`W3_imag,`W7_real,`W7_imag);
butterfly butterfly1077 (clk,temp_m5_4_5_r,temp_m5_4_5_i,temp_m5_4_21_r,temp_m5_4_21_i,temp_m5_20_5_r,temp_m5_20_5_i,temp_m5_20_21_r,temp_m5_20_21_i,temp_b5_4_5_r,temp_b5_4_5_i,temp_b5_4_21_r,temp_b5_4_21_i,temp_b5_20_5_r,temp_b5_20_5_i,temp_b5_20_21_r,temp_b5_20_21_i);
MULT MULT1078 (clk,temp_b4_4_6_r,temp_b4_4_6_i,temp_b4_4_22_r,temp_b4_4_22_i,temp_b4_20_6_r,temp_b4_20_6_i,temp_b4_20_22_r,temp_b4_20_22_i,temp_m5_4_6_r,temp_m5_4_6_i,temp_m5_4_22_r,temp_m5_4_22_i,temp_m5_20_6_r,temp_m5_20_6_i,temp_m5_20_22_r,temp_m5_20_22_i,`W5_real,`W5_imag,`W3_real,`W3_imag,`W8_real,`W8_imag);
butterfly butterfly1078 (clk,temp_m5_4_6_r,temp_m5_4_6_i,temp_m5_4_22_r,temp_m5_4_22_i,temp_m5_20_6_r,temp_m5_20_6_i,temp_m5_20_22_r,temp_m5_20_22_i,temp_b5_4_6_r,temp_b5_4_6_i,temp_b5_4_22_r,temp_b5_4_22_i,temp_b5_20_6_r,temp_b5_20_6_i,temp_b5_20_22_r,temp_b5_20_22_i);
MULT MULT1079 (clk,temp_b4_4_7_r,temp_b4_4_7_i,temp_b4_4_23_r,temp_b4_4_23_i,temp_b4_20_7_r,temp_b4_20_7_i,temp_b4_20_23_r,temp_b4_20_23_i,temp_m5_4_7_r,temp_m5_4_7_i,temp_m5_4_23_r,temp_m5_4_23_i,temp_m5_20_7_r,temp_m5_20_7_i,temp_m5_20_23_r,temp_m5_20_23_i,`W6_real,`W6_imag,`W3_real,`W3_imag,`W9_real,`W9_imag);
butterfly butterfly1079 (clk,temp_m5_4_7_r,temp_m5_4_7_i,temp_m5_4_23_r,temp_m5_4_23_i,temp_m5_20_7_r,temp_m5_20_7_i,temp_m5_20_23_r,temp_m5_20_23_i,temp_b5_4_7_r,temp_b5_4_7_i,temp_b5_4_23_r,temp_b5_4_23_i,temp_b5_20_7_r,temp_b5_20_7_i,temp_b5_20_23_r,temp_b5_20_23_i);
MULT MULT1080 (clk,temp_b4_4_8_r,temp_b4_4_8_i,temp_b4_4_24_r,temp_b4_4_24_i,temp_b4_20_8_r,temp_b4_20_8_i,temp_b4_20_24_r,temp_b4_20_24_i,temp_m5_4_8_r,temp_m5_4_8_i,temp_m5_4_24_r,temp_m5_4_24_i,temp_m5_20_8_r,temp_m5_20_8_i,temp_m5_20_24_r,temp_m5_20_24_i,`W7_real,`W7_imag,`W3_real,`W3_imag,`W10_real,`W10_imag);
butterfly butterfly1080 (clk,temp_m5_4_8_r,temp_m5_4_8_i,temp_m5_4_24_r,temp_m5_4_24_i,temp_m5_20_8_r,temp_m5_20_8_i,temp_m5_20_24_r,temp_m5_20_24_i,temp_b5_4_8_r,temp_b5_4_8_i,temp_b5_4_24_r,temp_b5_4_24_i,temp_b5_20_8_r,temp_b5_20_8_i,temp_b5_20_24_r,temp_b5_20_24_i);
MULT MULT1081 (clk,temp_b4_4_9_r,temp_b4_4_9_i,temp_b4_4_25_r,temp_b4_4_25_i,temp_b4_20_9_r,temp_b4_20_9_i,temp_b4_20_25_r,temp_b4_20_25_i,temp_m5_4_9_r,temp_m5_4_9_i,temp_m5_4_25_r,temp_m5_4_25_i,temp_m5_20_9_r,temp_m5_20_9_i,temp_m5_20_25_r,temp_m5_20_25_i,`W8_real,`W8_imag,`W3_real,`W3_imag,`W11_real,`W11_imag);
butterfly butterfly1081 (clk,temp_m5_4_9_r,temp_m5_4_9_i,temp_m5_4_25_r,temp_m5_4_25_i,temp_m5_20_9_r,temp_m5_20_9_i,temp_m5_20_25_r,temp_m5_20_25_i,temp_b5_4_9_r,temp_b5_4_9_i,temp_b5_4_25_r,temp_b5_4_25_i,temp_b5_20_9_r,temp_b5_20_9_i,temp_b5_20_25_r,temp_b5_20_25_i);
MULT MULT1082 (clk,temp_b4_4_10_r,temp_b4_4_10_i,temp_b4_4_26_r,temp_b4_4_26_i,temp_b4_20_10_r,temp_b4_20_10_i,temp_b4_20_26_r,temp_b4_20_26_i,temp_m5_4_10_r,temp_m5_4_10_i,temp_m5_4_26_r,temp_m5_4_26_i,temp_m5_20_10_r,temp_m5_20_10_i,temp_m5_20_26_r,temp_m5_20_26_i,`W9_real,`W9_imag,`W3_real,`W3_imag,`W12_real,`W12_imag);
butterfly butterfly1082 (clk,temp_m5_4_10_r,temp_m5_4_10_i,temp_m5_4_26_r,temp_m5_4_26_i,temp_m5_20_10_r,temp_m5_20_10_i,temp_m5_20_26_r,temp_m5_20_26_i,temp_b5_4_10_r,temp_b5_4_10_i,temp_b5_4_26_r,temp_b5_4_26_i,temp_b5_20_10_r,temp_b5_20_10_i,temp_b5_20_26_r,temp_b5_20_26_i);
MULT MULT1083 (clk,temp_b4_4_11_r,temp_b4_4_11_i,temp_b4_4_27_r,temp_b4_4_27_i,temp_b4_20_11_r,temp_b4_20_11_i,temp_b4_20_27_r,temp_b4_20_27_i,temp_m5_4_11_r,temp_m5_4_11_i,temp_m5_4_27_r,temp_m5_4_27_i,temp_m5_20_11_r,temp_m5_20_11_i,temp_m5_20_27_r,temp_m5_20_27_i,`W10_real,`W10_imag,`W3_real,`W3_imag,`W13_real,`W13_imag);
butterfly butterfly1083 (clk,temp_m5_4_11_r,temp_m5_4_11_i,temp_m5_4_27_r,temp_m5_4_27_i,temp_m5_20_11_r,temp_m5_20_11_i,temp_m5_20_27_r,temp_m5_20_27_i,temp_b5_4_11_r,temp_b5_4_11_i,temp_b5_4_27_r,temp_b5_4_27_i,temp_b5_20_11_r,temp_b5_20_11_i,temp_b5_20_27_r,temp_b5_20_27_i);
MULT MULT1084 (clk,temp_b4_4_12_r,temp_b4_4_12_i,temp_b4_4_28_r,temp_b4_4_28_i,temp_b4_20_12_r,temp_b4_20_12_i,temp_b4_20_28_r,temp_b4_20_28_i,temp_m5_4_12_r,temp_m5_4_12_i,temp_m5_4_28_r,temp_m5_4_28_i,temp_m5_20_12_r,temp_m5_20_12_i,temp_m5_20_28_r,temp_m5_20_28_i,`W11_real,`W11_imag,`W3_real,`W3_imag,`W14_real,`W14_imag);
butterfly butterfly1084 (clk,temp_m5_4_12_r,temp_m5_4_12_i,temp_m5_4_28_r,temp_m5_4_28_i,temp_m5_20_12_r,temp_m5_20_12_i,temp_m5_20_28_r,temp_m5_20_28_i,temp_b5_4_12_r,temp_b5_4_12_i,temp_b5_4_28_r,temp_b5_4_28_i,temp_b5_20_12_r,temp_b5_20_12_i,temp_b5_20_28_r,temp_b5_20_28_i);
MULT MULT1085 (clk,temp_b4_4_13_r,temp_b4_4_13_i,temp_b4_4_29_r,temp_b4_4_29_i,temp_b4_20_13_r,temp_b4_20_13_i,temp_b4_20_29_r,temp_b4_20_29_i,temp_m5_4_13_r,temp_m5_4_13_i,temp_m5_4_29_r,temp_m5_4_29_i,temp_m5_20_13_r,temp_m5_20_13_i,temp_m5_20_29_r,temp_m5_20_29_i,`W12_real,`W12_imag,`W3_real,`W3_imag,`W15_real,`W15_imag);
butterfly butterfly1085 (clk,temp_m5_4_13_r,temp_m5_4_13_i,temp_m5_4_29_r,temp_m5_4_29_i,temp_m5_20_13_r,temp_m5_20_13_i,temp_m5_20_29_r,temp_m5_20_29_i,temp_b5_4_13_r,temp_b5_4_13_i,temp_b5_4_29_r,temp_b5_4_29_i,temp_b5_20_13_r,temp_b5_20_13_i,temp_b5_20_29_r,temp_b5_20_29_i);
MULT MULT1086 (clk,temp_b4_4_14_r,temp_b4_4_14_i,temp_b4_4_30_r,temp_b4_4_30_i,temp_b4_20_14_r,temp_b4_20_14_i,temp_b4_20_30_r,temp_b4_20_30_i,temp_m5_4_14_r,temp_m5_4_14_i,temp_m5_4_30_r,temp_m5_4_30_i,temp_m5_20_14_r,temp_m5_20_14_i,temp_m5_20_30_r,temp_m5_20_30_i,`W13_real,`W13_imag,`W3_real,`W3_imag,`W16_real,`W16_imag);
butterfly butterfly1086 (clk,temp_m5_4_14_r,temp_m5_4_14_i,temp_m5_4_30_r,temp_m5_4_30_i,temp_m5_20_14_r,temp_m5_20_14_i,temp_m5_20_30_r,temp_m5_20_30_i,temp_b5_4_14_r,temp_b5_4_14_i,temp_b5_4_30_r,temp_b5_4_30_i,temp_b5_20_14_r,temp_b5_20_14_i,temp_b5_20_30_r,temp_b5_20_30_i);
MULT MULT1087 (clk,temp_b4_4_15_r,temp_b4_4_15_i,temp_b4_4_31_r,temp_b4_4_31_i,temp_b4_20_15_r,temp_b4_20_15_i,temp_b4_20_31_r,temp_b4_20_31_i,temp_m5_4_15_r,temp_m5_4_15_i,temp_m5_4_31_r,temp_m5_4_31_i,temp_m5_20_15_r,temp_m5_20_15_i,temp_m5_20_31_r,temp_m5_20_31_i,`W14_real,`W14_imag,`W3_real,`W3_imag,`W17_real,`W17_imag);
butterfly butterfly1087 (clk,temp_m5_4_15_r,temp_m5_4_15_i,temp_m5_4_31_r,temp_m5_4_31_i,temp_m5_20_15_r,temp_m5_20_15_i,temp_m5_20_31_r,temp_m5_20_31_i,temp_b5_4_15_r,temp_b5_4_15_i,temp_b5_4_31_r,temp_b5_4_31_i,temp_b5_20_15_r,temp_b5_20_15_i,temp_b5_20_31_r,temp_b5_20_31_i);
MULT MULT1088 (clk,temp_b4_4_16_r,temp_b4_4_16_i,temp_b4_4_32_r,temp_b4_4_32_i,temp_b4_20_16_r,temp_b4_20_16_i,temp_b4_20_32_r,temp_b4_20_32_i,temp_m5_4_16_r,temp_m5_4_16_i,temp_m5_4_32_r,temp_m5_4_32_i,temp_m5_20_16_r,temp_m5_20_16_i,temp_m5_20_32_r,temp_m5_20_32_i,`W15_real,`W15_imag,`W3_real,`W3_imag,`W18_real,`W18_imag);
butterfly butterfly1088 (clk,temp_m5_4_16_r,temp_m5_4_16_i,temp_m5_4_32_r,temp_m5_4_32_i,temp_m5_20_16_r,temp_m5_20_16_i,temp_m5_20_32_r,temp_m5_20_32_i,temp_b5_4_16_r,temp_b5_4_16_i,temp_b5_4_32_r,temp_b5_4_32_i,temp_b5_20_16_r,temp_b5_20_16_i,temp_b5_20_32_r,temp_b5_20_32_i);
MULT MULT1089 (clk,temp_b4_5_1_r,temp_b4_5_1_i,temp_b4_5_17_r,temp_b4_5_17_i,temp_b4_21_1_r,temp_b4_21_1_i,temp_b4_21_17_r,temp_b4_21_17_i,temp_m5_5_1_r,temp_m5_5_1_i,temp_m5_5_17_r,temp_m5_5_17_i,temp_m5_21_1_r,temp_m5_21_1_i,temp_m5_21_17_r,temp_m5_21_17_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly1089 (clk,temp_m5_5_1_r,temp_m5_5_1_i,temp_m5_5_17_r,temp_m5_5_17_i,temp_m5_21_1_r,temp_m5_21_1_i,temp_m5_21_17_r,temp_m5_21_17_i,temp_b5_5_1_r,temp_b5_5_1_i,temp_b5_5_17_r,temp_b5_5_17_i,temp_b5_21_1_r,temp_b5_21_1_i,temp_b5_21_17_r,temp_b5_21_17_i);
MULT MULT1090 (clk,temp_b4_5_2_r,temp_b4_5_2_i,temp_b4_5_18_r,temp_b4_5_18_i,temp_b4_21_2_r,temp_b4_21_2_i,temp_b4_21_18_r,temp_b4_21_18_i,temp_m5_5_2_r,temp_m5_5_2_i,temp_m5_5_18_r,temp_m5_5_18_i,temp_m5_21_2_r,temp_m5_21_2_i,temp_m5_21_18_r,temp_m5_21_18_i,`W1_real,`W1_imag,`W4_real,`W4_imag,`W5_real,`W5_imag);
butterfly butterfly1090 (clk,temp_m5_5_2_r,temp_m5_5_2_i,temp_m5_5_18_r,temp_m5_5_18_i,temp_m5_21_2_r,temp_m5_21_2_i,temp_m5_21_18_r,temp_m5_21_18_i,temp_b5_5_2_r,temp_b5_5_2_i,temp_b5_5_18_r,temp_b5_5_18_i,temp_b5_21_2_r,temp_b5_21_2_i,temp_b5_21_18_r,temp_b5_21_18_i);
MULT MULT1091 (clk,temp_b4_5_3_r,temp_b4_5_3_i,temp_b4_5_19_r,temp_b4_5_19_i,temp_b4_21_3_r,temp_b4_21_3_i,temp_b4_21_19_r,temp_b4_21_19_i,temp_m5_5_3_r,temp_m5_5_3_i,temp_m5_5_19_r,temp_m5_5_19_i,temp_m5_21_3_r,temp_m5_21_3_i,temp_m5_21_19_r,temp_m5_21_19_i,`W2_real,`W2_imag,`W4_real,`W4_imag,`W6_real,`W6_imag);
butterfly butterfly1091 (clk,temp_m5_5_3_r,temp_m5_5_3_i,temp_m5_5_19_r,temp_m5_5_19_i,temp_m5_21_3_r,temp_m5_21_3_i,temp_m5_21_19_r,temp_m5_21_19_i,temp_b5_5_3_r,temp_b5_5_3_i,temp_b5_5_19_r,temp_b5_5_19_i,temp_b5_21_3_r,temp_b5_21_3_i,temp_b5_21_19_r,temp_b5_21_19_i);
MULT MULT1092 (clk,temp_b4_5_4_r,temp_b4_5_4_i,temp_b4_5_20_r,temp_b4_5_20_i,temp_b4_21_4_r,temp_b4_21_4_i,temp_b4_21_20_r,temp_b4_21_20_i,temp_m5_5_4_r,temp_m5_5_4_i,temp_m5_5_20_r,temp_m5_5_20_i,temp_m5_21_4_r,temp_m5_21_4_i,temp_m5_21_20_r,temp_m5_21_20_i,`W3_real,`W3_imag,`W4_real,`W4_imag,`W7_real,`W7_imag);
butterfly butterfly1092 (clk,temp_m5_5_4_r,temp_m5_5_4_i,temp_m5_5_20_r,temp_m5_5_20_i,temp_m5_21_4_r,temp_m5_21_4_i,temp_m5_21_20_r,temp_m5_21_20_i,temp_b5_5_4_r,temp_b5_5_4_i,temp_b5_5_20_r,temp_b5_5_20_i,temp_b5_21_4_r,temp_b5_21_4_i,temp_b5_21_20_r,temp_b5_21_20_i);
MULT MULT1093 (clk,temp_b4_5_5_r,temp_b4_5_5_i,temp_b4_5_21_r,temp_b4_5_21_i,temp_b4_21_5_r,temp_b4_21_5_i,temp_b4_21_21_r,temp_b4_21_21_i,temp_m5_5_5_r,temp_m5_5_5_i,temp_m5_5_21_r,temp_m5_5_21_i,temp_m5_21_5_r,temp_m5_21_5_i,temp_m5_21_21_r,temp_m5_21_21_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly1093 (clk,temp_m5_5_5_r,temp_m5_5_5_i,temp_m5_5_21_r,temp_m5_5_21_i,temp_m5_21_5_r,temp_m5_21_5_i,temp_m5_21_21_r,temp_m5_21_21_i,temp_b5_5_5_r,temp_b5_5_5_i,temp_b5_5_21_r,temp_b5_5_21_i,temp_b5_21_5_r,temp_b5_21_5_i,temp_b5_21_21_r,temp_b5_21_21_i);
MULT MULT1094 (clk,temp_b4_5_6_r,temp_b4_5_6_i,temp_b4_5_22_r,temp_b4_5_22_i,temp_b4_21_6_r,temp_b4_21_6_i,temp_b4_21_22_r,temp_b4_21_22_i,temp_m5_5_6_r,temp_m5_5_6_i,temp_m5_5_22_r,temp_m5_5_22_i,temp_m5_21_6_r,temp_m5_21_6_i,temp_m5_21_22_r,temp_m5_21_22_i,`W5_real,`W5_imag,`W4_real,`W4_imag,`W9_real,`W9_imag);
butterfly butterfly1094 (clk,temp_m5_5_6_r,temp_m5_5_6_i,temp_m5_5_22_r,temp_m5_5_22_i,temp_m5_21_6_r,temp_m5_21_6_i,temp_m5_21_22_r,temp_m5_21_22_i,temp_b5_5_6_r,temp_b5_5_6_i,temp_b5_5_22_r,temp_b5_5_22_i,temp_b5_21_6_r,temp_b5_21_6_i,temp_b5_21_22_r,temp_b5_21_22_i);
MULT MULT1095 (clk,temp_b4_5_7_r,temp_b4_5_7_i,temp_b4_5_23_r,temp_b4_5_23_i,temp_b4_21_7_r,temp_b4_21_7_i,temp_b4_21_23_r,temp_b4_21_23_i,temp_m5_5_7_r,temp_m5_5_7_i,temp_m5_5_23_r,temp_m5_5_23_i,temp_m5_21_7_r,temp_m5_21_7_i,temp_m5_21_23_r,temp_m5_21_23_i,`W6_real,`W6_imag,`W4_real,`W4_imag,`W10_real,`W10_imag);
butterfly butterfly1095 (clk,temp_m5_5_7_r,temp_m5_5_7_i,temp_m5_5_23_r,temp_m5_5_23_i,temp_m5_21_7_r,temp_m5_21_7_i,temp_m5_21_23_r,temp_m5_21_23_i,temp_b5_5_7_r,temp_b5_5_7_i,temp_b5_5_23_r,temp_b5_5_23_i,temp_b5_21_7_r,temp_b5_21_7_i,temp_b5_21_23_r,temp_b5_21_23_i);
MULT MULT1096 (clk,temp_b4_5_8_r,temp_b4_5_8_i,temp_b4_5_24_r,temp_b4_5_24_i,temp_b4_21_8_r,temp_b4_21_8_i,temp_b4_21_24_r,temp_b4_21_24_i,temp_m5_5_8_r,temp_m5_5_8_i,temp_m5_5_24_r,temp_m5_5_24_i,temp_m5_21_8_r,temp_m5_21_8_i,temp_m5_21_24_r,temp_m5_21_24_i,`W7_real,`W7_imag,`W4_real,`W4_imag,`W11_real,`W11_imag);
butterfly butterfly1096 (clk,temp_m5_5_8_r,temp_m5_5_8_i,temp_m5_5_24_r,temp_m5_5_24_i,temp_m5_21_8_r,temp_m5_21_8_i,temp_m5_21_24_r,temp_m5_21_24_i,temp_b5_5_8_r,temp_b5_5_8_i,temp_b5_5_24_r,temp_b5_5_24_i,temp_b5_21_8_r,temp_b5_21_8_i,temp_b5_21_24_r,temp_b5_21_24_i);
MULT MULT1097 (clk,temp_b4_5_9_r,temp_b4_5_9_i,temp_b4_5_25_r,temp_b4_5_25_i,temp_b4_21_9_r,temp_b4_21_9_i,temp_b4_21_25_r,temp_b4_21_25_i,temp_m5_5_9_r,temp_m5_5_9_i,temp_m5_5_25_r,temp_m5_5_25_i,temp_m5_21_9_r,temp_m5_21_9_i,temp_m5_21_25_r,temp_m5_21_25_i,`W8_real,`W8_imag,`W4_real,`W4_imag,`W12_real,`W12_imag);
butterfly butterfly1097 (clk,temp_m5_5_9_r,temp_m5_5_9_i,temp_m5_5_25_r,temp_m5_5_25_i,temp_m5_21_9_r,temp_m5_21_9_i,temp_m5_21_25_r,temp_m5_21_25_i,temp_b5_5_9_r,temp_b5_5_9_i,temp_b5_5_25_r,temp_b5_5_25_i,temp_b5_21_9_r,temp_b5_21_9_i,temp_b5_21_25_r,temp_b5_21_25_i);
MULT MULT1098 (clk,temp_b4_5_10_r,temp_b4_5_10_i,temp_b4_5_26_r,temp_b4_5_26_i,temp_b4_21_10_r,temp_b4_21_10_i,temp_b4_21_26_r,temp_b4_21_26_i,temp_m5_5_10_r,temp_m5_5_10_i,temp_m5_5_26_r,temp_m5_5_26_i,temp_m5_21_10_r,temp_m5_21_10_i,temp_m5_21_26_r,temp_m5_21_26_i,`W9_real,`W9_imag,`W4_real,`W4_imag,`W13_real,`W13_imag);
butterfly butterfly1098 (clk,temp_m5_5_10_r,temp_m5_5_10_i,temp_m5_5_26_r,temp_m5_5_26_i,temp_m5_21_10_r,temp_m5_21_10_i,temp_m5_21_26_r,temp_m5_21_26_i,temp_b5_5_10_r,temp_b5_5_10_i,temp_b5_5_26_r,temp_b5_5_26_i,temp_b5_21_10_r,temp_b5_21_10_i,temp_b5_21_26_r,temp_b5_21_26_i);
MULT MULT1099 (clk,temp_b4_5_11_r,temp_b4_5_11_i,temp_b4_5_27_r,temp_b4_5_27_i,temp_b4_21_11_r,temp_b4_21_11_i,temp_b4_21_27_r,temp_b4_21_27_i,temp_m5_5_11_r,temp_m5_5_11_i,temp_m5_5_27_r,temp_m5_5_27_i,temp_m5_21_11_r,temp_m5_21_11_i,temp_m5_21_27_r,temp_m5_21_27_i,`W10_real,`W10_imag,`W4_real,`W4_imag,`W14_real,`W14_imag);
butterfly butterfly1099 (clk,temp_m5_5_11_r,temp_m5_5_11_i,temp_m5_5_27_r,temp_m5_5_27_i,temp_m5_21_11_r,temp_m5_21_11_i,temp_m5_21_27_r,temp_m5_21_27_i,temp_b5_5_11_r,temp_b5_5_11_i,temp_b5_5_27_r,temp_b5_5_27_i,temp_b5_21_11_r,temp_b5_21_11_i,temp_b5_21_27_r,temp_b5_21_27_i);
MULT MULT1100 (clk,temp_b4_5_12_r,temp_b4_5_12_i,temp_b4_5_28_r,temp_b4_5_28_i,temp_b4_21_12_r,temp_b4_21_12_i,temp_b4_21_28_r,temp_b4_21_28_i,temp_m5_5_12_r,temp_m5_5_12_i,temp_m5_5_28_r,temp_m5_5_28_i,temp_m5_21_12_r,temp_m5_21_12_i,temp_m5_21_28_r,temp_m5_21_28_i,`W11_real,`W11_imag,`W4_real,`W4_imag,`W15_real,`W15_imag);
butterfly butterfly1100 (clk,temp_m5_5_12_r,temp_m5_5_12_i,temp_m5_5_28_r,temp_m5_5_28_i,temp_m5_21_12_r,temp_m5_21_12_i,temp_m5_21_28_r,temp_m5_21_28_i,temp_b5_5_12_r,temp_b5_5_12_i,temp_b5_5_28_r,temp_b5_5_28_i,temp_b5_21_12_r,temp_b5_21_12_i,temp_b5_21_28_r,temp_b5_21_28_i);
MULT MULT1101 (clk,temp_b4_5_13_r,temp_b4_5_13_i,temp_b4_5_29_r,temp_b4_5_29_i,temp_b4_21_13_r,temp_b4_21_13_i,temp_b4_21_29_r,temp_b4_21_29_i,temp_m5_5_13_r,temp_m5_5_13_i,temp_m5_5_29_r,temp_m5_5_29_i,temp_m5_21_13_r,temp_m5_21_13_i,temp_m5_21_29_r,temp_m5_21_29_i,`W12_real,`W12_imag,`W4_real,`W4_imag,`W16_real,`W16_imag);
butterfly butterfly1101 (clk,temp_m5_5_13_r,temp_m5_5_13_i,temp_m5_5_29_r,temp_m5_5_29_i,temp_m5_21_13_r,temp_m5_21_13_i,temp_m5_21_29_r,temp_m5_21_29_i,temp_b5_5_13_r,temp_b5_5_13_i,temp_b5_5_29_r,temp_b5_5_29_i,temp_b5_21_13_r,temp_b5_21_13_i,temp_b5_21_29_r,temp_b5_21_29_i);
MULT MULT1102 (clk,temp_b4_5_14_r,temp_b4_5_14_i,temp_b4_5_30_r,temp_b4_5_30_i,temp_b4_21_14_r,temp_b4_21_14_i,temp_b4_21_30_r,temp_b4_21_30_i,temp_m5_5_14_r,temp_m5_5_14_i,temp_m5_5_30_r,temp_m5_5_30_i,temp_m5_21_14_r,temp_m5_21_14_i,temp_m5_21_30_r,temp_m5_21_30_i,`W13_real,`W13_imag,`W4_real,`W4_imag,`W17_real,`W17_imag);
butterfly butterfly1102 (clk,temp_m5_5_14_r,temp_m5_5_14_i,temp_m5_5_30_r,temp_m5_5_30_i,temp_m5_21_14_r,temp_m5_21_14_i,temp_m5_21_30_r,temp_m5_21_30_i,temp_b5_5_14_r,temp_b5_5_14_i,temp_b5_5_30_r,temp_b5_5_30_i,temp_b5_21_14_r,temp_b5_21_14_i,temp_b5_21_30_r,temp_b5_21_30_i);
MULT MULT1103 (clk,temp_b4_5_15_r,temp_b4_5_15_i,temp_b4_5_31_r,temp_b4_5_31_i,temp_b4_21_15_r,temp_b4_21_15_i,temp_b4_21_31_r,temp_b4_21_31_i,temp_m5_5_15_r,temp_m5_5_15_i,temp_m5_5_31_r,temp_m5_5_31_i,temp_m5_21_15_r,temp_m5_21_15_i,temp_m5_21_31_r,temp_m5_21_31_i,`W14_real,`W14_imag,`W4_real,`W4_imag,`W18_real,`W18_imag);
butterfly butterfly1103 (clk,temp_m5_5_15_r,temp_m5_5_15_i,temp_m5_5_31_r,temp_m5_5_31_i,temp_m5_21_15_r,temp_m5_21_15_i,temp_m5_21_31_r,temp_m5_21_31_i,temp_b5_5_15_r,temp_b5_5_15_i,temp_b5_5_31_r,temp_b5_5_31_i,temp_b5_21_15_r,temp_b5_21_15_i,temp_b5_21_31_r,temp_b5_21_31_i);
MULT MULT1104 (clk,temp_b4_5_16_r,temp_b4_5_16_i,temp_b4_5_32_r,temp_b4_5_32_i,temp_b4_21_16_r,temp_b4_21_16_i,temp_b4_21_32_r,temp_b4_21_32_i,temp_m5_5_16_r,temp_m5_5_16_i,temp_m5_5_32_r,temp_m5_5_32_i,temp_m5_21_16_r,temp_m5_21_16_i,temp_m5_21_32_r,temp_m5_21_32_i,`W15_real,`W15_imag,`W4_real,`W4_imag,`W19_real,`W19_imag);
butterfly butterfly1104 (clk,temp_m5_5_16_r,temp_m5_5_16_i,temp_m5_5_32_r,temp_m5_5_32_i,temp_m5_21_16_r,temp_m5_21_16_i,temp_m5_21_32_r,temp_m5_21_32_i,temp_b5_5_16_r,temp_b5_5_16_i,temp_b5_5_32_r,temp_b5_5_32_i,temp_b5_21_16_r,temp_b5_21_16_i,temp_b5_21_32_r,temp_b5_21_32_i);
MULT MULT1105 (clk,temp_b4_6_1_r,temp_b4_6_1_i,temp_b4_6_17_r,temp_b4_6_17_i,temp_b4_22_1_r,temp_b4_22_1_i,temp_b4_22_17_r,temp_b4_22_17_i,temp_m5_6_1_r,temp_m5_6_1_i,temp_m5_6_17_r,temp_m5_6_17_i,temp_m5_22_1_r,temp_m5_22_1_i,temp_m5_22_17_r,temp_m5_22_17_i,`W0_real,`W0_imag,`W5_real,`W5_imag,`W5_real,`W5_imag);
butterfly butterfly1105 (clk,temp_m5_6_1_r,temp_m5_6_1_i,temp_m5_6_17_r,temp_m5_6_17_i,temp_m5_22_1_r,temp_m5_22_1_i,temp_m5_22_17_r,temp_m5_22_17_i,temp_b5_6_1_r,temp_b5_6_1_i,temp_b5_6_17_r,temp_b5_6_17_i,temp_b5_22_1_r,temp_b5_22_1_i,temp_b5_22_17_r,temp_b5_22_17_i);
MULT MULT1106 (clk,temp_b4_6_2_r,temp_b4_6_2_i,temp_b4_6_18_r,temp_b4_6_18_i,temp_b4_22_2_r,temp_b4_22_2_i,temp_b4_22_18_r,temp_b4_22_18_i,temp_m5_6_2_r,temp_m5_6_2_i,temp_m5_6_18_r,temp_m5_6_18_i,temp_m5_22_2_r,temp_m5_22_2_i,temp_m5_22_18_r,temp_m5_22_18_i,`W1_real,`W1_imag,`W5_real,`W5_imag,`W6_real,`W6_imag);
butterfly butterfly1106 (clk,temp_m5_6_2_r,temp_m5_6_2_i,temp_m5_6_18_r,temp_m5_6_18_i,temp_m5_22_2_r,temp_m5_22_2_i,temp_m5_22_18_r,temp_m5_22_18_i,temp_b5_6_2_r,temp_b5_6_2_i,temp_b5_6_18_r,temp_b5_6_18_i,temp_b5_22_2_r,temp_b5_22_2_i,temp_b5_22_18_r,temp_b5_22_18_i);
MULT MULT1107 (clk,temp_b4_6_3_r,temp_b4_6_3_i,temp_b4_6_19_r,temp_b4_6_19_i,temp_b4_22_3_r,temp_b4_22_3_i,temp_b4_22_19_r,temp_b4_22_19_i,temp_m5_6_3_r,temp_m5_6_3_i,temp_m5_6_19_r,temp_m5_6_19_i,temp_m5_22_3_r,temp_m5_22_3_i,temp_m5_22_19_r,temp_m5_22_19_i,`W2_real,`W2_imag,`W5_real,`W5_imag,`W7_real,`W7_imag);
butterfly butterfly1107 (clk,temp_m5_6_3_r,temp_m5_6_3_i,temp_m5_6_19_r,temp_m5_6_19_i,temp_m5_22_3_r,temp_m5_22_3_i,temp_m5_22_19_r,temp_m5_22_19_i,temp_b5_6_3_r,temp_b5_6_3_i,temp_b5_6_19_r,temp_b5_6_19_i,temp_b5_22_3_r,temp_b5_22_3_i,temp_b5_22_19_r,temp_b5_22_19_i);
MULT MULT1108 (clk,temp_b4_6_4_r,temp_b4_6_4_i,temp_b4_6_20_r,temp_b4_6_20_i,temp_b4_22_4_r,temp_b4_22_4_i,temp_b4_22_20_r,temp_b4_22_20_i,temp_m5_6_4_r,temp_m5_6_4_i,temp_m5_6_20_r,temp_m5_6_20_i,temp_m5_22_4_r,temp_m5_22_4_i,temp_m5_22_20_r,temp_m5_22_20_i,`W3_real,`W3_imag,`W5_real,`W5_imag,`W8_real,`W8_imag);
butterfly butterfly1108 (clk,temp_m5_6_4_r,temp_m5_6_4_i,temp_m5_6_20_r,temp_m5_6_20_i,temp_m5_22_4_r,temp_m5_22_4_i,temp_m5_22_20_r,temp_m5_22_20_i,temp_b5_6_4_r,temp_b5_6_4_i,temp_b5_6_20_r,temp_b5_6_20_i,temp_b5_22_4_r,temp_b5_22_4_i,temp_b5_22_20_r,temp_b5_22_20_i);
MULT MULT1109 (clk,temp_b4_6_5_r,temp_b4_6_5_i,temp_b4_6_21_r,temp_b4_6_21_i,temp_b4_22_5_r,temp_b4_22_5_i,temp_b4_22_21_r,temp_b4_22_21_i,temp_m5_6_5_r,temp_m5_6_5_i,temp_m5_6_21_r,temp_m5_6_21_i,temp_m5_22_5_r,temp_m5_22_5_i,temp_m5_22_21_r,temp_m5_22_21_i,`W4_real,`W4_imag,`W5_real,`W5_imag,`W9_real,`W9_imag);
butterfly butterfly1109 (clk,temp_m5_6_5_r,temp_m5_6_5_i,temp_m5_6_21_r,temp_m5_6_21_i,temp_m5_22_5_r,temp_m5_22_5_i,temp_m5_22_21_r,temp_m5_22_21_i,temp_b5_6_5_r,temp_b5_6_5_i,temp_b5_6_21_r,temp_b5_6_21_i,temp_b5_22_5_r,temp_b5_22_5_i,temp_b5_22_21_r,temp_b5_22_21_i);
MULT MULT1110 (clk,temp_b4_6_6_r,temp_b4_6_6_i,temp_b4_6_22_r,temp_b4_6_22_i,temp_b4_22_6_r,temp_b4_22_6_i,temp_b4_22_22_r,temp_b4_22_22_i,temp_m5_6_6_r,temp_m5_6_6_i,temp_m5_6_22_r,temp_m5_6_22_i,temp_m5_22_6_r,temp_m5_22_6_i,temp_m5_22_22_r,temp_m5_22_22_i,`W5_real,`W5_imag,`W5_real,`W5_imag,`W10_real,`W10_imag);
butterfly butterfly1110 (clk,temp_m5_6_6_r,temp_m5_6_6_i,temp_m5_6_22_r,temp_m5_6_22_i,temp_m5_22_6_r,temp_m5_22_6_i,temp_m5_22_22_r,temp_m5_22_22_i,temp_b5_6_6_r,temp_b5_6_6_i,temp_b5_6_22_r,temp_b5_6_22_i,temp_b5_22_6_r,temp_b5_22_6_i,temp_b5_22_22_r,temp_b5_22_22_i);
MULT MULT1111 (clk,temp_b4_6_7_r,temp_b4_6_7_i,temp_b4_6_23_r,temp_b4_6_23_i,temp_b4_22_7_r,temp_b4_22_7_i,temp_b4_22_23_r,temp_b4_22_23_i,temp_m5_6_7_r,temp_m5_6_7_i,temp_m5_6_23_r,temp_m5_6_23_i,temp_m5_22_7_r,temp_m5_22_7_i,temp_m5_22_23_r,temp_m5_22_23_i,`W6_real,`W6_imag,`W5_real,`W5_imag,`W11_real,`W11_imag);
butterfly butterfly1111 (clk,temp_m5_6_7_r,temp_m5_6_7_i,temp_m5_6_23_r,temp_m5_6_23_i,temp_m5_22_7_r,temp_m5_22_7_i,temp_m5_22_23_r,temp_m5_22_23_i,temp_b5_6_7_r,temp_b5_6_7_i,temp_b5_6_23_r,temp_b5_6_23_i,temp_b5_22_7_r,temp_b5_22_7_i,temp_b5_22_23_r,temp_b5_22_23_i);
MULT MULT1112 (clk,temp_b4_6_8_r,temp_b4_6_8_i,temp_b4_6_24_r,temp_b4_6_24_i,temp_b4_22_8_r,temp_b4_22_8_i,temp_b4_22_24_r,temp_b4_22_24_i,temp_m5_6_8_r,temp_m5_6_8_i,temp_m5_6_24_r,temp_m5_6_24_i,temp_m5_22_8_r,temp_m5_22_8_i,temp_m5_22_24_r,temp_m5_22_24_i,`W7_real,`W7_imag,`W5_real,`W5_imag,`W12_real,`W12_imag);
butterfly butterfly1112 (clk,temp_m5_6_8_r,temp_m5_6_8_i,temp_m5_6_24_r,temp_m5_6_24_i,temp_m5_22_8_r,temp_m5_22_8_i,temp_m5_22_24_r,temp_m5_22_24_i,temp_b5_6_8_r,temp_b5_6_8_i,temp_b5_6_24_r,temp_b5_6_24_i,temp_b5_22_8_r,temp_b5_22_8_i,temp_b5_22_24_r,temp_b5_22_24_i);
MULT MULT1113 (clk,temp_b4_6_9_r,temp_b4_6_9_i,temp_b4_6_25_r,temp_b4_6_25_i,temp_b4_22_9_r,temp_b4_22_9_i,temp_b4_22_25_r,temp_b4_22_25_i,temp_m5_6_9_r,temp_m5_6_9_i,temp_m5_6_25_r,temp_m5_6_25_i,temp_m5_22_9_r,temp_m5_22_9_i,temp_m5_22_25_r,temp_m5_22_25_i,`W8_real,`W8_imag,`W5_real,`W5_imag,`W13_real,`W13_imag);
butterfly butterfly1113 (clk,temp_m5_6_9_r,temp_m5_6_9_i,temp_m5_6_25_r,temp_m5_6_25_i,temp_m5_22_9_r,temp_m5_22_9_i,temp_m5_22_25_r,temp_m5_22_25_i,temp_b5_6_9_r,temp_b5_6_9_i,temp_b5_6_25_r,temp_b5_6_25_i,temp_b5_22_9_r,temp_b5_22_9_i,temp_b5_22_25_r,temp_b5_22_25_i);
MULT MULT1114 (clk,temp_b4_6_10_r,temp_b4_6_10_i,temp_b4_6_26_r,temp_b4_6_26_i,temp_b4_22_10_r,temp_b4_22_10_i,temp_b4_22_26_r,temp_b4_22_26_i,temp_m5_6_10_r,temp_m5_6_10_i,temp_m5_6_26_r,temp_m5_6_26_i,temp_m5_22_10_r,temp_m5_22_10_i,temp_m5_22_26_r,temp_m5_22_26_i,`W9_real,`W9_imag,`W5_real,`W5_imag,`W14_real,`W14_imag);
butterfly butterfly1114 (clk,temp_m5_6_10_r,temp_m5_6_10_i,temp_m5_6_26_r,temp_m5_6_26_i,temp_m5_22_10_r,temp_m5_22_10_i,temp_m5_22_26_r,temp_m5_22_26_i,temp_b5_6_10_r,temp_b5_6_10_i,temp_b5_6_26_r,temp_b5_6_26_i,temp_b5_22_10_r,temp_b5_22_10_i,temp_b5_22_26_r,temp_b5_22_26_i);
MULT MULT1115 (clk,temp_b4_6_11_r,temp_b4_6_11_i,temp_b4_6_27_r,temp_b4_6_27_i,temp_b4_22_11_r,temp_b4_22_11_i,temp_b4_22_27_r,temp_b4_22_27_i,temp_m5_6_11_r,temp_m5_6_11_i,temp_m5_6_27_r,temp_m5_6_27_i,temp_m5_22_11_r,temp_m5_22_11_i,temp_m5_22_27_r,temp_m5_22_27_i,`W10_real,`W10_imag,`W5_real,`W5_imag,`W15_real,`W15_imag);
butterfly butterfly1115 (clk,temp_m5_6_11_r,temp_m5_6_11_i,temp_m5_6_27_r,temp_m5_6_27_i,temp_m5_22_11_r,temp_m5_22_11_i,temp_m5_22_27_r,temp_m5_22_27_i,temp_b5_6_11_r,temp_b5_6_11_i,temp_b5_6_27_r,temp_b5_6_27_i,temp_b5_22_11_r,temp_b5_22_11_i,temp_b5_22_27_r,temp_b5_22_27_i);
MULT MULT1116 (clk,temp_b4_6_12_r,temp_b4_6_12_i,temp_b4_6_28_r,temp_b4_6_28_i,temp_b4_22_12_r,temp_b4_22_12_i,temp_b4_22_28_r,temp_b4_22_28_i,temp_m5_6_12_r,temp_m5_6_12_i,temp_m5_6_28_r,temp_m5_6_28_i,temp_m5_22_12_r,temp_m5_22_12_i,temp_m5_22_28_r,temp_m5_22_28_i,`W11_real,`W11_imag,`W5_real,`W5_imag,`W16_real,`W16_imag);
butterfly butterfly1116 (clk,temp_m5_6_12_r,temp_m5_6_12_i,temp_m5_6_28_r,temp_m5_6_28_i,temp_m5_22_12_r,temp_m5_22_12_i,temp_m5_22_28_r,temp_m5_22_28_i,temp_b5_6_12_r,temp_b5_6_12_i,temp_b5_6_28_r,temp_b5_6_28_i,temp_b5_22_12_r,temp_b5_22_12_i,temp_b5_22_28_r,temp_b5_22_28_i);
MULT MULT1117 (clk,temp_b4_6_13_r,temp_b4_6_13_i,temp_b4_6_29_r,temp_b4_6_29_i,temp_b4_22_13_r,temp_b4_22_13_i,temp_b4_22_29_r,temp_b4_22_29_i,temp_m5_6_13_r,temp_m5_6_13_i,temp_m5_6_29_r,temp_m5_6_29_i,temp_m5_22_13_r,temp_m5_22_13_i,temp_m5_22_29_r,temp_m5_22_29_i,`W12_real,`W12_imag,`W5_real,`W5_imag,`W17_real,`W17_imag);
butterfly butterfly1117 (clk,temp_m5_6_13_r,temp_m5_6_13_i,temp_m5_6_29_r,temp_m5_6_29_i,temp_m5_22_13_r,temp_m5_22_13_i,temp_m5_22_29_r,temp_m5_22_29_i,temp_b5_6_13_r,temp_b5_6_13_i,temp_b5_6_29_r,temp_b5_6_29_i,temp_b5_22_13_r,temp_b5_22_13_i,temp_b5_22_29_r,temp_b5_22_29_i);
MULT MULT1118 (clk,temp_b4_6_14_r,temp_b4_6_14_i,temp_b4_6_30_r,temp_b4_6_30_i,temp_b4_22_14_r,temp_b4_22_14_i,temp_b4_22_30_r,temp_b4_22_30_i,temp_m5_6_14_r,temp_m5_6_14_i,temp_m5_6_30_r,temp_m5_6_30_i,temp_m5_22_14_r,temp_m5_22_14_i,temp_m5_22_30_r,temp_m5_22_30_i,`W13_real,`W13_imag,`W5_real,`W5_imag,`W18_real,`W18_imag);
butterfly butterfly1118 (clk,temp_m5_6_14_r,temp_m5_6_14_i,temp_m5_6_30_r,temp_m5_6_30_i,temp_m5_22_14_r,temp_m5_22_14_i,temp_m5_22_30_r,temp_m5_22_30_i,temp_b5_6_14_r,temp_b5_6_14_i,temp_b5_6_30_r,temp_b5_6_30_i,temp_b5_22_14_r,temp_b5_22_14_i,temp_b5_22_30_r,temp_b5_22_30_i);
MULT MULT1119 (clk,temp_b4_6_15_r,temp_b4_6_15_i,temp_b4_6_31_r,temp_b4_6_31_i,temp_b4_22_15_r,temp_b4_22_15_i,temp_b4_22_31_r,temp_b4_22_31_i,temp_m5_6_15_r,temp_m5_6_15_i,temp_m5_6_31_r,temp_m5_6_31_i,temp_m5_22_15_r,temp_m5_22_15_i,temp_m5_22_31_r,temp_m5_22_31_i,`W14_real,`W14_imag,`W5_real,`W5_imag,`W19_real,`W19_imag);
butterfly butterfly1119 (clk,temp_m5_6_15_r,temp_m5_6_15_i,temp_m5_6_31_r,temp_m5_6_31_i,temp_m5_22_15_r,temp_m5_22_15_i,temp_m5_22_31_r,temp_m5_22_31_i,temp_b5_6_15_r,temp_b5_6_15_i,temp_b5_6_31_r,temp_b5_6_31_i,temp_b5_22_15_r,temp_b5_22_15_i,temp_b5_22_31_r,temp_b5_22_31_i);
MULT MULT1120 (clk,temp_b4_6_16_r,temp_b4_6_16_i,temp_b4_6_32_r,temp_b4_6_32_i,temp_b4_22_16_r,temp_b4_22_16_i,temp_b4_22_32_r,temp_b4_22_32_i,temp_m5_6_16_r,temp_m5_6_16_i,temp_m5_6_32_r,temp_m5_6_32_i,temp_m5_22_16_r,temp_m5_22_16_i,temp_m5_22_32_r,temp_m5_22_32_i,`W15_real,`W15_imag,`W5_real,`W5_imag,`W20_real,`W20_imag);
butterfly butterfly1120 (clk,temp_m5_6_16_r,temp_m5_6_16_i,temp_m5_6_32_r,temp_m5_6_32_i,temp_m5_22_16_r,temp_m5_22_16_i,temp_m5_22_32_r,temp_m5_22_32_i,temp_b5_6_16_r,temp_b5_6_16_i,temp_b5_6_32_r,temp_b5_6_32_i,temp_b5_22_16_r,temp_b5_22_16_i,temp_b5_22_32_r,temp_b5_22_32_i);
MULT MULT1121 (clk,temp_b4_7_1_r,temp_b4_7_1_i,temp_b4_7_17_r,temp_b4_7_17_i,temp_b4_23_1_r,temp_b4_23_1_i,temp_b4_23_17_r,temp_b4_23_17_i,temp_m5_7_1_r,temp_m5_7_1_i,temp_m5_7_17_r,temp_m5_7_17_i,temp_m5_23_1_r,temp_m5_23_1_i,temp_m5_23_17_r,temp_m5_23_17_i,`W0_real,`W0_imag,`W6_real,`W6_imag,`W6_real,`W6_imag);
butterfly butterfly1121 (clk,temp_m5_7_1_r,temp_m5_7_1_i,temp_m5_7_17_r,temp_m5_7_17_i,temp_m5_23_1_r,temp_m5_23_1_i,temp_m5_23_17_r,temp_m5_23_17_i,temp_b5_7_1_r,temp_b5_7_1_i,temp_b5_7_17_r,temp_b5_7_17_i,temp_b5_23_1_r,temp_b5_23_1_i,temp_b5_23_17_r,temp_b5_23_17_i);
MULT MULT1122 (clk,temp_b4_7_2_r,temp_b4_7_2_i,temp_b4_7_18_r,temp_b4_7_18_i,temp_b4_23_2_r,temp_b4_23_2_i,temp_b4_23_18_r,temp_b4_23_18_i,temp_m5_7_2_r,temp_m5_7_2_i,temp_m5_7_18_r,temp_m5_7_18_i,temp_m5_23_2_r,temp_m5_23_2_i,temp_m5_23_18_r,temp_m5_23_18_i,`W1_real,`W1_imag,`W6_real,`W6_imag,`W7_real,`W7_imag);
butterfly butterfly1122 (clk,temp_m5_7_2_r,temp_m5_7_2_i,temp_m5_7_18_r,temp_m5_7_18_i,temp_m5_23_2_r,temp_m5_23_2_i,temp_m5_23_18_r,temp_m5_23_18_i,temp_b5_7_2_r,temp_b5_7_2_i,temp_b5_7_18_r,temp_b5_7_18_i,temp_b5_23_2_r,temp_b5_23_2_i,temp_b5_23_18_r,temp_b5_23_18_i);
MULT MULT1123 (clk,temp_b4_7_3_r,temp_b4_7_3_i,temp_b4_7_19_r,temp_b4_7_19_i,temp_b4_23_3_r,temp_b4_23_3_i,temp_b4_23_19_r,temp_b4_23_19_i,temp_m5_7_3_r,temp_m5_7_3_i,temp_m5_7_19_r,temp_m5_7_19_i,temp_m5_23_3_r,temp_m5_23_3_i,temp_m5_23_19_r,temp_m5_23_19_i,`W2_real,`W2_imag,`W6_real,`W6_imag,`W8_real,`W8_imag);
butterfly butterfly1123 (clk,temp_m5_7_3_r,temp_m5_7_3_i,temp_m5_7_19_r,temp_m5_7_19_i,temp_m5_23_3_r,temp_m5_23_3_i,temp_m5_23_19_r,temp_m5_23_19_i,temp_b5_7_3_r,temp_b5_7_3_i,temp_b5_7_19_r,temp_b5_7_19_i,temp_b5_23_3_r,temp_b5_23_3_i,temp_b5_23_19_r,temp_b5_23_19_i);
MULT MULT1124 (clk,temp_b4_7_4_r,temp_b4_7_4_i,temp_b4_7_20_r,temp_b4_7_20_i,temp_b4_23_4_r,temp_b4_23_4_i,temp_b4_23_20_r,temp_b4_23_20_i,temp_m5_7_4_r,temp_m5_7_4_i,temp_m5_7_20_r,temp_m5_7_20_i,temp_m5_23_4_r,temp_m5_23_4_i,temp_m5_23_20_r,temp_m5_23_20_i,`W3_real,`W3_imag,`W6_real,`W6_imag,`W9_real,`W9_imag);
butterfly butterfly1124 (clk,temp_m5_7_4_r,temp_m5_7_4_i,temp_m5_7_20_r,temp_m5_7_20_i,temp_m5_23_4_r,temp_m5_23_4_i,temp_m5_23_20_r,temp_m5_23_20_i,temp_b5_7_4_r,temp_b5_7_4_i,temp_b5_7_20_r,temp_b5_7_20_i,temp_b5_23_4_r,temp_b5_23_4_i,temp_b5_23_20_r,temp_b5_23_20_i);
MULT MULT1125 (clk,temp_b4_7_5_r,temp_b4_7_5_i,temp_b4_7_21_r,temp_b4_7_21_i,temp_b4_23_5_r,temp_b4_23_5_i,temp_b4_23_21_r,temp_b4_23_21_i,temp_m5_7_5_r,temp_m5_7_5_i,temp_m5_7_21_r,temp_m5_7_21_i,temp_m5_23_5_r,temp_m5_23_5_i,temp_m5_23_21_r,temp_m5_23_21_i,`W4_real,`W4_imag,`W6_real,`W6_imag,`W10_real,`W10_imag);
butterfly butterfly1125 (clk,temp_m5_7_5_r,temp_m5_7_5_i,temp_m5_7_21_r,temp_m5_7_21_i,temp_m5_23_5_r,temp_m5_23_5_i,temp_m5_23_21_r,temp_m5_23_21_i,temp_b5_7_5_r,temp_b5_7_5_i,temp_b5_7_21_r,temp_b5_7_21_i,temp_b5_23_5_r,temp_b5_23_5_i,temp_b5_23_21_r,temp_b5_23_21_i);
MULT MULT1126 (clk,temp_b4_7_6_r,temp_b4_7_6_i,temp_b4_7_22_r,temp_b4_7_22_i,temp_b4_23_6_r,temp_b4_23_6_i,temp_b4_23_22_r,temp_b4_23_22_i,temp_m5_7_6_r,temp_m5_7_6_i,temp_m5_7_22_r,temp_m5_7_22_i,temp_m5_23_6_r,temp_m5_23_6_i,temp_m5_23_22_r,temp_m5_23_22_i,`W5_real,`W5_imag,`W6_real,`W6_imag,`W11_real,`W11_imag);
butterfly butterfly1126 (clk,temp_m5_7_6_r,temp_m5_7_6_i,temp_m5_7_22_r,temp_m5_7_22_i,temp_m5_23_6_r,temp_m5_23_6_i,temp_m5_23_22_r,temp_m5_23_22_i,temp_b5_7_6_r,temp_b5_7_6_i,temp_b5_7_22_r,temp_b5_7_22_i,temp_b5_23_6_r,temp_b5_23_6_i,temp_b5_23_22_r,temp_b5_23_22_i);
MULT MULT1127 (clk,temp_b4_7_7_r,temp_b4_7_7_i,temp_b4_7_23_r,temp_b4_7_23_i,temp_b4_23_7_r,temp_b4_23_7_i,temp_b4_23_23_r,temp_b4_23_23_i,temp_m5_7_7_r,temp_m5_7_7_i,temp_m5_7_23_r,temp_m5_7_23_i,temp_m5_23_7_r,temp_m5_23_7_i,temp_m5_23_23_r,temp_m5_23_23_i,`W6_real,`W6_imag,`W6_real,`W6_imag,`W12_real,`W12_imag);
butterfly butterfly1127 (clk,temp_m5_7_7_r,temp_m5_7_7_i,temp_m5_7_23_r,temp_m5_7_23_i,temp_m5_23_7_r,temp_m5_23_7_i,temp_m5_23_23_r,temp_m5_23_23_i,temp_b5_7_7_r,temp_b5_7_7_i,temp_b5_7_23_r,temp_b5_7_23_i,temp_b5_23_7_r,temp_b5_23_7_i,temp_b5_23_23_r,temp_b5_23_23_i);
MULT MULT1128 (clk,temp_b4_7_8_r,temp_b4_7_8_i,temp_b4_7_24_r,temp_b4_7_24_i,temp_b4_23_8_r,temp_b4_23_8_i,temp_b4_23_24_r,temp_b4_23_24_i,temp_m5_7_8_r,temp_m5_7_8_i,temp_m5_7_24_r,temp_m5_7_24_i,temp_m5_23_8_r,temp_m5_23_8_i,temp_m5_23_24_r,temp_m5_23_24_i,`W7_real,`W7_imag,`W6_real,`W6_imag,`W13_real,`W13_imag);
butterfly butterfly1128 (clk,temp_m5_7_8_r,temp_m5_7_8_i,temp_m5_7_24_r,temp_m5_7_24_i,temp_m5_23_8_r,temp_m5_23_8_i,temp_m5_23_24_r,temp_m5_23_24_i,temp_b5_7_8_r,temp_b5_7_8_i,temp_b5_7_24_r,temp_b5_7_24_i,temp_b5_23_8_r,temp_b5_23_8_i,temp_b5_23_24_r,temp_b5_23_24_i);
MULT MULT1129 (clk,temp_b4_7_9_r,temp_b4_7_9_i,temp_b4_7_25_r,temp_b4_7_25_i,temp_b4_23_9_r,temp_b4_23_9_i,temp_b4_23_25_r,temp_b4_23_25_i,temp_m5_7_9_r,temp_m5_7_9_i,temp_m5_7_25_r,temp_m5_7_25_i,temp_m5_23_9_r,temp_m5_23_9_i,temp_m5_23_25_r,temp_m5_23_25_i,`W8_real,`W8_imag,`W6_real,`W6_imag,`W14_real,`W14_imag);
butterfly butterfly1129 (clk,temp_m5_7_9_r,temp_m5_7_9_i,temp_m5_7_25_r,temp_m5_7_25_i,temp_m5_23_9_r,temp_m5_23_9_i,temp_m5_23_25_r,temp_m5_23_25_i,temp_b5_7_9_r,temp_b5_7_9_i,temp_b5_7_25_r,temp_b5_7_25_i,temp_b5_23_9_r,temp_b5_23_9_i,temp_b5_23_25_r,temp_b5_23_25_i);
MULT MULT1130 (clk,temp_b4_7_10_r,temp_b4_7_10_i,temp_b4_7_26_r,temp_b4_7_26_i,temp_b4_23_10_r,temp_b4_23_10_i,temp_b4_23_26_r,temp_b4_23_26_i,temp_m5_7_10_r,temp_m5_7_10_i,temp_m5_7_26_r,temp_m5_7_26_i,temp_m5_23_10_r,temp_m5_23_10_i,temp_m5_23_26_r,temp_m5_23_26_i,`W9_real,`W9_imag,`W6_real,`W6_imag,`W15_real,`W15_imag);
butterfly butterfly1130 (clk,temp_m5_7_10_r,temp_m5_7_10_i,temp_m5_7_26_r,temp_m5_7_26_i,temp_m5_23_10_r,temp_m5_23_10_i,temp_m5_23_26_r,temp_m5_23_26_i,temp_b5_7_10_r,temp_b5_7_10_i,temp_b5_7_26_r,temp_b5_7_26_i,temp_b5_23_10_r,temp_b5_23_10_i,temp_b5_23_26_r,temp_b5_23_26_i);
MULT MULT1131 (clk,temp_b4_7_11_r,temp_b4_7_11_i,temp_b4_7_27_r,temp_b4_7_27_i,temp_b4_23_11_r,temp_b4_23_11_i,temp_b4_23_27_r,temp_b4_23_27_i,temp_m5_7_11_r,temp_m5_7_11_i,temp_m5_7_27_r,temp_m5_7_27_i,temp_m5_23_11_r,temp_m5_23_11_i,temp_m5_23_27_r,temp_m5_23_27_i,`W10_real,`W10_imag,`W6_real,`W6_imag,`W16_real,`W16_imag);
butterfly butterfly1131 (clk,temp_m5_7_11_r,temp_m5_7_11_i,temp_m5_7_27_r,temp_m5_7_27_i,temp_m5_23_11_r,temp_m5_23_11_i,temp_m5_23_27_r,temp_m5_23_27_i,temp_b5_7_11_r,temp_b5_7_11_i,temp_b5_7_27_r,temp_b5_7_27_i,temp_b5_23_11_r,temp_b5_23_11_i,temp_b5_23_27_r,temp_b5_23_27_i);
MULT MULT1132 (clk,temp_b4_7_12_r,temp_b4_7_12_i,temp_b4_7_28_r,temp_b4_7_28_i,temp_b4_23_12_r,temp_b4_23_12_i,temp_b4_23_28_r,temp_b4_23_28_i,temp_m5_7_12_r,temp_m5_7_12_i,temp_m5_7_28_r,temp_m5_7_28_i,temp_m5_23_12_r,temp_m5_23_12_i,temp_m5_23_28_r,temp_m5_23_28_i,`W11_real,`W11_imag,`W6_real,`W6_imag,`W17_real,`W17_imag);
butterfly butterfly1132 (clk,temp_m5_7_12_r,temp_m5_7_12_i,temp_m5_7_28_r,temp_m5_7_28_i,temp_m5_23_12_r,temp_m5_23_12_i,temp_m5_23_28_r,temp_m5_23_28_i,temp_b5_7_12_r,temp_b5_7_12_i,temp_b5_7_28_r,temp_b5_7_28_i,temp_b5_23_12_r,temp_b5_23_12_i,temp_b5_23_28_r,temp_b5_23_28_i);
MULT MULT1133 (clk,temp_b4_7_13_r,temp_b4_7_13_i,temp_b4_7_29_r,temp_b4_7_29_i,temp_b4_23_13_r,temp_b4_23_13_i,temp_b4_23_29_r,temp_b4_23_29_i,temp_m5_7_13_r,temp_m5_7_13_i,temp_m5_7_29_r,temp_m5_7_29_i,temp_m5_23_13_r,temp_m5_23_13_i,temp_m5_23_29_r,temp_m5_23_29_i,`W12_real,`W12_imag,`W6_real,`W6_imag,`W18_real,`W18_imag);
butterfly butterfly1133 (clk,temp_m5_7_13_r,temp_m5_7_13_i,temp_m5_7_29_r,temp_m5_7_29_i,temp_m5_23_13_r,temp_m5_23_13_i,temp_m5_23_29_r,temp_m5_23_29_i,temp_b5_7_13_r,temp_b5_7_13_i,temp_b5_7_29_r,temp_b5_7_29_i,temp_b5_23_13_r,temp_b5_23_13_i,temp_b5_23_29_r,temp_b5_23_29_i);
MULT MULT1134 (clk,temp_b4_7_14_r,temp_b4_7_14_i,temp_b4_7_30_r,temp_b4_7_30_i,temp_b4_23_14_r,temp_b4_23_14_i,temp_b4_23_30_r,temp_b4_23_30_i,temp_m5_7_14_r,temp_m5_7_14_i,temp_m5_7_30_r,temp_m5_7_30_i,temp_m5_23_14_r,temp_m5_23_14_i,temp_m5_23_30_r,temp_m5_23_30_i,`W13_real,`W13_imag,`W6_real,`W6_imag,`W19_real,`W19_imag);
butterfly butterfly1134 (clk,temp_m5_7_14_r,temp_m5_7_14_i,temp_m5_7_30_r,temp_m5_7_30_i,temp_m5_23_14_r,temp_m5_23_14_i,temp_m5_23_30_r,temp_m5_23_30_i,temp_b5_7_14_r,temp_b5_7_14_i,temp_b5_7_30_r,temp_b5_7_30_i,temp_b5_23_14_r,temp_b5_23_14_i,temp_b5_23_30_r,temp_b5_23_30_i);
MULT MULT1135 (clk,temp_b4_7_15_r,temp_b4_7_15_i,temp_b4_7_31_r,temp_b4_7_31_i,temp_b4_23_15_r,temp_b4_23_15_i,temp_b4_23_31_r,temp_b4_23_31_i,temp_m5_7_15_r,temp_m5_7_15_i,temp_m5_7_31_r,temp_m5_7_31_i,temp_m5_23_15_r,temp_m5_23_15_i,temp_m5_23_31_r,temp_m5_23_31_i,`W14_real,`W14_imag,`W6_real,`W6_imag,`W20_real,`W20_imag);
butterfly butterfly1135 (clk,temp_m5_7_15_r,temp_m5_7_15_i,temp_m5_7_31_r,temp_m5_7_31_i,temp_m5_23_15_r,temp_m5_23_15_i,temp_m5_23_31_r,temp_m5_23_31_i,temp_b5_7_15_r,temp_b5_7_15_i,temp_b5_7_31_r,temp_b5_7_31_i,temp_b5_23_15_r,temp_b5_23_15_i,temp_b5_23_31_r,temp_b5_23_31_i);
MULT MULT1136 (clk,temp_b4_7_16_r,temp_b4_7_16_i,temp_b4_7_32_r,temp_b4_7_32_i,temp_b4_23_16_r,temp_b4_23_16_i,temp_b4_23_32_r,temp_b4_23_32_i,temp_m5_7_16_r,temp_m5_7_16_i,temp_m5_7_32_r,temp_m5_7_32_i,temp_m5_23_16_r,temp_m5_23_16_i,temp_m5_23_32_r,temp_m5_23_32_i,`W15_real,`W15_imag,`W6_real,`W6_imag,`W21_real,`W21_imag);
butterfly butterfly1136 (clk,temp_m5_7_16_r,temp_m5_7_16_i,temp_m5_7_32_r,temp_m5_7_32_i,temp_m5_23_16_r,temp_m5_23_16_i,temp_m5_23_32_r,temp_m5_23_32_i,temp_b5_7_16_r,temp_b5_7_16_i,temp_b5_7_32_r,temp_b5_7_32_i,temp_b5_23_16_r,temp_b5_23_16_i,temp_b5_23_32_r,temp_b5_23_32_i);
MULT MULT1137 (clk,temp_b4_8_1_r,temp_b4_8_1_i,temp_b4_8_17_r,temp_b4_8_17_i,temp_b4_24_1_r,temp_b4_24_1_i,temp_b4_24_17_r,temp_b4_24_17_i,temp_m5_8_1_r,temp_m5_8_1_i,temp_m5_8_17_r,temp_m5_8_17_i,temp_m5_24_1_r,temp_m5_24_1_i,temp_m5_24_17_r,temp_m5_24_17_i,`W0_real,`W0_imag,`W7_real,`W7_imag,`W7_real,`W7_imag);
butterfly butterfly1137 (clk,temp_m5_8_1_r,temp_m5_8_1_i,temp_m5_8_17_r,temp_m5_8_17_i,temp_m5_24_1_r,temp_m5_24_1_i,temp_m5_24_17_r,temp_m5_24_17_i,temp_b5_8_1_r,temp_b5_8_1_i,temp_b5_8_17_r,temp_b5_8_17_i,temp_b5_24_1_r,temp_b5_24_1_i,temp_b5_24_17_r,temp_b5_24_17_i);
MULT MULT1138 (clk,temp_b4_8_2_r,temp_b4_8_2_i,temp_b4_8_18_r,temp_b4_8_18_i,temp_b4_24_2_r,temp_b4_24_2_i,temp_b4_24_18_r,temp_b4_24_18_i,temp_m5_8_2_r,temp_m5_8_2_i,temp_m5_8_18_r,temp_m5_8_18_i,temp_m5_24_2_r,temp_m5_24_2_i,temp_m5_24_18_r,temp_m5_24_18_i,`W1_real,`W1_imag,`W7_real,`W7_imag,`W8_real,`W8_imag);
butterfly butterfly1138 (clk,temp_m5_8_2_r,temp_m5_8_2_i,temp_m5_8_18_r,temp_m5_8_18_i,temp_m5_24_2_r,temp_m5_24_2_i,temp_m5_24_18_r,temp_m5_24_18_i,temp_b5_8_2_r,temp_b5_8_2_i,temp_b5_8_18_r,temp_b5_8_18_i,temp_b5_24_2_r,temp_b5_24_2_i,temp_b5_24_18_r,temp_b5_24_18_i);
MULT MULT1139 (clk,temp_b4_8_3_r,temp_b4_8_3_i,temp_b4_8_19_r,temp_b4_8_19_i,temp_b4_24_3_r,temp_b4_24_3_i,temp_b4_24_19_r,temp_b4_24_19_i,temp_m5_8_3_r,temp_m5_8_3_i,temp_m5_8_19_r,temp_m5_8_19_i,temp_m5_24_3_r,temp_m5_24_3_i,temp_m5_24_19_r,temp_m5_24_19_i,`W2_real,`W2_imag,`W7_real,`W7_imag,`W9_real,`W9_imag);
butterfly butterfly1139 (clk,temp_m5_8_3_r,temp_m5_8_3_i,temp_m5_8_19_r,temp_m5_8_19_i,temp_m5_24_3_r,temp_m5_24_3_i,temp_m5_24_19_r,temp_m5_24_19_i,temp_b5_8_3_r,temp_b5_8_3_i,temp_b5_8_19_r,temp_b5_8_19_i,temp_b5_24_3_r,temp_b5_24_3_i,temp_b5_24_19_r,temp_b5_24_19_i);
MULT MULT1140 (clk,temp_b4_8_4_r,temp_b4_8_4_i,temp_b4_8_20_r,temp_b4_8_20_i,temp_b4_24_4_r,temp_b4_24_4_i,temp_b4_24_20_r,temp_b4_24_20_i,temp_m5_8_4_r,temp_m5_8_4_i,temp_m5_8_20_r,temp_m5_8_20_i,temp_m5_24_4_r,temp_m5_24_4_i,temp_m5_24_20_r,temp_m5_24_20_i,`W3_real,`W3_imag,`W7_real,`W7_imag,`W10_real,`W10_imag);
butterfly butterfly1140 (clk,temp_m5_8_4_r,temp_m5_8_4_i,temp_m5_8_20_r,temp_m5_8_20_i,temp_m5_24_4_r,temp_m5_24_4_i,temp_m5_24_20_r,temp_m5_24_20_i,temp_b5_8_4_r,temp_b5_8_4_i,temp_b5_8_20_r,temp_b5_8_20_i,temp_b5_24_4_r,temp_b5_24_4_i,temp_b5_24_20_r,temp_b5_24_20_i);
MULT MULT1141 (clk,temp_b4_8_5_r,temp_b4_8_5_i,temp_b4_8_21_r,temp_b4_8_21_i,temp_b4_24_5_r,temp_b4_24_5_i,temp_b4_24_21_r,temp_b4_24_21_i,temp_m5_8_5_r,temp_m5_8_5_i,temp_m5_8_21_r,temp_m5_8_21_i,temp_m5_24_5_r,temp_m5_24_5_i,temp_m5_24_21_r,temp_m5_24_21_i,`W4_real,`W4_imag,`W7_real,`W7_imag,`W11_real,`W11_imag);
butterfly butterfly1141 (clk,temp_m5_8_5_r,temp_m5_8_5_i,temp_m5_8_21_r,temp_m5_8_21_i,temp_m5_24_5_r,temp_m5_24_5_i,temp_m5_24_21_r,temp_m5_24_21_i,temp_b5_8_5_r,temp_b5_8_5_i,temp_b5_8_21_r,temp_b5_8_21_i,temp_b5_24_5_r,temp_b5_24_5_i,temp_b5_24_21_r,temp_b5_24_21_i);
MULT MULT1142 (clk,temp_b4_8_6_r,temp_b4_8_6_i,temp_b4_8_22_r,temp_b4_8_22_i,temp_b4_24_6_r,temp_b4_24_6_i,temp_b4_24_22_r,temp_b4_24_22_i,temp_m5_8_6_r,temp_m5_8_6_i,temp_m5_8_22_r,temp_m5_8_22_i,temp_m5_24_6_r,temp_m5_24_6_i,temp_m5_24_22_r,temp_m5_24_22_i,`W5_real,`W5_imag,`W7_real,`W7_imag,`W12_real,`W12_imag);
butterfly butterfly1142 (clk,temp_m5_8_6_r,temp_m5_8_6_i,temp_m5_8_22_r,temp_m5_8_22_i,temp_m5_24_6_r,temp_m5_24_6_i,temp_m5_24_22_r,temp_m5_24_22_i,temp_b5_8_6_r,temp_b5_8_6_i,temp_b5_8_22_r,temp_b5_8_22_i,temp_b5_24_6_r,temp_b5_24_6_i,temp_b5_24_22_r,temp_b5_24_22_i);
MULT MULT1143 (clk,temp_b4_8_7_r,temp_b4_8_7_i,temp_b4_8_23_r,temp_b4_8_23_i,temp_b4_24_7_r,temp_b4_24_7_i,temp_b4_24_23_r,temp_b4_24_23_i,temp_m5_8_7_r,temp_m5_8_7_i,temp_m5_8_23_r,temp_m5_8_23_i,temp_m5_24_7_r,temp_m5_24_7_i,temp_m5_24_23_r,temp_m5_24_23_i,`W6_real,`W6_imag,`W7_real,`W7_imag,`W13_real,`W13_imag);
butterfly butterfly1143 (clk,temp_m5_8_7_r,temp_m5_8_7_i,temp_m5_8_23_r,temp_m5_8_23_i,temp_m5_24_7_r,temp_m5_24_7_i,temp_m5_24_23_r,temp_m5_24_23_i,temp_b5_8_7_r,temp_b5_8_7_i,temp_b5_8_23_r,temp_b5_8_23_i,temp_b5_24_7_r,temp_b5_24_7_i,temp_b5_24_23_r,temp_b5_24_23_i);
MULT MULT1144 (clk,temp_b4_8_8_r,temp_b4_8_8_i,temp_b4_8_24_r,temp_b4_8_24_i,temp_b4_24_8_r,temp_b4_24_8_i,temp_b4_24_24_r,temp_b4_24_24_i,temp_m5_8_8_r,temp_m5_8_8_i,temp_m5_8_24_r,temp_m5_8_24_i,temp_m5_24_8_r,temp_m5_24_8_i,temp_m5_24_24_r,temp_m5_24_24_i,`W7_real,`W7_imag,`W7_real,`W7_imag,`W14_real,`W14_imag);
butterfly butterfly1144 (clk,temp_m5_8_8_r,temp_m5_8_8_i,temp_m5_8_24_r,temp_m5_8_24_i,temp_m5_24_8_r,temp_m5_24_8_i,temp_m5_24_24_r,temp_m5_24_24_i,temp_b5_8_8_r,temp_b5_8_8_i,temp_b5_8_24_r,temp_b5_8_24_i,temp_b5_24_8_r,temp_b5_24_8_i,temp_b5_24_24_r,temp_b5_24_24_i);
MULT MULT1145 (clk,temp_b4_8_9_r,temp_b4_8_9_i,temp_b4_8_25_r,temp_b4_8_25_i,temp_b4_24_9_r,temp_b4_24_9_i,temp_b4_24_25_r,temp_b4_24_25_i,temp_m5_8_9_r,temp_m5_8_9_i,temp_m5_8_25_r,temp_m5_8_25_i,temp_m5_24_9_r,temp_m5_24_9_i,temp_m5_24_25_r,temp_m5_24_25_i,`W8_real,`W8_imag,`W7_real,`W7_imag,`W15_real,`W15_imag);
butterfly butterfly1145 (clk,temp_m5_8_9_r,temp_m5_8_9_i,temp_m5_8_25_r,temp_m5_8_25_i,temp_m5_24_9_r,temp_m5_24_9_i,temp_m5_24_25_r,temp_m5_24_25_i,temp_b5_8_9_r,temp_b5_8_9_i,temp_b5_8_25_r,temp_b5_8_25_i,temp_b5_24_9_r,temp_b5_24_9_i,temp_b5_24_25_r,temp_b5_24_25_i);
MULT MULT1146 (clk,temp_b4_8_10_r,temp_b4_8_10_i,temp_b4_8_26_r,temp_b4_8_26_i,temp_b4_24_10_r,temp_b4_24_10_i,temp_b4_24_26_r,temp_b4_24_26_i,temp_m5_8_10_r,temp_m5_8_10_i,temp_m5_8_26_r,temp_m5_8_26_i,temp_m5_24_10_r,temp_m5_24_10_i,temp_m5_24_26_r,temp_m5_24_26_i,`W9_real,`W9_imag,`W7_real,`W7_imag,`W16_real,`W16_imag);
butterfly butterfly1146 (clk,temp_m5_8_10_r,temp_m5_8_10_i,temp_m5_8_26_r,temp_m5_8_26_i,temp_m5_24_10_r,temp_m5_24_10_i,temp_m5_24_26_r,temp_m5_24_26_i,temp_b5_8_10_r,temp_b5_8_10_i,temp_b5_8_26_r,temp_b5_8_26_i,temp_b5_24_10_r,temp_b5_24_10_i,temp_b5_24_26_r,temp_b5_24_26_i);
MULT MULT1147 (clk,temp_b4_8_11_r,temp_b4_8_11_i,temp_b4_8_27_r,temp_b4_8_27_i,temp_b4_24_11_r,temp_b4_24_11_i,temp_b4_24_27_r,temp_b4_24_27_i,temp_m5_8_11_r,temp_m5_8_11_i,temp_m5_8_27_r,temp_m5_8_27_i,temp_m5_24_11_r,temp_m5_24_11_i,temp_m5_24_27_r,temp_m5_24_27_i,`W10_real,`W10_imag,`W7_real,`W7_imag,`W17_real,`W17_imag);
butterfly butterfly1147 (clk,temp_m5_8_11_r,temp_m5_8_11_i,temp_m5_8_27_r,temp_m5_8_27_i,temp_m5_24_11_r,temp_m5_24_11_i,temp_m5_24_27_r,temp_m5_24_27_i,temp_b5_8_11_r,temp_b5_8_11_i,temp_b5_8_27_r,temp_b5_8_27_i,temp_b5_24_11_r,temp_b5_24_11_i,temp_b5_24_27_r,temp_b5_24_27_i);
MULT MULT1148 (clk,temp_b4_8_12_r,temp_b4_8_12_i,temp_b4_8_28_r,temp_b4_8_28_i,temp_b4_24_12_r,temp_b4_24_12_i,temp_b4_24_28_r,temp_b4_24_28_i,temp_m5_8_12_r,temp_m5_8_12_i,temp_m5_8_28_r,temp_m5_8_28_i,temp_m5_24_12_r,temp_m5_24_12_i,temp_m5_24_28_r,temp_m5_24_28_i,`W11_real,`W11_imag,`W7_real,`W7_imag,`W18_real,`W18_imag);
butterfly butterfly1148 (clk,temp_m5_8_12_r,temp_m5_8_12_i,temp_m5_8_28_r,temp_m5_8_28_i,temp_m5_24_12_r,temp_m5_24_12_i,temp_m5_24_28_r,temp_m5_24_28_i,temp_b5_8_12_r,temp_b5_8_12_i,temp_b5_8_28_r,temp_b5_8_28_i,temp_b5_24_12_r,temp_b5_24_12_i,temp_b5_24_28_r,temp_b5_24_28_i);
MULT MULT1149 (clk,temp_b4_8_13_r,temp_b4_8_13_i,temp_b4_8_29_r,temp_b4_8_29_i,temp_b4_24_13_r,temp_b4_24_13_i,temp_b4_24_29_r,temp_b4_24_29_i,temp_m5_8_13_r,temp_m5_8_13_i,temp_m5_8_29_r,temp_m5_8_29_i,temp_m5_24_13_r,temp_m5_24_13_i,temp_m5_24_29_r,temp_m5_24_29_i,`W12_real,`W12_imag,`W7_real,`W7_imag,`W19_real,`W19_imag);
butterfly butterfly1149 (clk,temp_m5_8_13_r,temp_m5_8_13_i,temp_m5_8_29_r,temp_m5_8_29_i,temp_m5_24_13_r,temp_m5_24_13_i,temp_m5_24_29_r,temp_m5_24_29_i,temp_b5_8_13_r,temp_b5_8_13_i,temp_b5_8_29_r,temp_b5_8_29_i,temp_b5_24_13_r,temp_b5_24_13_i,temp_b5_24_29_r,temp_b5_24_29_i);
MULT MULT1150 (clk,temp_b4_8_14_r,temp_b4_8_14_i,temp_b4_8_30_r,temp_b4_8_30_i,temp_b4_24_14_r,temp_b4_24_14_i,temp_b4_24_30_r,temp_b4_24_30_i,temp_m5_8_14_r,temp_m5_8_14_i,temp_m5_8_30_r,temp_m5_8_30_i,temp_m5_24_14_r,temp_m5_24_14_i,temp_m5_24_30_r,temp_m5_24_30_i,`W13_real,`W13_imag,`W7_real,`W7_imag,`W20_real,`W20_imag);
butterfly butterfly1150 (clk,temp_m5_8_14_r,temp_m5_8_14_i,temp_m5_8_30_r,temp_m5_8_30_i,temp_m5_24_14_r,temp_m5_24_14_i,temp_m5_24_30_r,temp_m5_24_30_i,temp_b5_8_14_r,temp_b5_8_14_i,temp_b5_8_30_r,temp_b5_8_30_i,temp_b5_24_14_r,temp_b5_24_14_i,temp_b5_24_30_r,temp_b5_24_30_i);
MULT MULT1151 (clk,temp_b4_8_15_r,temp_b4_8_15_i,temp_b4_8_31_r,temp_b4_8_31_i,temp_b4_24_15_r,temp_b4_24_15_i,temp_b4_24_31_r,temp_b4_24_31_i,temp_m5_8_15_r,temp_m5_8_15_i,temp_m5_8_31_r,temp_m5_8_31_i,temp_m5_24_15_r,temp_m5_24_15_i,temp_m5_24_31_r,temp_m5_24_31_i,`W14_real,`W14_imag,`W7_real,`W7_imag,`W21_real,`W21_imag);
butterfly butterfly1151 (clk,temp_m5_8_15_r,temp_m5_8_15_i,temp_m5_8_31_r,temp_m5_8_31_i,temp_m5_24_15_r,temp_m5_24_15_i,temp_m5_24_31_r,temp_m5_24_31_i,temp_b5_8_15_r,temp_b5_8_15_i,temp_b5_8_31_r,temp_b5_8_31_i,temp_b5_24_15_r,temp_b5_24_15_i,temp_b5_24_31_r,temp_b5_24_31_i);
MULT MULT1152 (clk,temp_b4_8_16_r,temp_b4_8_16_i,temp_b4_8_32_r,temp_b4_8_32_i,temp_b4_24_16_r,temp_b4_24_16_i,temp_b4_24_32_r,temp_b4_24_32_i,temp_m5_8_16_r,temp_m5_8_16_i,temp_m5_8_32_r,temp_m5_8_32_i,temp_m5_24_16_r,temp_m5_24_16_i,temp_m5_24_32_r,temp_m5_24_32_i,`W15_real,`W15_imag,`W7_real,`W7_imag,`W22_real,`W22_imag);
butterfly butterfly1152 (clk,temp_m5_8_16_r,temp_m5_8_16_i,temp_m5_8_32_r,temp_m5_8_32_i,temp_m5_24_16_r,temp_m5_24_16_i,temp_m5_24_32_r,temp_m5_24_32_i,temp_b5_8_16_r,temp_b5_8_16_i,temp_b5_8_32_r,temp_b5_8_32_i,temp_b5_24_16_r,temp_b5_24_16_i,temp_b5_24_32_r,temp_b5_24_32_i);
MULT MULT1153 (clk,temp_b4_9_1_r,temp_b4_9_1_i,temp_b4_9_17_r,temp_b4_9_17_i,temp_b4_25_1_r,temp_b4_25_1_i,temp_b4_25_17_r,temp_b4_25_17_i,temp_m5_9_1_r,temp_m5_9_1_i,temp_m5_9_17_r,temp_m5_9_17_i,temp_m5_25_1_r,temp_m5_25_1_i,temp_m5_25_17_r,temp_m5_25_17_i,`W0_real,`W0_imag,`W8_real,`W8_imag,`W8_real,`W8_imag);
butterfly butterfly1153 (clk,temp_m5_9_1_r,temp_m5_9_1_i,temp_m5_9_17_r,temp_m5_9_17_i,temp_m5_25_1_r,temp_m5_25_1_i,temp_m5_25_17_r,temp_m5_25_17_i,temp_b5_9_1_r,temp_b5_9_1_i,temp_b5_9_17_r,temp_b5_9_17_i,temp_b5_25_1_r,temp_b5_25_1_i,temp_b5_25_17_r,temp_b5_25_17_i);
MULT MULT1154 (clk,temp_b4_9_2_r,temp_b4_9_2_i,temp_b4_9_18_r,temp_b4_9_18_i,temp_b4_25_2_r,temp_b4_25_2_i,temp_b4_25_18_r,temp_b4_25_18_i,temp_m5_9_2_r,temp_m5_9_2_i,temp_m5_9_18_r,temp_m5_9_18_i,temp_m5_25_2_r,temp_m5_25_2_i,temp_m5_25_18_r,temp_m5_25_18_i,`W1_real,`W1_imag,`W8_real,`W8_imag,`W9_real,`W9_imag);
butterfly butterfly1154 (clk,temp_m5_9_2_r,temp_m5_9_2_i,temp_m5_9_18_r,temp_m5_9_18_i,temp_m5_25_2_r,temp_m5_25_2_i,temp_m5_25_18_r,temp_m5_25_18_i,temp_b5_9_2_r,temp_b5_9_2_i,temp_b5_9_18_r,temp_b5_9_18_i,temp_b5_25_2_r,temp_b5_25_2_i,temp_b5_25_18_r,temp_b5_25_18_i);
MULT MULT1155 (clk,temp_b4_9_3_r,temp_b4_9_3_i,temp_b4_9_19_r,temp_b4_9_19_i,temp_b4_25_3_r,temp_b4_25_3_i,temp_b4_25_19_r,temp_b4_25_19_i,temp_m5_9_3_r,temp_m5_9_3_i,temp_m5_9_19_r,temp_m5_9_19_i,temp_m5_25_3_r,temp_m5_25_3_i,temp_m5_25_19_r,temp_m5_25_19_i,`W2_real,`W2_imag,`W8_real,`W8_imag,`W10_real,`W10_imag);
butterfly butterfly1155 (clk,temp_m5_9_3_r,temp_m5_9_3_i,temp_m5_9_19_r,temp_m5_9_19_i,temp_m5_25_3_r,temp_m5_25_3_i,temp_m5_25_19_r,temp_m5_25_19_i,temp_b5_9_3_r,temp_b5_9_3_i,temp_b5_9_19_r,temp_b5_9_19_i,temp_b5_25_3_r,temp_b5_25_3_i,temp_b5_25_19_r,temp_b5_25_19_i);
MULT MULT1156 (clk,temp_b4_9_4_r,temp_b4_9_4_i,temp_b4_9_20_r,temp_b4_9_20_i,temp_b4_25_4_r,temp_b4_25_4_i,temp_b4_25_20_r,temp_b4_25_20_i,temp_m5_9_4_r,temp_m5_9_4_i,temp_m5_9_20_r,temp_m5_9_20_i,temp_m5_25_4_r,temp_m5_25_4_i,temp_m5_25_20_r,temp_m5_25_20_i,`W3_real,`W3_imag,`W8_real,`W8_imag,`W11_real,`W11_imag);
butterfly butterfly1156 (clk,temp_m5_9_4_r,temp_m5_9_4_i,temp_m5_9_20_r,temp_m5_9_20_i,temp_m5_25_4_r,temp_m5_25_4_i,temp_m5_25_20_r,temp_m5_25_20_i,temp_b5_9_4_r,temp_b5_9_4_i,temp_b5_9_20_r,temp_b5_9_20_i,temp_b5_25_4_r,temp_b5_25_4_i,temp_b5_25_20_r,temp_b5_25_20_i);
MULT MULT1157 (clk,temp_b4_9_5_r,temp_b4_9_5_i,temp_b4_9_21_r,temp_b4_9_21_i,temp_b4_25_5_r,temp_b4_25_5_i,temp_b4_25_21_r,temp_b4_25_21_i,temp_m5_9_5_r,temp_m5_9_5_i,temp_m5_9_21_r,temp_m5_9_21_i,temp_m5_25_5_r,temp_m5_25_5_i,temp_m5_25_21_r,temp_m5_25_21_i,`W4_real,`W4_imag,`W8_real,`W8_imag,`W12_real,`W12_imag);
butterfly butterfly1157 (clk,temp_m5_9_5_r,temp_m5_9_5_i,temp_m5_9_21_r,temp_m5_9_21_i,temp_m5_25_5_r,temp_m5_25_5_i,temp_m5_25_21_r,temp_m5_25_21_i,temp_b5_9_5_r,temp_b5_9_5_i,temp_b5_9_21_r,temp_b5_9_21_i,temp_b5_25_5_r,temp_b5_25_5_i,temp_b5_25_21_r,temp_b5_25_21_i);
MULT MULT1158 (clk,temp_b4_9_6_r,temp_b4_9_6_i,temp_b4_9_22_r,temp_b4_9_22_i,temp_b4_25_6_r,temp_b4_25_6_i,temp_b4_25_22_r,temp_b4_25_22_i,temp_m5_9_6_r,temp_m5_9_6_i,temp_m5_9_22_r,temp_m5_9_22_i,temp_m5_25_6_r,temp_m5_25_6_i,temp_m5_25_22_r,temp_m5_25_22_i,`W5_real,`W5_imag,`W8_real,`W8_imag,`W13_real,`W13_imag);
butterfly butterfly1158 (clk,temp_m5_9_6_r,temp_m5_9_6_i,temp_m5_9_22_r,temp_m5_9_22_i,temp_m5_25_6_r,temp_m5_25_6_i,temp_m5_25_22_r,temp_m5_25_22_i,temp_b5_9_6_r,temp_b5_9_6_i,temp_b5_9_22_r,temp_b5_9_22_i,temp_b5_25_6_r,temp_b5_25_6_i,temp_b5_25_22_r,temp_b5_25_22_i);
MULT MULT1159 (clk,temp_b4_9_7_r,temp_b4_9_7_i,temp_b4_9_23_r,temp_b4_9_23_i,temp_b4_25_7_r,temp_b4_25_7_i,temp_b4_25_23_r,temp_b4_25_23_i,temp_m5_9_7_r,temp_m5_9_7_i,temp_m5_9_23_r,temp_m5_9_23_i,temp_m5_25_7_r,temp_m5_25_7_i,temp_m5_25_23_r,temp_m5_25_23_i,`W6_real,`W6_imag,`W8_real,`W8_imag,`W14_real,`W14_imag);
butterfly butterfly1159 (clk,temp_m5_9_7_r,temp_m5_9_7_i,temp_m5_9_23_r,temp_m5_9_23_i,temp_m5_25_7_r,temp_m5_25_7_i,temp_m5_25_23_r,temp_m5_25_23_i,temp_b5_9_7_r,temp_b5_9_7_i,temp_b5_9_23_r,temp_b5_9_23_i,temp_b5_25_7_r,temp_b5_25_7_i,temp_b5_25_23_r,temp_b5_25_23_i);
MULT MULT1160 (clk,temp_b4_9_8_r,temp_b4_9_8_i,temp_b4_9_24_r,temp_b4_9_24_i,temp_b4_25_8_r,temp_b4_25_8_i,temp_b4_25_24_r,temp_b4_25_24_i,temp_m5_9_8_r,temp_m5_9_8_i,temp_m5_9_24_r,temp_m5_9_24_i,temp_m5_25_8_r,temp_m5_25_8_i,temp_m5_25_24_r,temp_m5_25_24_i,`W7_real,`W7_imag,`W8_real,`W8_imag,`W15_real,`W15_imag);
butterfly butterfly1160 (clk,temp_m5_9_8_r,temp_m5_9_8_i,temp_m5_9_24_r,temp_m5_9_24_i,temp_m5_25_8_r,temp_m5_25_8_i,temp_m5_25_24_r,temp_m5_25_24_i,temp_b5_9_8_r,temp_b5_9_8_i,temp_b5_9_24_r,temp_b5_9_24_i,temp_b5_25_8_r,temp_b5_25_8_i,temp_b5_25_24_r,temp_b5_25_24_i);
MULT MULT1161 (clk,temp_b4_9_9_r,temp_b4_9_9_i,temp_b4_9_25_r,temp_b4_9_25_i,temp_b4_25_9_r,temp_b4_25_9_i,temp_b4_25_25_r,temp_b4_25_25_i,temp_m5_9_9_r,temp_m5_9_9_i,temp_m5_9_25_r,temp_m5_9_25_i,temp_m5_25_9_r,temp_m5_25_9_i,temp_m5_25_25_r,temp_m5_25_25_i,`W8_real,`W8_imag,`W8_real,`W8_imag,`W16_real,`W16_imag);
butterfly butterfly1161 (clk,temp_m5_9_9_r,temp_m5_9_9_i,temp_m5_9_25_r,temp_m5_9_25_i,temp_m5_25_9_r,temp_m5_25_9_i,temp_m5_25_25_r,temp_m5_25_25_i,temp_b5_9_9_r,temp_b5_9_9_i,temp_b5_9_25_r,temp_b5_9_25_i,temp_b5_25_9_r,temp_b5_25_9_i,temp_b5_25_25_r,temp_b5_25_25_i);
MULT MULT1162 (clk,temp_b4_9_10_r,temp_b4_9_10_i,temp_b4_9_26_r,temp_b4_9_26_i,temp_b4_25_10_r,temp_b4_25_10_i,temp_b4_25_26_r,temp_b4_25_26_i,temp_m5_9_10_r,temp_m5_9_10_i,temp_m5_9_26_r,temp_m5_9_26_i,temp_m5_25_10_r,temp_m5_25_10_i,temp_m5_25_26_r,temp_m5_25_26_i,`W9_real,`W9_imag,`W8_real,`W8_imag,`W17_real,`W17_imag);
butterfly butterfly1162 (clk,temp_m5_9_10_r,temp_m5_9_10_i,temp_m5_9_26_r,temp_m5_9_26_i,temp_m5_25_10_r,temp_m5_25_10_i,temp_m5_25_26_r,temp_m5_25_26_i,temp_b5_9_10_r,temp_b5_9_10_i,temp_b5_9_26_r,temp_b5_9_26_i,temp_b5_25_10_r,temp_b5_25_10_i,temp_b5_25_26_r,temp_b5_25_26_i);
MULT MULT1163 (clk,temp_b4_9_11_r,temp_b4_9_11_i,temp_b4_9_27_r,temp_b4_9_27_i,temp_b4_25_11_r,temp_b4_25_11_i,temp_b4_25_27_r,temp_b4_25_27_i,temp_m5_9_11_r,temp_m5_9_11_i,temp_m5_9_27_r,temp_m5_9_27_i,temp_m5_25_11_r,temp_m5_25_11_i,temp_m5_25_27_r,temp_m5_25_27_i,`W10_real,`W10_imag,`W8_real,`W8_imag,`W18_real,`W18_imag);
butterfly butterfly1163 (clk,temp_m5_9_11_r,temp_m5_9_11_i,temp_m5_9_27_r,temp_m5_9_27_i,temp_m5_25_11_r,temp_m5_25_11_i,temp_m5_25_27_r,temp_m5_25_27_i,temp_b5_9_11_r,temp_b5_9_11_i,temp_b5_9_27_r,temp_b5_9_27_i,temp_b5_25_11_r,temp_b5_25_11_i,temp_b5_25_27_r,temp_b5_25_27_i);
MULT MULT1164 (clk,temp_b4_9_12_r,temp_b4_9_12_i,temp_b4_9_28_r,temp_b4_9_28_i,temp_b4_25_12_r,temp_b4_25_12_i,temp_b4_25_28_r,temp_b4_25_28_i,temp_m5_9_12_r,temp_m5_9_12_i,temp_m5_9_28_r,temp_m5_9_28_i,temp_m5_25_12_r,temp_m5_25_12_i,temp_m5_25_28_r,temp_m5_25_28_i,`W11_real,`W11_imag,`W8_real,`W8_imag,`W19_real,`W19_imag);
butterfly butterfly1164 (clk,temp_m5_9_12_r,temp_m5_9_12_i,temp_m5_9_28_r,temp_m5_9_28_i,temp_m5_25_12_r,temp_m5_25_12_i,temp_m5_25_28_r,temp_m5_25_28_i,temp_b5_9_12_r,temp_b5_9_12_i,temp_b5_9_28_r,temp_b5_9_28_i,temp_b5_25_12_r,temp_b5_25_12_i,temp_b5_25_28_r,temp_b5_25_28_i);
MULT MULT1165 (clk,temp_b4_9_13_r,temp_b4_9_13_i,temp_b4_9_29_r,temp_b4_9_29_i,temp_b4_25_13_r,temp_b4_25_13_i,temp_b4_25_29_r,temp_b4_25_29_i,temp_m5_9_13_r,temp_m5_9_13_i,temp_m5_9_29_r,temp_m5_9_29_i,temp_m5_25_13_r,temp_m5_25_13_i,temp_m5_25_29_r,temp_m5_25_29_i,`W12_real,`W12_imag,`W8_real,`W8_imag,`W20_real,`W20_imag);
butterfly butterfly1165 (clk,temp_m5_9_13_r,temp_m5_9_13_i,temp_m5_9_29_r,temp_m5_9_29_i,temp_m5_25_13_r,temp_m5_25_13_i,temp_m5_25_29_r,temp_m5_25_29_i,temp_b5_9_13_r,temp_b5_9_13_i,temp_b5_9_29_r,temp_b5_9_29_i,temp_b5_25_13_r,temp_b5_25_13_i,temp_b5_25_29_r,temp_b5_25_29_i);
MULT MULT1166 (clk,temp_b4_9_14_r,temp_b4_9_14_i,temp_b4_9_30_r,temp_b4_9_30_i,temp_b4_25_14_r,temp_b4_25_14_i,temp_b4_25_30_r,temp_b4_25_30_i,temp_m5_9_14_r,temp_m5_9_14_i,temp_m5_9_30_r,temp_m5_9_30_i,temp_m5_25_14_r,temp_m5_25_14_i,temp_m5_25_30_r,temp_m5_25_30_i,`W13_real,`W13_imag,`W8_real,`W8_imag,`W21_real,`W21_imag);
butterfly butterfly1166 (clk,temp_m5_9_14_r,temp_m5_9_14_i,temp_m5_9_30_r,temp_m5_9_30_i,temp_m5_25_14_r,temp_m5_25_14_i,temp_m5_25_30_r,temp_m5_25_30_i,temp_b5_9_14_r,temp_b5_9_14_i,temp_b5_9_30_r,temp_b5_9_30_i,temp_b5_25_14_r,temp_b5_25_14_i,temp_b5_25_30_r,temp_b5_25_30_i);
MULT MULT1167 (clk,temp_b4_9_15_r,temp_b4_9_15_i,temp_b4_9_31_r,temp_b4_9_31_i,temp_b4_25_15_r,temp_b4_25_15_i,temp_b4_25_31_r,temp_b4_25_31_i,temp_m5_9_15_r,temp_m5_9_15_i,temp_m5_9_31_r,temp_m5_9_31_i,temp_m5_25_15_r,temp_m5_25_15_i,temp_m5_25_31_r,temp_m5_25_31_i,`W14_real,`W14_imag,`W8_real,`W8_imag,`W22_real,`W22_imag);
butterfly butterfly1167 (clk,temp_m5_9_15_r,temp_m5_9_15_i,temp_m5_9_31_r,temp_m5_9_31_i,temp_m5_25_15_r,temp_m5_25_15_i,temp_m5_25_31_r,temp_m5_25_31_i,temp_b5_9_15_r,temp_b5_9_15_i,temp_b5_9_31_r,temp_b5_9_31_i,temp_b5_25_15_r,temp_b5_25_15_i,temp_b5_25_31_r,temp_b5_25_31_i);
MULT MULT1168 (clk,temp_b4_9_16_r,temp_b4_9_16_i,temp_b4_9_32_r,temp_b4_9_32_i,temp_b4_25_16_r,temp_b4_25_16_i,temp_b4_25_32_r,temp_b4_25_32_i,temp_m5_9_16_r,temp_m5_9_16_i,temp_m5_9_32_r,temp_m5_9_32_i,temp_m5_25_16_r,temp_m5_25_16_i,temp_m5_25_32_r,temp_m5_25_32_i,`W15_real,`W15_imag,`W8_real,`W8_imag,`W23_real,`W23_imag);
butterfly butterfly1168 (clk,temp_m5_9_16_r,temp_m5_9_16_i,temp_m5_9_32_r,temp_m5_9_32_i,temp_m5_25_16_r,temp_m5_25_16_i,temp_m5_25_32_r,temp_m5_25_32_i,temp_b5_9_16_r,temp_b5_9_16_i,temp_b5_9_32_r,temp_b5_9_32_i,temp_b5_25_16_r,temp_b5_25_16_i,temp_b5_25_32_r,temp_b5_25_32_i);
MULT MULT1169 (clk,temp_b4_10_1_r,temp_b4_10_1_i,temp_b4_10_17_r,temp_b4_10_17_i,temp_b4_26_1_r,temp_b4_26_1_i,temp_b4_26_17_r,temp_b4_26_17_i,temp_m5_10_1_r,temp_m5_10_1_i,temp_m5_10_17_r,temp_m5_10_17_i,temp_m5_26_1_r,temp_m5_26_1_i,temp_m5_26_17_r,temp_m5_26_17_i,`W0_real,`W0_imag,`W9_real,`W9_imag,`W9_real,`W9_imag);
butterfly butterfly1169 (clk,temp_m5_10_1_r,temp_m5_10_1_i,temp_m5_10_17_r,temp_m5_10_17_i,temp_m5_26_1_r,temp_m5_26_1_i,temp_m5_26_17_r,temp_m5_26_17_i,temp_b5_10_1_r,temp_b5_10_1_i,temp_b5_10_17_r,temp_b5_10_17_i,temp_b5_26_1_r,temp_b5_26_1_i,temp_b5_26_17_r,temp_b5_26_17_i);
MULT MULT1170 (clk,temp_b4_10_2_r,temp_b4_10_2_i,temp_b4_10_18_r,temp_b4_10_18_i,temp_b4_26_2_r,temp_b4_26_2_i,temp_b4_26_18_r,temp_b4_26_18_i,temp_m5_10_2_r,temp_m5_10_2_i,temp_m5_10_18_r,temp_m5_10_18_i,temp_m5_26_2_r,temp_m5_26_2_i,temp_m5_26_18_r,temp_m5_26_18_i,`W1_real,`W1_imag,`W9_real,`W9_imag,`W10_real,`W10_imag);
butterfly butterfly1170 (clk,temp_m5_10_2_r,temp_m5_10_2_i,temp_m5_10_18_r,temp_m5_10_18_i,temp_m5_26_2_r,temp_m5_26_2_i,temp_m5_26_18_r,temp_m5_26_18_i,temp_b5_10_2_r,temp_b5_10_2_i,temp_b5_10_18_r,temp_b5_10_18_i,temp_b5_26_2_r,temp_b5_26_2_i,temp_b5_26_18_r,temp_b5_26_18_i);
MULT MULT1171 (clk,temp_b4_10_3_r,temp_b4_10_3_i,temp_b4_10_19_r,temp_b4_10_19_i,temp_b4_26_3_r,temp_b4_26_3_i,temp_b4_26_19_r,temp_b4_26_19_i,temp_m5_10_3_r,temp_m5_10_3_i,temp_m5_10_19_r,temp_m5_10_19_i,temp_m5_26_3_r,temp_m5_26_3_i,temp_m5_26_19_r,temp_m5_26_19_i,`W2_real,`W2_imag,`W9_real,`W9_imag,`W11_real,`W11_imag);
butterfly butterfly1171 (clk,temp_m5_10_3_r,temp_m5_10_3_i,temp_m5_10_19_r,temp_m5_10_19_i,temp_m5_26_3_r,temp_m5_26_3_i,temp_m5_26_19_r,temp_m5_26_19_i,temp_b5_10_3_r,temp_b5_10_3_i,temp_b5_10_19_r,temp_b5_10_19_i,temp_b5_26_3_r,temp_b5_26_3_i,temp_b5_26_19_r,temp_b5_26_19_i);
MULT MULT1172 (clk,temp_b4_10_4_r,temp_b4_10_4_i,temp_b4_10_20_r,temp_b4_10_20_i,temp_b4_26_4_r,temp_b4_26_4_i,temp_b4_26_20_r,temp_b4_26_20_i,temp_m5_10_4_r,temp_m5_10_4_i,temp_m5_10_20_r,temp_m5_10_20_i,temp_m5_26_4_r,temp_m5_26_4_i,temp_m5_26_20_r,temp_m5_26_20_i,`W3_real,`W3_imag,`W9_real,`W9_imag,`W12_real,`W12_imag);
butterfly butterfly1172 (clk,temp_m5_10_4_r,temp_m5_10_4_i,temp_m5_10_20_r,temp_m5_10_20_i,temp_m5_26_4_r,temp_m5_26_4_i,temp_m5_26_20_r,temp_m5_26_20_i,temp_b5_10_4_r,temp_b5_10_4_i,temp_b5_10_20_r,temp_b5_10_20_i,temp_b5_26_4_r,temp_b5_26_4_i,temp_b5_26_20_r,temp_b5_26_20_i);
MULT MULT1173 (clk,temp_b4_10_5_r,temp_b4_10_5_i,temp_b4_10_21_r,temp_b4_10_21_i,temp_b4_26_5_r,temp_b4_26_5_i,temp_b4_26_21_r,temp_b4_26_21_i,temp_m5_10_5_r,temp_m5_10_5_i,temp_m5_10_21_r,temp_m5_10_21_i,temp_m5_26_5_r,temp_m5_26_5_i,temp_m5_26_21_r,temp_m5_26_21_i,`W4_real,`W4_imag,`W9_real,`W9_imag,`W13_real,`W13_imag);
butterfly butterfly1173 (clk,temp_m5_10_5_r,temp_m5_10_5_i,temp_m5_10_21_r,temp_m5_10_21_i,temp_m5_26_5_r,temp_m5_26_5_i,temp_m5_26_21_r,temp_m5_26_21_i,temp_b5_10_5_r,temp_b5_10_5_i,temp_b5_10_21_r,temp_b5_10_21_i,temp_b5_26_5_r,temp_b5_26_5_i,temp_b5_26_21_r,temp_b5_26_21_i);
MULT MULT1174 (clk,temp_b4_10_6_r,temp_b4_10_6_i,temp_b4_10_22_r,temp_b4_10_22_i,temp_b4_26_6_r,temp_b4_26_6_i,temp_b4_26_22_r,temp_b4_26_22_i,temp_m5_10_6_r,temp_m5_10_6_i,temp_m5_10_22_r,temp_m5_10_22_i,temp_m5_26_6_r,temp_m5_26_6_i,temp_m5_26_22_r,temp_m5_26_22_i,`W5_real,`W5_imag,`W9_real,`W9_imag,`W14_real,`W14_imag);
butterfly butterfly1174 (clk,temp_m5_10_6_r,temp_m5_10_6_i,temp_m5_10_22_r,temp_m5_10_22_i,temp_m5_26_6_r,temp_m5_26_6_i,temp_m5_26_22_r,temp_m5_26_22_i,temp_b5_10_6_r,temp_b5_10_6_i,temp_b5_10_22_r,temp_b5_10_22_i,temp_b5_26_6_r,temp_b5_26_6_i,temp_b5_26_22_r,temp_b5_26_22_i);
MULT MULT1175 (clk,temp_b4_10_7_r,temp_b4_10_7_i,temp_b4_10_23_r,temp_b4_10_23_i,temp_b4_26_7_r,temp_b4_26_7_i,temp_b4_26_23_r,temp_b4_26_23_i,temp_m5_10_7_r,temp_m5_10_7_i,temp_m5_10_23_r,temp_m5_10_23_i,temp_m5_26_7_r,temp_m5_26_7_i,temp_m5_26_23_r,temp_m5_26_23_i,`W6_real,`W6_imag,`W9_real,`W9_imag,`W15_real,`W15_imag);
butterfly butterfly1175 (clk,temp_m5_10_7_r,temp_m5_10_7_i,temp_m5_10_23_r,temp_m5_10_23_i,temp_m5_26_7_r,temp_m5_26_7_i,temp_m5_26_23_r,temp_m5_26_23_i,temp_b5_10_7_r,temp_b5_10_7_i,temp_b5_10_23_r,temp_b5_10_23_i,temp_b5_26_7_r,temp_b5_26_7_i,temp_b5_26_23_r,temp_b5_26_23_i);
MULT MULT1176 (clk,temp_b4_10_8_r,temp_b4_10_8_i,temp_b4_10_24_r,temp_b4_10_24_i,temp_b4_26_8_r,temp_b4_26_8_i,temp_b4_26_24_r,temp_b4_26_24_i,temp_m5_10_8_r,temp_m5_10_8_i,temp_m5_10_24_r,temp_m5_10_24_i,temp_m5_26_8_r,temp_m5_26_8_i,temp_m5_26_24_r,temp_m5_26_24_i,`W7_real,`W7_imag,`W9_real,`W9_imag,`W16_real,`W16_imag);
butterfly butterfly1176 (clk,temp_m5_10_8_r,temp_m5_10_8_i,temp_m5_10_24_r,temp_m5_10_24_i,temp_m5_26_8_r,temp_m5_26_8_i,temp_m5_26_24_r,temp_m5_26_24_i,temp_b5_10_8_r,temp_b5_10_8_i,temp_b5_10_24_r,temp_b5_10_24_i,temp_b5_26_8_r,temp_b5_26_8_i,temp_b5_26_24_r,temp_b5_26_24_i);
MULT MULT1177 (clk,temp_b4_10_9_r,temp_b4_10_9_i,temp_b4_10_25_r,temp_b4_10_25_i,temp_b4_26_9_r,temp_b4_26_9_i,temp_b4_26_25_r,temp_b4_26_25_i,temp_m5_10_9_r,temp_m5_10_9_i,temp_m5_10_25_r,temp_m5_10_25_i,temp_m5_26_9_r,temp_m5_26_9_i,temp_m5_26_25_r,temp_m5_26_25_i,`W8_real,`W8_imag,`W9_real,`W9_imag,`W17_real,`W17_imag);
butterfly butterfly1177 (clk,temp_m5_10_9_r,temp_m5_10_9_i,temp_m5_10_25_r,temp_m5_10_25_i,temp_m5_26_9_r,temp_m5_26_9_i,temp_m5_26_25_r,temp_m5_26_25_i,temp_b5_10_9_r,temp_b5_10_9_i,temp_b5_10_25_r,temp_b5_10_25_i,temp_b5_26_9_r,temp_b5_26_9_i,temp_b5_26_25_r,temp_b5_26_25_i);
MULT MULT1178 (clk,temp_b4_10_10_r,temp_b4_10_10_i,temp_b4_10_26_r,temp_b4_10_26_i,temp_b4_26_10_r,temp_b4_26_10_i,temp_b4_26_26_r,temp_b4_26_26_i,temp_m5_10_10_r,temp_m5_10_10_i,temp_m5_10_26_r,temp_m5_10_26_i,temp_m5_26_10_r,temp_m5_26_10_i,temp_m5_26_26_r,temp_m5_26_26_i,`W9_real,`W9_imag,`W9_real,`W9_imag,`W18_real,`W18_imag);
butterfly butterfly1178 (clk,temp_m5_10_10_r,temp_m5_10_10_i,temp_m5_10_26_r,temp_m5_10_26_i,temp_m5_26_10_r,temp_m5_26_10_i,temp_m5_26_26_r,temp_m5_26_26_i,temp_b5_10_10_r,temp_b5_10_10_i,temp_b5_10_26_r,temp_b5_10_26_i,temp_b5_26_10_r,temp_b5_26_10_i,temp_b5_26_26_r,temp_b5_26_26_i);
MULT MULT1179 (clk,temp_b4_10_11_r,temp_b4_10_11_i,temp_b4_10_27_r,temp_b4_10_27_i,temp_b4_26_11_r,temp_b4_26_11_i,temp_b4_26_27_r,temp_b4_26_27_i,temp_m5_10_11_r,temp_m5_10_11_i,temp_m5_10_27_r,temp_m5_10_27_i,temp_m5_26_11_r,temp_m5_26_11_i,temp_m5_26_27_r,temp_m5_26_27_i,`W10_real,`W10_imag,`W9_real,`W9_imag,`W19_real,`W19_imag);
butterfly butterfly1179 (clk,temp_m5_10_11_r,temp_m5_10_11_i,temp_m5_10_27_r,temp_m5_10_27_i,temp_m5_26_11_r,temp_m5_26_11_i,temp_m5_26_27_r,temp_m5_26_27_i,temp_b5_10_11_r,temp_b5_10_11_i,temp_b5_10_27_r,temp_b5_10_27_i,temp_b5_26_11_r,temp_b5_26_11_i,temp_b5_26_27_r,temp_b5_26_27_i);
MULT MULT1180 (clk,temp_b4_10_12_r,temp_b4_10_12_i,temp_b4_10_28_r,temp_b4_10_28_i,temp_b4_26_12_r,temp_b4_26_12_i,temp_b4_26_28_r,temp_b4_26_28_i,temp_m5_10_12_r,temp_m5_10_12_i,temp_m5_10_28_r,temp_m5_10_28_i,temp_m5_26_12_r,temp_m5_26_12_i,temp_m5_26_28_r,temp_m5_26_28_i,`W11_real,`W11_imag,`W9_real,`W9_imag,`W20_real,`W20_imag);
butterfly butterfly1180 (clk,temp_m5_10_12_r,temp_m5_10_12_i,temp_m5_10_28_r,temp_m5_10_28_i,temp_m5_26_12_r,temp_m5_26_12_i,temp_m5_26_28_r,temp_m5_26_28_i,temp_b5_10_12_r,temp_b5_10_12_i,temp_b5_10_28_r,temp_b5_10_28_i,temp_b5_26_12_r,temp_b5_26_12_i,temp_b5_26_28_r,temp_b5_26_28_i);
MULT MULT1181 (clk,temp_b4_10_13_r,temp_b4_10_13_i,temp_b4_10_29_r,temp_b4_10_29_i,temp_b4_26_13_r,temp_b4_26_13_i,temp_b4_26_29_r,temp_b4_26_29_i,temp_m5_10_13_r,temp_m5_10_13_i,temp_m5_10_29_r,temp_m5_10_29_i,temp_m5_26_13_r,temp_m5_26_13_i,temp_m5_26_29_r,temp_m5_26_29_i,`W12_real,`W12_imag,`W9_real,`W9_imag,`W21_real,`W21_imag);
butterfly butterfly1181 (clk,temp_m5_10_13_r,temp_m5_10_13_i,temp_m5_10_29_r,temp_m5_10_29_i,temp_m5_26_13_r,temp_m5_26_13_i,temp_m5_26_29_r,temp_m5_26_29_i,temp_b5_10_13_r,temp_b5_10_13_i,temp_b5_10_29_r,temp_b5_10_29_i,temp_b5_26_13_r,temp_b5_26_13_i,temp_b5_26_29_r,temp_b5_26_29_i);
MULT MULT1182 (clk,temp_b4_10_14_r,temp_b4_10_14_i,temp_b4_10_30_r,temp_b4_10_30_i,temp_b4_26_14_r,temp_b4_26_14_i,temp_b4_26_30_r,temp_b4_26_30_i,temp_m5_10_14_r,temp_m5_10_14_i,temp_m5_10_30_r,temp_m5_10_30_i,temp_m5_26_14_r,temp_m5_26_14_i,temp_m5_26_30_r,temp_m5_26_30_i,`W13_real,`W13_imag,`W9_real,`W9_imag,`W22_real,`W22_imag);
butterfly butterfly1182 (clk,temp_m5_10_14_r,temp_m5_10_14_i,temp_m5_10_30_r,temp_m5_10_30_i,temp_m5_26_14_r,temp_m5_26_14_i,temp_m5_26_30_r,temp_m5_26_30_i,temp_b5_10_14_r,temp_b5_10_14_i,temp_b5_10_30_r,temp_b5_10_30_i,temp_b5_26_14_r,temp_b5_26_14_i,temp_b5_26_30_r,temp_b5_26_30_i);
MULT MULT1183 (clk,temp_b4_10_15_r,temp_b4_10_15_i,temp_b4_10_31_r,temp_b4_10_31_i,temp_b4_26_15_r,temp_b4_26_15_i,temp_b4_26_31_r,temp_b4_26_31_i,temp_m5_10_15_r,temp_m5_10_15_i,temp_m5_10_31_r,temp_m5_10_31_i,temp_m5_26_15_r,temp_m5_26_15_i,temp_m5_26_31_r,temp_m5_26_31_i,`W14_real,`W14_imag,`W9_real,`W9_imag,`W23_real,`W23_imag);
butterfly butterfly1183 (clk,temp_m5_10_15_r,temp_m5_10_15_i,temp_m5_10_31_r,temp_m5_10_31_i,temp_m5_26_15_r,temp_m5_26_15_i,temp_m5_26_31_r,temp_m5_26_31_i,temp_b5_10_15_r,temp_b5_10_15_i,temp_b5_10_31_r,temp_b5_10_31_i,temp_b5_26_15_r,temp_b5_26_15_i,temp_b5_26_31_r,temp_b5_26_31_i);
MULT MULT1184 (clk,temp_b4_10_16_r,temp_b4_10_16_i,temp_b4_10_32_r,temp_b4_10_32_i,temp_b4_26_16_r,temp_b4_26_16_i,temp_b4_26_32_r,temp_b4_26_32_i,temp_m5_10_16_r,temp_m5_10_16_i,temp_m5_10_32_r,temp_m5_10_32_i,temp_m5_26_16_r,temp_m5_26_16_i,temp_m5_26_32_r,temp_m5_26_32_i,`W15_real,`W15_imag,`W9_real,`W9_imag,`W24_real,`W24_imag);
butterfly butterfly1184 (clk,temp_m5_10_16_r,temp_m5_10_16_i,temp_m5_10_32_r,temp_m5_10_32_i,temp_m5_26_16_r,temp_m5_26_16_i,temp_m5_26_32_r,temp_m5_26_32_i,temp_b5_10_16_r,temp_b5_10_16_i,temp_b5_10_32_r,temp_b5_10_32_i,temp_b5_26_16_r,temp_b5_26_16_i,temp_b5_26_32_r,temp_b5_26_32_i);
MULT MULT1185 (clk,temp_b4_11_1_r,temp_b4_11_1_i,temp_b4_11_17_r,temp_b4_11_17_i,temp_b4_27_1_r,temp_b4_27_1_i,temp_b4_27_17_r,temp_b4_27_17_i,temp_m5_11_1_r,temp_m5_11_1_i,temp_m5_11_17_r,temp_m5_11_17_i,temp_m5_27_1_r,temp_m5_27_1_i,temp_m5_27_17_r,temp_m5_27_17_i,`W0_real,`W0_imag,`W10_real,`W10_imag,`W10_real,`W10_imag);
butterfly butterfly1185 (clk,temp_m5_11_1_r,temp_m5_11_1_i,temp_m5_11_17_r,temp_m5_11_17_i,temp_m5_27_1_r,temp_m5_27_1_i,temp_m5_27_17_r,temp_m5_27_17_i,temp_b5_11_1_r,temp_b5_11_1_i,temp_b5_11_17_r,temp_b5_11_17_i,temp_b5_27_1_r,temp_b5_27_1_i,temp_b5_27_17_r,temp_b5_27_17_i);
MULT MULT1186 (clk,temp_b4_11_2_r,temp_b4_11_2_i,temp_b4_11_18_r,temp_b4_11_18_i,temp_b4_27_2_r,temp_b4_27_2_i,temp_b4_27_18_r,temp_b4_27_18_i,temp_m5_11_2_r,temp_m5_11_2_i,temp_m5_11_18_r,temp_m5_11_18_i,temp_m5_27_2_r,temp_m5_27_2_i,temp_m5_27_18_r,temp_m5_27_18_i,`W1_real,`W1_imag,`W10_real,`W10_imag,`W11_real,`W11_imag);
butterfly butterfly1186 (clk,temp_m5_11_2_r,temp_m5_11_2_i,temp_m5_11_18_r,temp_m5_11_18_i,temp_m5_27_2_r,temp_m5_27_2_i,temp_m5_27_18_r,temp_m5_27_18_i,temp_b5_11_2_r,temp_b5_11_2_i,temp_b5_11_18_r,temp_b5_11_18_i,temp_b5_27_2_r,temp_b5_27_2_i,temp_b5_27_18_r,temp_b5_27_18_i);
MULT MULT1187 (clk,temp_b4_11_3_r,temp_b4_11_3_i,temp_b4_11_19_r,temp_b4_11_19_i,temp_b4_27_3_r,temp_b4_27_3_i,temp_b4_27_19_r,temp_b4_27_19_i,temp_m5_11_3_r,temp_m5_11_3_i,temp_m5_11_19_r,temp_m5_11_19_i,temp_m5_27_3_r,temp_m5_27_3_i,temp_m5_27_19_r,temp_m5_27_19_i,`W2_real,`W2_imag,`W10_real,`W10_imag,`W12_real,`W12_imag);
butterfly butterfly1187 (clk,temp_m5_11_3_r,temp_m5_11_3_i,temp_m5_11_19_r,temp_m5_11_19_i,temp_m5_27_3_r,temp_m5_27_3_i,temp_m5_27_19_r,temp_m5_27_19_i,temp_b5_11_3_r,temp_b5_11_3_i,temp_b5_11_19_r,temp_b5_11_19_i,temp_b5_27_3_r,temp_b5_27_3_i,temp_b5_27_19_r,temp_b5_27_19_i);
MULT MULT1188 (clk,temp_b4_11_4_r,temp_b4_11_4_i,temp_b4_11_20_r,temp_b4_11_20_i,temp_b4_27_4_r,temp_b4_27_4_i,temp_b4_27_20_r,temp_b4_27_20_i,temp_m5_11_4_r,temp_m5_11_4_i,temp_m5_11_20_r,temp_m5_11_20_i,temp_m5_27_4_r,temp_m5_27_4_i,temp_m5_27_20_r,temp_m5_27_20_i,`W3_real,`W3_imag,`W10_real,`W10_imag,`W13_real,`W13_imag);
butterfly butterfly1188 (clk,temp_m5_11_4_r,temp_m5_11_4_i,temp_m5_11_20_r,temp_m5_11_20_i,temp_m5_27_4_r,temp_m5_27_4_i,temp_m5_27_20_r,temp_m5_27_20_i,temp_b5_11_4_r,temp_b5_11_4_i,temp_b5_11_20_r,temp_b5_11_20_i,temp_b5_27_4_r,temp_b5_27_4_i,temp_b5_27_20_r,temp_b5_27_20_i);
MULT MULT1189 (clk,temp_b4_11_5_r,temp_b4_11_5_i,temp_b4_11_21_r,temp_b4_11_21_i,temp_b4_27_5_r,temp_b4_27_5_i,temp_b4_27_21_r,temp_b4_27_21_i,temp_m5_11_5_r,temp_m5_11_5_i,temp_m5_11_21_r,temp_m5_11_21_i,temp_m5_27_5_r,temp_m5_27_5_i,temp_m5_27_21_r,temp_m5_27_21_i,`W4_real,`W4_imag,`W10_real,`W10_imag,`W14_real,`W14_imag);
butterfly butterfly1189 (clk,temp_m5_11_5_r,temp_m5_11_5_i,temp_m5_11_21_r,temp_m5_11_21_i,temp_m5_27_5_r,temp_m5_27_5_i,temp_m5_27_21_r,temp_m5_27_21_i,temp_b5_11_5_r,temp_b5_11_5_i,temp_b5_11_21_r,temp_b5_11_21_i,temp_b5_27_5_r,temp_b5_27_5_i,temp_b5_27_21_r,temp_b5_27_21_i);
MULT MULT1190 (clk,temp_b4_11_6_r,temp_b4_11_6_i,temp_b4_11_22_r,temp_b4_11_22_i,temp_b4_27_6_r,temp_b4_27_6_i,temp_b4_27_22_r,temp_b4_27_22_i,temp_m5_11_6_r,temp_m5_11_6_i,temp_m5_11_22_r,temp_m5_11_22_i,temp_m5_27_6_r,temp_m5_27_6_i,temp_m5_27_22_r,temp_m5_27_22_i,`W5_real,`W5_imag,`W10_real,`W10_imag,`W15_real,`W15_imag);
butterfly butterfly1190 (clk,temp_m5_11_6_r,temp_m5_11_6_i,temp_m5_11_22_r,temp_m5_11_22_i,temp_m5_27_6_r,temp_m5_27_6_i,temp_m5_27_22_r,temp_m5_27_22_i,temp_b5_11_6_r,temp_b5_11_6_i,temp_b5_11_22_r,temp_b5_11_22_i,temp_b5_27_6_r,temp_b5_27_6_i,temp_b5_27_22_r,temp_b5_27_22_i);
MULT MULT1191 (clk,temp_b4_11_7_r,temp_b4_11_7_i,temp_b4_11_23_r,temp_b4_11_23_i,temp_b4_27_7_r,temp_b4_27_7_i,temp_b4_27_23_r,temp_b4_27_23_i,temp_m5_11_7_r,temp_m5_11_7_i,temp_m5_11_23_r,temp_m5_11_23_i,temp_m5_27_7_r,temp_m5_27_7_i,temp_m5_27_23_r,temp_m5_27_23_i,`W6_real,`W6_imag,`W10_real,`W10_imag,`W16_real,`W16_imag);
butterfly butterfly1191 (clk,temp_m5_11_7_r,temp_m5_11_7_i,temp_m5_11_23_r,temp_m5_11_23_i,temp_m5_27_7_r,temp_m5_27_7_i,temp_m5_27_23_r,temp_m5_27_23_i,temp_b5_11_7_r,temp_b5_11_7_i,temp_b5_11_23_r,temp_b5_11_23_i,temp_b5_27_7_r,temp_b5_27_7_i,temp_b5_27_23_r,temp_b5_27_23_i);
MULT MULT1192 (clk,temp_b4_11_8_r,temp_b4_11_8_i,temp_b4_11_24_r,temp_b4_11_24_i,temp_b4_27_8_r,temp_b4_27_8_i,temp_b4_27_24_r,temp_b4_27_24_i,temp_m5_11_8_r,temp_m5_11_8_i,temp_m5_11_24_r,temp_m5_11_24_i,temp_m5_27_8_r,temp_m5_27_8_i,temp_m5_27_24_r,temp_m5_27_24_i,`W7_real,`W7_imag,`W10_real,`W10_imag,`W17_real,`W17_imag);
butterfly butterfly1192 (clk,temp_m5_11_8_r,temp_m5_11_8_i,temp_m5_11_24_r,temp_m5_11_24_i,temp_m5_27_8_r,temp_m5_27_8_i,temp_m5_27_24_r,temp_m5_27_24_i,temp_b5_11_8_r,temp_b5_11_8_i,temp_b5_11_24_r,temp_b5_11_24_i,temp_b5_27_8_r,temp_b5_27_8_i,temp_b5_27_24_r,temp_b5_27_24_i);
MULT MULT1193 (clk,temp_b4_11_9_r,temp_b4_11_9_i,temp_b4_11_25_r,temp_b4_11_25_i,temp_b4_27_9_r,temp_b4_27_9_i,temp_b4_27_25_r,temp_b4_27_25_i,temp_m5_11_9_r,temp_m5_11_9_i,temp_m5_11_25_r,temp_m5_11_25_i,temp_m5_27_9_r,temp_m5_27_9_i,temp_m5_27_25_r,temp_m5_27_25_i,`W8_real,`W8_imag,`W10_real,`W10_imag,`W18_real,`W18_imag);
butterfly butterfly1193 (clk,temp_m5_11_9_r,temp_m5_11_9_i,temp_m5_11_25_r,temp_m5_11_25_i,temp_m5_27_9_r,temp_m5_27_9_i,temp_m5_27_25_r,temp_m5_27_25_i,temp_b5_11_9_r,temp_b5_11_9_i,temp_b5_11_25_r,temp_b5_11_25_i,temp_b5_27_9_r,temp_b5_27_9_i,temp_b5_27_25_r,temp_b5_27_25_i);
MULT MULT1194 (clk,temp_b4_11_10_r,temp_b4_11_10_i,temp_b4_11_26_r,temp_b4_11_26_i,temp_b4_27_10_r,temp_b4_27_10_i,temp_b4_27_26_r,temp_b4_27_26_i,temp_m5_11_10_r,temp_m5_11_10_i,temp_m5_11_26_r,temp_m5_11_26_i,temp_m5_27_10_r,temp_m5_27_10_i,temp_m5_27_26_r,temp_m5_27_26_i,`W9_real,`W9_imag,`W10_real,`W10_imag,`W19_real,`W19_imag);
butterfly butterfly1194 (clk,temp_m5_11_10_r,temp_m5_11_10_i,temp_m5_11_26_r,temp_m5_11_26_i,temp_m5_27_10_r,temp_m5_27_10_i,temp_m5_27_26_r,temp_m5_27_26_i,temp_b5_11_10_r,temp_b5_11_10_i,temp_b5_11_26_r,temp_b5_11_26_i,temp_b5_27_10_r,temp_b5_27_10_i,temp_b5_27_26_r,temp_b5_27_26_i);
MULT MULT1195 (clk,temp_b4_11_11_r,temp_b4_11_11_i,temp_b4_11_27_r,temp_b4_11_27_i,temp_b4_27_11_r,temp_b4_27_11_i,temp_b4_27_27_r,temp_b4_27_27_i,temp_m5_11_11_r,temp_m5_11_11_i,temp_m5_11_27_r,temp_m5_11_27_i,temp_m5_27_11_r,temp_m5_27_11_i,temp_m5_27_27_r,temp_m5_27_27_i,`W10_real,`W10_imag,`W10_real,`W10_imag,`W20_real,`W20_imag);
butterfly butterfly1195 (clk,temp_m5_11_11_r,temp_m5_11_11_i,temp_m5_11_27_r,temp_m5_11_27_i,temp_m5_27_11_r,temp_m5_27_11_i,temp_m5_27_27_r,temp_m5_27_27_i,temp_b5_11_11_r,temp_b5_11_11_i,temp_b5_11_27_r,temp_b5_11_27_i,temp_b5_27_11_r,temp_b5_27_11_i,temp_b5_27_27_r,temp_b5_27_27_i);
MULT MULT1196 (clk,temp_b4_11_12_r,temp_b4_11_12_i,temp_b4_11_28_r,temp_b4_11_28_i,temp_b4_27_12_r,temp_b4_27_12_i,temp_b4_27_28_r,temp_b4_27_28_i,temp_m5_11_12_r,temp_m5_11_12_i,temp_m5_11_28_r,temp_m5_11_28_i,temp_m5_27_12_r,temp_m5_27_12_i,temp_m5_27_28_r,temp_m5_27_28_i,`W11_real,`W11_imag,`W10_real,`W10_imag,`W21_real,`W21_imag);
butterfly butterfly1196 (clk,temp_m5_11_12_r,temp_m5_11_12_i,temp_m5_11_28_r,temp_m5_11_28_i,temp_m5_27_12_r,temp_m5_27_12_i,temp_m5_27_28_r,temp_m5_27_28_i,temp_b5_11_12_r,temp_b5_11_12_i,temp_b5_11_28_r,temp_b5_11_28_i,temp_b5_27_12_r,temp_b5_27_12_i,temp_b5_27_28_r,temp_b5_27_28_i);
MULT MULT1197 (clk,temp_b4_11_13_r,temp_b4_11_13_i,temp_b4_11_29_r,temp_b4_11_29_i,temp_b4_27_13_r,temp_b4_27_13_i,temp_b4_27_29_r,temp_b4_27_29_i,temp_m5_11_13_r,temp_m5_11_13_i,temp_m5_11_29_r,temp_m5_11_29_i,temp_m5_27_13_r,temp_m5_27_13_i,temp_m5_27_29_r,temp_m5_27_29_i,`W12_real,`W12_imag,`W10_real,`W10_imag,`W22_real,`W22_imag);
butterfly butterfly1197 (clk,temp_m5_11_13_r,temp_m5_11_13_i,temp_m5_11_29_r,temp_m5_11_29_i,temp_m5_27_13_r,temp_m5_27_13_i,temp_m5_27_29_r,temp_m5_27_29_i,temp_b5_11_13_r,temp_b5_11_13_i,temp_b5_11_29_r,temp_b5_11_29_i,temp_b5_27_13_r,temp_b5_27_13_i,temp_b5_27_29_r,temp_b5_27_29_i);
MULT MULT1198 (clk,temp_b4_11_14_r,temp_b4_11_14_i,temp_b4_11_30_r,temp_b4_11_30_i,temp_b4_27_14_r,temp_b4_27_14_i,temp_b4_27_30_r,temp_b4_27_30_i,temp_m5_11_14_r,temp_m5_11_14_i,temp_m5_11_30_r,temp_m5_11_30_i,temp_m5_27_14_r,temp_m5_27_14_i,temp_m5_27_30_r,temp_m5_27_30_i,`W13_real,`W13_imag,`W10_real,`W10_imag,`W23_real,`W23_imag);
butterfly butterfly1198 (clk,temp_m5_11_14_r,temp_m5_11_14_i,temp_m5_11_30_r,temp_m5_11_30_i,temp_m5_27_14_r,temp_m5_27_14_i,temp_m5_27_30_r,temp_m5_27_30_i,temp_b5_11_14_r,temp_b5_11_14_i,temp_b5_11_30_r,temp_b5_11_30_i,temp_b5_27_14_r,temp_b5_27_14_i,temp_b5_27_30_r,temp_b5_27_30_i);
MULT MULT1199 (clk,temp_b4_11_15_r,temp_b4_11_15_i,temp_b4_11_31_r,temp_b4_11_31_i,temp_b4_27_15_r,temp_b4_27_15_i,temp_b4_27_31_r,temp_b4_27_31_i,temp_m5_11_15_r,temp_m5_11_15_i,temp_m5_11_31_r,temp_m5_11_31_i,temp_m5_27_15_r,temp_m5_27_15_i,temp_m5_27_31_r,temp_m5_27_31_i,`W14_real,`W14_imag,`W10_real,`W10_imag,`W24_real,`W24_imag);
butterfly butterfly1199 (clk,temp_m5_11_15_r,temp_m5_11_15_i,temp_m5_11_31_r,temp_m5_11_31_i,temp_m5_27_15_r,temp_m5_27_15_i,temp_m5_27_31_r,temp_m5_27_31_i,temp_b5_11_15_r,temp_b5_11_15_i,temp_b5_11_31_r,temp_b5_11_31_i,temp_b5_27_15_r,temp_b5_27_15_i,temp_b5_27_31_r,temp_b5_27_31_i);
MULT MULT1200 (clk,temp_b4_11_16_r,temp_b4_11_16_i,temp_b4_11_32_r,temp_b4_11_32_i,temp_b4_27_16_r,temp_b4_27_16_i,temp_b4_27_32_r,temp_b4_27_32_i,temp_m5_11_16_r,temp_m5_11_16_i,temp_m5_11_32_r,temp_m5_11_32_i,temp_m5_27_16_r,temp_m5_27_16_i,temp_m5_27_32_r,temp_m5_27_32_i,`W15_real,`W15_imag,`W10_real,`W10_imag,`W25_real,`W25_imag);
butterfly butterfly1200 (clk,temp_m5_11_16_r,temp_m5_11_16_i,temp_m5_11_32_r,temp_m5_11_32_i,temp_m5_27_16_r,temp_m5_27_16_i,temp_m5_27_32_r,temp_m5_27_32_i,temp_b5_11_16_r,temp_b5_11_16_i,temp_b5_11_32_r,temp_b5_11_32_i,temp_b5_27_16_r,temp_b5_27_16_i,temp_b5_27_32_r,temp_b5_27_32_i);
MULT MULT1201 (clk,temp_b4_12_1_r,temp_b4_12_1_i,temp_b4_12_17_r,temp_b4_12_17_i,temp_b4_28_1_r,temp_b4_28_1_i,temp_b4_28_17_r,temp_b4_28_17_i,temp_m5_12_1_r,temp_m5_12_1_i,temp_m5_12_17_r,temp_m5_12_17_i,temp_m5_28_1_r,temp_m5_28_1_i,temp_m5_28_17_r,temp_m5_28_17_i,`W0_real,`W0_imag,`W11_real,`W11_imag,`W11_real,`W11_imag);
butterfly butterfly1201 (clk,temp_m5_12_1_r,temp_m5_12_1_i,temp_m5_12_17_r,temp_m5_12_17_i,temp_m5_28_1_r,temp_m5_28_1_i,temp_m5_28_17_r,temp_m5_28_17_i,temp_b5_12_1_r,temp_b5_12_1_i,temp_b5_12_17_r,temp_b5_12_17_i,temp_b5_28_1_r,temp_b5_28_1_i,temp_b5_28_17_r,temp_b5_28_17_i);
MULT MULT1202 (clk,temp_b4_12_2_r,temp_b4_12_2_i,temp_b4_12_18_r,temp_b4_12_18_i,temp_b4_28_2_r,temp_b4_28_2_i,temp_b4_28_18_r,temp_b4_28_18_i,temp_m5_12_2_r,temp_m5_12_2_i,temp_m5_12_18_r,temp_m5_12_18_i,temp_m5_28_2_r,temp_m5_28_2_i,temp_m5_28_18_r,temp_m5_28_18_i,`W1_real,`W1_imag,`W11_real,`W11_imag,`W12_real,`W12_imag);
butterfly butterfly1202 (clk,temp_m5_12_2_r,temp_m5_12_2_i,temp_m5_12_18_r,temp_m5_12_18_i,temp_m5_28_2_r,temp_m5_28_2_i,temp_m5_28_18_r,temp_m5_28_18_i,temp_b5_12_2_r,temp_b5_12_2_i,temp_b5_12_18_r,temp_b5_12_18_i,temp_b5_28_2_r,temp_b5_28_2_i,temp_b5_28_18_r,temp_b5_28_18_i);
MULT MULT1203 (clk,temp_b4_12_3_r,temp_b4_12_3_i,temp_b4_12_19_r,temp_b4_12_19_i,temp_b4_28_3_r,temp_b4_28_3_i,temp_b4_28_19_r,temp_b4_28_19_i,temp_m5_12_3_r,temp_m5_12_3_i,temp_m5_12_19_r,temp_m5_12_19_i,temp_m5_28_3_r,temp_m5_28_3_i,temp_m5_28_19_r,temp_m5_28_19_i,`W2_real,`W2_imag,`W11_real,`W11_imag,`W13_real,`W13_imag);
butterfly butterfly1203 (clk,temp_m5_12_3_r,temp_m5_12_3_i,temp_m5_12_19_r,temp_m5_12_19_i,temp_m5_28_3_r,temp_m5_28_3_i,temp_m5_28_19_r,temp_m5_28_19_i,temp_b5_12_3_r,temp_b5_12_3_i,temp_b5_12_19_r,temp_b5_12_19_i,temp_b5_28_3_r,temp_b5_28_3_i,temp_b5_28_19_r,temp_b5_28_19_i);
MULT MULT1204 (clk,temp_b4_12_4_r,temp_b4_12_4_i,temp_b4_12_20_r,temp_b4_12_20_i,temp_b4_28_4_r,temp_b4_28_4_i,temp_b4_28_20_r,temp_b4_28_20_i,temp_m5_12_4_r,temp_m5_12_4_i,temp_m5_12_20_r,temp_m5_12_20_i,temp_m5_28_4_r,temp_m5_28_4_i,temp_m5_28_20_r,temp_m5_28_20_i,`W3_real,`W3_imag,`W11_real,`W11_imag,`W14_real,`W14_imag);
butterfly butterfly1204 (clk,temp_m5_12_4_r,temp_m5_12_4_i,temp_m5_12_20_r,temp_m5_12_20_i,temp_m5_28_4_r,temp_m5_28_4_i,temp_m5_28_20_r,temp_m5_28_20_i,temp_b5_12_4_r,temp_b5_12_4_i,temp_b5_12_20_r,temp_b5_12_20_i,temp_b5_28_4_r,temp_b5_28_4_i,temp_b5_28_20_r,temp_b5_28_20_i);
MULT MULT1205 (clk,temp_b4_12_5_r,temp_b4_12_5_i,temp_b4_12_21_r,temp_b4_12_21_i,temp_b4_28_5_r,temp_b4_28_5_i,temp_b4_28_21_r,temp_b4_28_21_i,temp_m5_12_5_r,temp_m5_12_5_i,temp_m5_12_21_r,temp_m5_12_21_i,temp_m5_28_5_r,temp_m5_28_5_i,temp_m5_28_21_r,temp_m5_28_21_i,`W4_real,`W4_imag,`W11_real,`W11_imag,`W15_real,`W15_imag);
butterfly butterfly1205 (clk,temp_m5_12_5_r,temp_m5_12_5_i,temp_m5_12_21_r,temp_m5_12_21_i,temp_m5_28_5_r,temp_m5_28_5_i,temp_m5_28_21_r,temp_m5_28_21_i,temp_b5_12_5_r,temp_b5_12_5_i,temp_b5_12_21_r,temp_b5_12_21_i,temp_b5_28_5_r,temp_b5_28_5_i,temp_b5_28_21_r,temp_b5_28_21_i);
MULT MULT1206 (clk,temp_b4_12_6_r,temp_b4_12_6_i,temp_b4_12_22_r,temp_b4_12_22_i,temp_b4_28_6_r,temp_b4_28_6_i,temp_b4_28_22_r,temp_b4_28_22_i,temp_m5_12_6_r,temp_m5_12_6_i,temp_m5_12_22_r,temp_m5_12_22_i,temp_m5_28_6_r,temp_m5_28_6_i,temp_m5_28_22_r,temp_m5_28_22_i,`W5_real,`W5_imag,`W11_real,`W11_imag,`W16_real,`W16_imag);
butterfly butterfly1206 (clk,temp_m5_12_6_r,temp_m5_12_6_i,temp_m5_12_22_r,temp_m5_12_22_i,temp_m5_28_6_r,temp_m5_28_6_i,temp_m5_28_22_r,temp_m5_28_22_i,temp_b5_12_6_r,temp_b5_12_6_i,temp_b5_12_22_r,temp_b5_12_22_i,temp_b5_28_6_r,temp_b5_28_6_i,temp_b5_28_22_r,temp_b5_28_22_i);
MULT MULT1207 (clk,temp_b4_12_7_r,temp_b4_12_7_i,temp_b4_12_23_r,temp_b4_12_23_i,temp_b4_28_7_r,temp_b4_28_7_i,temp_b4_28_23_r,temp_b4_28_23_i,temp_m5_12_7_r,temp_m5_12_7_i,temp_m5_12_23_r,temp_m5_12_23_i,temp_m5_28_7_r,temp_m5_28_7_i,temp_m5_28_23_r,temp_m5_28_23_i,`W6_real,`W6_imag,`W11_real,`W11_imag,`W17_real,`W17_imag);
butterfly butterfly1207 (clk,temp_m5_12_7_r,temp_m5_12_7_i,temp_m5_12_23_r,temp_m5_12_23_i,temp_m5_28_7_r,temp_m5_28_7_i,temp_m5_28_23_r,temp_m5_28_23_i,temp_b5_12_7_r,temp_b5_12_7_i,temp_b5_12_23_r,temp_b5_12_23_i,temp_b5_28_7_r,temp_b5_28_7_i,temp_b5_28_23_r,temp_b5_28_23_i);
MULT MULT1208 (clk,temp_b4_12_8_r,temp_b4_12_8_i,temp_b4_12_24_r,temp_b4_12_24_i,temp_b4_28_8_r,temp_b4_28_8_i,temp_b4_28_24_r,temp_b4_28_24_i,temp_m5_12_8_r,temp_m5_12_8_i,temp_m5_12_24_r,temp_m5_12_24_i,temp_m5_28_8_r,temp_m5_28_8_i,temp_m5_28_24_r,temp_m5_28_24_i,`W7_real,`W7_imag,`W11_real,`W11_imag,`W18_real,`W18_imag);
butterfly butterfly1208 (clk,temp_m5_12_8_r,temp_m5_12_8_i,temp_m5_12_24_r,temp_m5_12_24_i,temp_m5_28_8_r,temp_m5_28_8_i,temp_m5_28_24_r,temp_m5_28_24_i,temp_b5_12_8_r,temp_b5_12_8_i,temp_b5_12_24_r,temp_b5_12_24_i,temp_b5_28_8_r,temp_b5_28_8_i,temp_b5_28_24_r,temp_b5_28_24_i);
MULT MULT1209 (clk,temp_b4_12_9_r,temp_b4_12_9_i,temp_b4_12_25_r,temp_b4_12_25_i,temp_b4_28_9_r,temp_b4_28_9_i,temp_b4_28_25_r,temp_b4_28_25_i,temp_m5_12_9_r,temp_m5_12_9_i,temp_m5_12_25_r,temp_m5_12_25_i,temp_m5_28_9_r,temp_m5_28_9_i,temp_m5_28_25_r,temp_m5_28_25_i,`W8_real,`W8_imag,`W11_real,`W11_imag,`W19_real,`W19_imag);
butterfly butterfly1209 (clk,temp_m5_12_9_r,temp_m5_12_9_i,temp_m5_12_25_r,temp_m5_12_25_i,temp_m5_28_9_r,temp_m5_28_9_i,temp_m5_28_25_r,temp_m5_28_25_i,temp_b5_12_9_r,temp_b5_12_9_i,temp_b5_12_25_r,temp_b5_12_25_i,temp_b5_28_9_r,temp_b5_28_9_i,temp_b5_28_25_r,temp_b5_28_25_i);
MULT MULT1210 (clk,temp_b4_12_10_r,temp_b4_12_10_i,temp_b4_12_26_r,temp_b4_12_26_i,temp_b4_28_10_r,temp_b4_28_10_i,temp_b4_28_26_r,temp_b4_28_26_i,temp_m5_12_10_r,temp_m5_12_10_i,temp_m5_12_26_r,temp_m5_12_26_i,temp_m5_28_10_r,temp_m5_28_10_i,temp_m5_28_26_r,temp_m5_28_26_i,`W9_real,`W9_imag,`W11_real,`W11_imag,`W20_real,`W20_imag);
butterfly butterfly1210 (clk,temp_m5_12_10_r,temp_m5_12_10_i,temp_m5_12_26_r,temp_m5_12_26_i,temp_m5_28_10_r,temp_m5_28_10_i,temp_m5_28_26_r,temp_m5_28_26_i,temp_b5_12_10_r,temp_b5_12_10_i,temp_b5_12_26_r,temp_b5_12_26_i,temp_b5_28_10_r,temp_b5_28_10_i,temp_b5_28_26_r,temp_b5_28_26_i);
MULT MULT1211 (clk,temp_b4_12_11_r,temp_b4_12_11_i,temp_b4_12_27_r,temp_b4_12_27_i,temp_b4_28_11_r,temp_b4_28_11_i,temp_b4_28_27_r,temp_b4_28_27_i,temp_m5_12_11_r,temp_m5_12_11_i,temp_m5_12_27_r,temp_m5_12_27_i,temp_m5_28_11_r,temp_m5_28_11_i,temp_m5_28_27_r,temp_m5_28_27_i,`W10_real,`W10_imag,`W11_real,`W11_imag,`W21_real,`W21_imag);
butterfly butterfly1211 (clk,temp_m5_12_11_r,temp_m5_12_11_i,temp_m5_12_27_r,temp_m5_12_27_i,temp_m5_28_11_r,temp_m5_28_11_i,temp_m5_28_27_r,temp_m5_28_27_i,temp_b5_12_11_r,temp_b5_12_11_i,temp_b5_12_27_r,temp_b5_12_27_i,temp_b5_28_11_r,temp_b5_28_11_i,temp_b5_28_27_r,temp_b5_28_27_i);
MULT MULT1212 (clk,temp_b4_12_12_r,temp_b4_12_12_i,temp_b4_12_28_r,temp_b4_12_28_i,temp_b4_28_12_r,temp_b4_28_12_i,temp_b4_28_28_r,temp_b4_28_28_i,temp_m5_12_12_r,temp_m5_12_12_i,temp_m5_12_28_r,temp_m5_12_28_i,temp_m5_28_12_r,temp_m5_28_12_i,temp_m5_28_28_r,temp_m5_28_28_i,`W11_real,`W11_imag,`W11_real,`W11_imag,`W22_real,`W22_imag);
butterfly butterfly1212 (clk,temp_m5_12_12_r,temp_m5_12_12_i,temp_m5_12_28_r,temp_m5_12_28_i,temp_m5_28_12_r,temp_m5_28_12_i,temp_m5_28_28_r,temp_m5_28_28_i,temp_b5_12_12_r,temp_b5_12_12_i,temp_b5_12_28_r,temp_b5_12_28_i,temp_b5_28_12_r,temp_b5_28_12_i,temp_b5_28_28_r,temp_b5_28_28_i);
MULT MULT1213 (clk,temp_b4_12_13_r,temp_b4_12_13_i,temp_b4_12_29_r,temp_b4_12_29_i,temp_b4_28_13_r,temp_b4_28_13_i,temp_b4_28_29_r,temp_b4_28_29_i,temp_m5_12_13_r,temp_m5_12_13_i,temp_m5_12_29_r,temp_m5_12_29_i,temp_m5_28_13_r,temp_m5_28_13_i,temp_m5_28_29_r,temp_m5_28_29_i,`W12_real,`W12_imag,`W11_real,`W11_imag,`W23_real,`W23_imag);
butterfly butterfly1213 (clk,temp_m5_12_13_r,temp_m5_12_13_i,temp_m5_12_29_r,temp_m5_12_29_i,temp_m5_28_13_r,temp_m5_28_13_i,temp_m5_28_29_r,temp_m5_28_29_i,temp_b5_12_13_r,temp_b5_12_13_i,temp_b5_12_29_r,temp_b5_12_29_i,temp_b5_28_13_r,temp_b5_28_13_i,temp_b5_28_29_r,temp_b5_28_29_i);
MULT MULT1214 (clk,temp_b4_12_14_r,temp_b4_12_14_i,temp_b4_12_30_r,temp_b4_12_30_i,temp_b4_28_14_r,temp_b4_28_14_i,temp_b4_28_30_r,temp_b4_28_30_i,temp_m5_12_14_r,temp_m5_12_14_i,temp_m5_12_30_r,temp_m5_12_30_i,temp_m5_28_14_r,temp_m5_28_14_i,temp_m5_28_30_r,temp_m5_28_30_i,`W13_real,`W13_imag,`W11_real,`W11_imag,`W24_real,`W24_imag);
butterfly butterfly1214 (clk,temp_m5_12_14_r,temp_m5_12_14_i,temp_m5_12_30_r,temp_m5_12_30_i,temp_m5_28_14_r,temp_m5_28_14_i,temp_m5_28_30_r,temp_m5_28_30_i,temp_b5_12_14_r,temp_b5_12_14_i,temp_b5_12_30_r,temp_b5_12_30_i,temp_b5_28_14_r,temp_b5_28_14_i,temp_b5_28_30_r,temp_b5_28_30_i);
MULT MULT1215 (clk,temp_b4_12_15_r,temp_b4_12_15_i,temp_b4_12_31_r,temp_b4_12_31_i,temp_b4_28_15_r,temp_b4_28_15_i,temp_b4_28_31_r,temp_b4_28_31_i,temp_m5_12_15_r,temp_m5_12_15_i,temp_m5_12_31_r,temp_m5_12_31_i,temp_m5_28_15_r,temp_m5_28_15_i,temp_m5_28_31_r,temp_m5_28_31_i,`W14_real,`W14_imag,`W11_real,`W11_imag,`W25_real,`W25_imag);
butterfly butterfly1215 (clk,temp_m5_12_15_r,temp_m5_12_15_i,temp_m5_12_31_r,temp_m5_12_31_i,temp_m5_28_15_r,temp_m5_28_15_i,temp_m5_28_31_r,temp_m5_28_31_i,temp_b5_12_15_r,temp_b5_12_15_i,temp_b5_12_31_r,temp_b5_12_31_i,temp_b5_28_15_r,temp_b5_28_15_i,temp_b5_28_31_r,temp_b5_28_31_i);
MULT MULT1216 (clk,temp_b4_12_16_r,temp_b4_12_16_i,temp_b4_12_32_r,temp_b4_12_32_i,temp_b4_28_16_r,temp_b4_28_16_i,temp_b4_28_32_r,temp_b4_28_32_i,temp_m5_12_16_r,temp_m5_12_16_i,temp_m5_12_32_r,temp_m5_12_32_i,temp_m5_28_16_r,temp_m5_28_16_i,temp_m5_28_32_r,temp_m5_28_32_i,`W15_real,`W15_imag,`W11_real,`W11_imag,`W26_real,`W26_imag);
butterfly butterfly1216 (clk,temp_m5_12_16_r,temp_m5_12_16_i,temp_m5_12_32_r,temp_m5_12_32_i,temp_m5_28_16_r,temp_m5_28_16_i,temp_m5_28_32_r,temp_m5_28_32_i,temp_b5_12_16_r,temp_b5_12_16_i,temp_b5_12_32_r,temp_b5_12_32_i,temp_b5_28_16_r,temp_b5_28_16_i,temp_b5_28_32_r,temp_b5_28_32_i);
MULT MULT1217 (clk,temp_b4_13_1_r,temp_b4_13_1_i,temp_b4_13_17_r,temp_b4_13_17_i,temp_b4_29_1_r,temp_b4_29_1_i,temp_b4_29_17_r,temp_b4_29_17_i,temp_m5_13_1_r,temp_m5_13_1_i,temp_m5_13_17_r,temp_m5_13_17_i,temp_m5_29_1_r,temp_m5_29_1_i,temp_m5_29_17_r,temp_m5_29_17_i,`W0_real,`W0_imag,`W12_real,`W12_imag,`W12_real,`W12_imag);
butterfly butterfly1217 (clk,temp_m5_13_1_r,temp_m5_13_1_i,temp_m5_13_17_r,temp_m5_13_17_i,temp_m5_29_1_r,temp_m5_29_1_i,temp_m5_29_17_r,temp_m5_29_17_i,temp_b5_13_1_r,temp_b5_13_1_i,temp_b5_13_17_r,temp_b5_13_17_i,temp_b5_29_1_r,temp_b5_29_1_i,temp_b5_29_17_r,temp_b5_29_17_i);
MULT MULT1218 (clk,temp_b4_13_2_r,temp_b4_13_2_i,temp_b4_13_18_r,temp_b4_13_18_i,temp_b4_29_2_r,temp_b4_29_2_i,temp_b4_29_18_r,temp_b4_29_18_i,temp_m5_13_2_r,temp_m5_13_2_i,temp_m5_13_18_r,temp_m5_13_18_i,temp_m5_29_2_r,temp_m5_29_2_i,temp_m5_29_18_r,temp_m5_29_18_i,`W1_real,`W1_imag,`W12_real,`W12_imag,`W13_real,`W13_imag);
butterfly butterfly1218 (clk,temp_m5_13_2_r,temp_m5_13_2_i,temp_m5_13_18_r,temp_m5_13_18_i,temp_m5_29_2_r,temp_m5_29_2_i,temp_m5_29_18_r,temp_m5_29_18_i,temp_b5_13_2_r,temp_b5_13_2_i,temp_b5_13_18_r,temp_b5_13_18_i,temp_b5_29_2_r,temp_b5_29_2_i,temp_b5_29_18_r,temp_b5_29_18_i);
MULT MULT1219 (clk,temp_b4_13_3_r,temp_b4_13_3_i,temp_b4_13_19_r,temp_b4_13_19_i,temp_b4_29_3_r,temp_b4_29_3_i,temp_b4_29_19_r,temp_b4_29_19_i,temp_m5_13_3_r,temp_m5_13_3_i,temp_m5_13_19_r,temp_m5_13_19_i,temp_m5_29_3_r,temp_m5_29_3_i,temp_m5_29_19_r,temp_m5_29_19_i,`W2_real,`W2_imag,`W12_real,`W12_imag,`W14_real,`W14_imag);
butterfly butterfly1219 (clk,temp_m5_13_3_r,temp_m5_13_3_i,temp_m5_13_19_r,temp_m5_13_19_i,temp_m5_29_3_r,temp_m5_29_3_i,temp_m5_29_19_r,temp_m5_29_19_i,temp_b5_13_3_r,temp_b5_13_3_i,temp_b5_13_19_r,temp_b5_13_19_i,temp_b5_29_3_r,temp_b5_29_3_i,temp_b5_29_19_r,temp_b5_29_19_i);
MULT MULT1220 (clk,temp_b4_13_4_r,temp_b4_13_4_i,temp_b4_13_20_r,temp_b4_13_20_i,temp_b4_29_4_r,temp_b4_29_4_i,temp_b4_29_20_r,temp_b4_29_20_i,temp_m5_13_4_r,temp_m5_13_4_i,temp_m5_13_20_r,temp_m5_13_20_i,temp_m5_29_4_r,temp_m5_29_4_i,temp_m5_29_20_r,temp_m5_29_20_i,`W3_real,`W3_imag,`W12_real,`W12_imag,`W15_real,`W15_imag);
butterfly butterfly1220 (clk,temp_m5_13_4_r,temp_m5_13_4_i,temp_m5_13_20_r,temp_m5_13_20_i,temp_m5_29_4_r,temp_m5_29_4_i,temp_m5_29_20_r,temp_m5_29_20_i,temp_b5_13_4_r,temp_b5_13_4_i,temp_b5_13_20_r,temp_b5_13_20_i,temp_b5_29_4_r,temp_b5_29_4_i,temp_b5_29_20_r,temp_b5_29_20_i);
MULT MULT1221 (clk,temp_b4_13_5_r,temp_b4_13_5_i,temp_b4_13_21_r,temp_b4_13_21_i,temp_b4_29_5_r,temp_b4_29_5_i,temp_b4_29_21_r,temp_b4_29_21_i,temp_m5_13_5_r,temp_m5_13_5_i,temp_m5_13_21_r,temp_m5_13_21_i,temp_m5_29_5_r,temp_m5_29_5_i,temp_m5_29_21_r,temp_m5_29_21_i,`W4_real,`W4_imag,`W12_real,`W12_imag,`W16_real,`W16_imag);
butterfly butterfly1221 (clk,temp_m5_13_5_r,temp_m5_13_5_i,temp_m5_13_21_r,temp_m5_13_21_i,temp_m5_29_5_r,temp_m5_29_5_i,temp_m5_29_21_r,temp_m5_29_21_i,temp_b5_13_5_r,temp_b5_13_5_i,temp_b5_13_21_r,temp_b5_13_21_i,temp_b5_29_5_r,temp_b5_29_5_i,temp_b5_29_21_r,temp_b5_29_21_i);
MULT MULT1222 (clk,temp_b4_13_6_r,temp_b4_13_6_i,temp_b4_13_22_r,temp_b4_13_22_i,temp_b4_29_6_r,temp_b4_29_6_i,temp_b4_29_22_r,temp_b4_29_22_i,temp_m5_13_6_r,temp_m5_13_6_i,temp_m5_13_22_r,temp_m5_13_22_i,temp_m5_29_6_r,temp_m5_29_6_i,temp_m5_29_22_r,temp_m5_29_22_i,`W5_real,`W5_imag,`W12_real,`W12_imag,`W17_real,`W17_imag);
butterfly butterfly1222 (clk,temp_m5_13_6_r,temp_m5_13_6_i,temp_m5_13_22_r,temp_m5_13_22_i,temp_m5_29_6_r,temp_m5_29_6_i,temp_m5_29_22_r,temp_m5_29_22_i,temp_b5_13_6_r,temp_b5_13_6_i,temp_b5_13_22_r,temp_b5_13_22_i,temp_b5_29_6_r,temp_b5_29_6_i,temp_b5_29_22_r,temp_b5_29_22_i);
MULT MULT1223 (clk,temp_b4_13_7_r,temp_b4_13_7_i,temp_b4_13_23_r,temp_b4_13_23_i,temp_b4_29_7_r,temp_b4_29_7_i,temp_b4_29_23_r,temp_b4_29_23_i,temp_m5_13_7_r,temp_m5_13_7_i,temp_m5_13_23_r,temp_m5_13_23_i,temp_m5_29_7_r,temp_m5_29_7_i,temp_m5_29_23_r,temp_m5_29_23_i,`W6_real,`W6_imag,`W12_real,`W12_imag,`W18_real,`W18_imag);
butterfly butterfly1223 (clk,temp_m5_13_7_r,temp_m5_13_7_i,temp_m5_13_23_r,temp_m5_13_23_i,temp_m5_29_7_r,temp_m5_29_7_i,temp_m5_29_23_r,temp_m5_29_23_i,temp_b5_13_7_r,temp_b5_13_7_i,temp_b5_13_23_r,temp_b5_13_23_i,temp_b5_29_7_r,temp_b5_29_7_i,temp_b5_29_23_r,temp_b5_29_23_i);
MULT MULT1224 (clk,temp_b4_13_8_r,temp_b4_13_8_i,temp_b4_13_24_r,temp_b4_13_24_i,temp_b4_29_8_r,temp_b4_29_8_i,temp_b4_29_24_r,temp_b4_29_24_i,temp_m5_13_8_r,temp_m5_13_8_i,temp_m5_13_24_r,temp_m5_13_24_i,temp_m5_29_8_r,temp_m5_29_8_i,temp_m5_29_24_r,temp_m5_29_24_i,`W7_real,`W7_imag,`W12_real,`W12_imag,`W19_real,`W19_imag);
butterfly butterfly1224 (clk,temp_m5_13_8_r,temp_m5_13_8_i,temp_m5_13_24_r,temp_m5_13_24_i,temp_m5_29_8_r,temp_m5_29_8_i,temp_m5_29_24_r,temp_m5_29_24_i,temp_b5_13_8_r,temp_b5_13_8_i,temp_b5_13_24_r,temp_b5_13_24_i,temp_b5_29_8_r,temp_b5_29_8_i,temp_b5_29_24_r,temp_b5_29_24_i);
MULT MULT1225 (clk,temp_b4_13_9_r,temp_b4_13_9_i,temp_b4_13_25_r,temp_b4_13_25_i,temp_b4_29_9_r,temp_b4_29_9_i,temp_b4_29_25_r,temp_b4_29_25_i,temp_m5_13_9_r,temp_m5_13_9_i,temp_m5_13_25_r,temp_m5_13_25_i,temp_m5_29_9_r,temp_m5_29_9_i,temp_m5_29_25_r,temp_m5_29_25_i,`W8_real,`W8_imag,`W12_real,`W12_imag,`W20_real,`W20_imag);
butterfly butterfly1225 (clk,temp_m5_13_9_r,temp_m5_13_9_i,temp_m5_13_25_r,temp_m5_13_25_i,temp_m5_29_9_r,temp_m5_29_9_i,temp_m5_29_25_r,temp_m5_29_25_i,temp_b5_13_9_r,temp_b5_13_9_i,temp_b5_13_25_r,temp_b5_13_25_i,temp_b5_29_9_r,temp_b5_29_9_i,temp_b5_29_25_r,temp_b5_29_25_i);
MULT MULT1226 (clk,temp_b4_13_10_r,temp_b4_13_10_i,temp_b4_13_26_r,temp_b4_13_26_i,temp_b4_29_10_r,temp_b4_29_10_i,temp_b4_29_26_r,temp_b4_29_26_i,temp_m5_13_10_r,temp_m5_13_10_i,temp_m5_13_26_r,temp_m5_13_26_i,temp_m5_29_10_r,temp_m5_29_10_i,temp_m5_29_26_r,temp_m5_29_26_i,`W9_real,`W9_imag,`W12_real,`W12_imag,`W21_real,`W21_imag);
butterfly butterfly1226 (clk,temp_m5_13_10_r,temp_m5_13_10_i,temp_m5_13_26_r,temp_m5_13_26_i,temp_m5_29_10_r,temp_m5_29_10_i,temp_m5_29_26_r,temp_m5_29_26_i,temp_b5_13_10_r,temp_b5_13_10_i,temp_b5_13_26_r,temp_b5_13_26_i,temp_b5_29_10_r,temp_b5_29_10_i,temp_b5_29_26_r,temp_b5_29_26_i);
MULT MULT1227 (clk,temp_b4_13_11_r,temp_b4_13_11_i,temp_b4_13_27_r,temp_b4_13_27_i,temp_b4_29_11_r,temp_b4_29_11_i,temp_b4_29_27_r,temp_b4_29_27_i,temp_m5_13_11_r,temp_m5_13_11_i,temp_m5_13_27_r,temp_m5_13_27_i,temp_m5_29_11_r,temp_m5_29_11_i,temp_m5_29_27_r,temp_m5_29_27_i,`W10_real,`W10_imag,`W12_real,`W12_imag,`W22_real,`W22_imag);
butterfly butterfly1227 (clk,temp_m5_13_11_r,temp_m5_13_11_i,temp_m5_13_27_r,temp_m5_13_27_i,temp_m5_29_11_r,temp_m5_29_11_i,temp_m5_29_27_r,temp_m5_29_27_i,temp_b5_13_11_r,temp_b5_13_11_i,temp_b5_13_27_r,temp_b5_13_27_i,temp_b5_29_11_r,temp_b5_29_11_i,temp_b5_29_27_r,temp_b5_29_27_i);
MULT MULT1228 (clk,temp_b4_13_12_r,temp_b4_13_12_i,temp_b4_13_28_r,temp_b4_13_28_i,temp_b4_29_12_r,temp_b4_29_12_i,temp_b4_29_28_r,temp_b4_29_28_i,temp_m5_13_12_r,temp_m5_13_12_i,temp_m5_13_28_r,temp_m5_13_28_i,temp_m5_29_12_r,temp_m5_29_12_i,temp_m5_29_28_r,temp_m5_29_28_i,`W11_real,`W11_imag,`W12_real,`W12_imag,`W23_real,`W23_imag);
butterfly butterfly1228 (clk,temp_m5_13_12_r,temp_m5_13_12_i,temp_m5_13_28_r,temp_m5_13_28_i,temp_m5_29_12_r,temp_m5_29_12_i,temp_m5_29_28_r,temp_m5_29_28_i,temp_b5_13_12_r,temp_b5_13_12_i,temp_b5_13_28_r,temp_b5_13_28_i,temp_b5_29_12_r,temp_b5_29_12_i,temp_b5_29_28_r,temp_b5_29_28_i);
MULT MULT1229 (clk,temp_b4_13_13_r,temp_b4_13_13_i,temp_b4_13_29_r,temp_b4_13_29_i,temp_b4_29_13_r,temp_b4_29_13_i,temp_b4_29_29_r,temp_b4_29_29_i,temp_m5_13_13_r,temp_m5_13_13_i,temp_m5_13_29_r,temp_m5_13_29_i,temp_m5_29_13_r,temp_m5_29_13_i,temp_m5_29_29_r,temp_m5_29_29_i,`W12_real,`W12_imag,`W12_real,`W12_imag,`W24_real,`W24_imag);
butterfly butterfly1229 (clk,temp_m5_13_13_r,temp_m5_13_13_i,temp_m5_13_29_r,temp_m5_13_29_i,temp_m5_29_13_r,temp_m5_29_13_i,temp_m5_29_29_r,temp_m5_29_29_i,temp_b5_13_13_r,temp_b5_13_13_i,temp_b5_13_29_r,temp_b5_13_29_i,temp_b5_29_13_r,temp_b5_29_13_i,temp_b5_29_29_r,temp_b5_29_29_i);
MULT MULT1230 (clk,temp_b4_13_14_r,temp_b4_13_14_i,temp_b4_13_30_r,temp_b4_13_30_i,temp_b4_29_14_r,temp_b4_29_14_i,temp_b4_29_30_r,temp_b4_29_30_i,temp_m5_13_14_r,temp_m5_13_14_i,temp_m5_13_30_r,temp_m5_13_30_i,temp_m5_29_14_r,temp_m5_29_14_i,temp_m5_29_30_r,temp_m5_29_30_i,`W13_real,`W13_imag,`W12_real,`W12_imag,`W25_real,`W25_imag);
butterfly butterfly1230 (clk,temp_m5_13_14_r,temp_m5_13_14_i,temp_m5_13_30_r,temp_m5_13_30_i,temp_m5_29_14_r,temp_m5_29_14_i,temp_m5_29_30_r,temp_m5_29_30_i,temp_b5_13_14_r,temp_b5_13_14_i,temp_b5_13_30_r,temp_b5_13_30_i,temp_b5_29_14_r,temp_b5_29_14_i,temp_b5_29_30_r,temp_b5_29_30_i);
MULT MULT1231 (clk,temp_b4_13_15_r,temp_b4_13_15_i,temp_b4_13_31_r,temp_b4_13_31_i,temp_b4_29_15_r,temp_b4_29_15_i,temp_b4_29_31_r,temp_b4_29_31_i,temp_m5_13_15_r,temp_m5_13_15_i,temp_m5_13_31_r,temp_m5_13_31_i,temp_m5_29_15_r,temp_m5_29_15_i,temp_m5_29_31_r,temp_m5_29_31_i,`W14_real,`W14_imag,`W12_real,`W12_imag,`W26_real,`W26_imag);
butterfly butterfly1231 (clk,temp_m5_13_15_r,temp_m5_13_15_i,temp_m5_13_31_r,temp_m5_13_31_i,temp_m5_29_15_r,temp_m5_29_15_i,temp_m5_29_31_r,temp_m5_29_31_i,temp_b5_13_15_r,temp_b5_13_15_i,temp_b5_13_31_r,temp_b5_13_31_i,temp_b5_29_15_r,temp_b5_29_15_i,temp_b5_29_31_r,temp_b5_29_31_i);
MULT MULT1232 (clk,temp_b4_13_16_r,temp_b4_13_16_i,temp_b4_13_32_r,temp_b4_13_32_i,temp_b4_29_16_r,temp_b4_29_16_i,temp_b4_29_32_r,temp_b4_29_32_i,temp_m5_13_16_r,temp_m5_13_16_i,temp_m5_13_32_r,temp_m5_13_32_i,temp_m5_29_16_r,temp_m5_29_16_i,temp_m5_29_32_r,temp_m5_29_32_i,`W15_real,`W15_imag,`W12_real,`W12_imag,`W27_real,`W27_imag);
butterfly butterfly1232 (clk,temp_m5_13_16_r,temp_m5_13_16_i,temp_m5_13_32_r,temp_m5_13_32_i,temp_m5_29_16_r,temp_m5_29_16_i,temp_m5_29_32_r,temp_m5_29_32_i,temp_b5_13_16_r,temp_b5_13_16_i,temp_b5_13_32_r,temp_b5_13_32_i,temp_b5_29_16_r,temp_b5_29_16_i,temp_b5_29_32_r,temp_b5_29_32_i);
MULT MULT1233 (clk,temp_b4_14_1_r,temp_b4_14_1_i,temp_b4_14_17_r,temp_b4_14_17_i,temp_b4_30_1_r,temp_b4_30_1_i,temp_b4_30_17_r,temp_b4_30_17_i,temp_m5_14_1_r,temp_m5_14_1_i,temp_m5_14_17_r,temp_m5_14_17_i,temp_m5_30_1_r,temp_m5_30_1_i,temp_m5_30_17_r,temp_m5_30_17_i,`W0_real,`W0_imag,`W13_real,`W13_imag,`W13_real,`W13_imag);
butterfly butterfly1233 (clk,temp_m5_14_1_r,temp_m5_14_1_i,temp_m5_14_17_r,temp_m5_14_17_i,temp_m5_30_1_r,temp_m5_30_1_i,temp_m5_30_17_r,temp_m5_30_17_i,temp_b5_14_1_r,temp_b5_14_1_i,temp_b5_14_17_r,temp_b5_14_17_i,temp_b5_30_1_r,temp_b5_30_1_i,temp_b5_30_17_r,temp_b5_30_17_i);
MULT MULT1234 (clk,temp_b4_14_2_r,temp_b4_14_2_i,temp_b4_14_18_r,temp_b4_14_18_i,temp_b4_30_2_r,temp_b4_30_2_i,temp_b4_30_18_r,temp_b4_30_18_i,temp_m5_14_2_r,temp_m5_14_2_i,temp_m5_14_18_r,temp_m5_14_18_i,temp_m5_30_2_r,temp_m5_30_2_i,temp_m5_30_18_r,temp_m5_30_18_i,`W1_real,`W1_imag,`W13_real,`W13_imag,`W14_real,`W14_imag);
butterfly butterfly1234 (clk,temp_m5_14_2_r,temp_m5_14_2_i,temp_m5_14_18_r,temp_m5_14_18_i,temp_m5_30_2_r,temp_m5_30_2_i,temp_m5_30_18_r,temp_m5_30_18_i,temp_b5_14_2_r,temp_b5_14_2_i,temp_b5_14_18_r,temp_b5_14_18_i,temp_b5_30_2_r,temp_b5_30_2_i,temp_b5_30_18_r,temp_b5_30_18_i);
MULT MULT1235 (clk,temp_b4_14_3_r,temp_b4_14_3_i,temp_b4_14_19_r,temp_b4_14_19_i,temp_b4_30_3_r,temp_b4_30_3_i,temp_b4_30_19_r,temp_b4_30_19_i,temp_m5_14_3_r,temp_m5_14_3_i,temp_m5_14_19_r,temp_m5_14_19_i,temp_m5_30_3_r,temp_m5_30_3_i,temp_m5_30_19_r,temp_m5_30_19_i,`W2_real,`W2_imag,`W13_real,`W13_imag,`W15_real,`W15_imag);
butterfly butterfly1235 (clk,temp_m5_14_3_r,temp_m5_14_3_i,temp_m5_14_19_r,temp_m5_14_19_i,temp_m5_30_3_r,temp_m5_30_3_i,temp_m5_30_19_r,temp_m5_30_19_i,temp_b5_14_3_r,temp_b5_14_3_i,temp_b5_14_19_r,temp_b5_14_19_i,temp_b5_30_3_r,temp_b5_30_3_i,temp_b5_30_19_r,temp_b5_30_19_i);
MULT MULT1236 (clk,temp_b4_14_4_r,temp_b4_14_4_i,temp_b4_14_20_r,temp_b4_14_20_i,temp_b4_30_4_r,temp_b4_30_4_i,temp_b4_30_20_r,temp_b4_30_20_i,temp_m5_14_4_r,temp_m5_14_4_i,temp_m5_14_20_r,temp_m5_14_20_i,temp_m5_30_4_r,temp_m5_30_4_i,temp_m5_30_20_r,temp_m5_30_20_i,`W3_real,`W3_imag,`W13_real,`W13_imag,`W16_real,`W16_imag);
butterfly butterfly1236 (clk,temp_m5_14_4_r,temp_m5_14_4_i,temp_m5_14_20_r,temp_m5_14_20_i,temp_m5_30_4_r,temp_m5_30_4_i,temp_m5_30_20_r,temp_m5_30_20_i,temp_b5_14_4_r,temp_b5_14_4_i,temp_b5_14_20_r,temp_b5_14_20_i,temp_b5_30_4_r,temp_b5_30_4_i,temp_b5_30_20_r,temp_b5_30_20_i);
MULT MULT1237 (clk,temp_b4_14_5_r,temp_b4_14_5_i,temp_b4_14_21_r,temp_b4_14_21_i,temp_b4_30_5_r,temp_b4_30_5_i,temp_b4_30_21_r,temp_b4_30_21_i,temp_m5_14_5_r,temp_m5_14_5_i,temp_m5_14_21_r,temp_m5_14_21_i,temp_m5_30_5_r,temp_m5_30_5_i,temp_m5_30_21_r,temp_m5_30_21_i,`W4_real,`W4_imag,`W13_real,`W13_imag,`W17_real,`W17_imag);
butterfly butterfly1237 (clk,temp_m5_14_5_r,temp_m5_14_5_i,temp_m5_14_21_r,temp_m5_14_21_i,temp_m5_30_5_r,temp_m5_30_5_i,temp_m5_30_21_r,temp_m5_30_21_i,temp_b5_14_5_r,temp_b5_14_5_i,temp_b5_14_21_r,temp_b5_14_21_i,temp_b5_30_5_r,temp_b5_30_5_i,temp_b5_30_21_r,temp_b5_30_21_i);
MULT MULT1238 (clk,temp_b4_14_6_r,temp_b4_14_6_i,temp_b4_14_22_r,temp_b4_14_22_i,temp_b4_30_6_r,temp_b4_30_6_i,temp_b4_30_22_r,temp_b4_30_22_i,temp_m5_14_6_r,temp_m5_14_6_i,temp_m5_14_22_r,temp_m5_14_22_i,temp_m5_30_6_r,temp_m5_30_6_i,temp_m5_30_22_r,temp_m5_30_22_i,`W5_real,`W5_imag,`W13_real,`W13_imag,`W18_real,`W18_imag);
butterfly butterfly1238 (clk,temp_m5_14_6_r,temp_m5_14_6_i,temp_m5_14_22_r,temp_m5_14_22_i,temp_m5_30_6_r,temp_m5_30_6_i,temp_m5_30_22_r,temp_m5_30_22_i,temp_b5_14_6_r,temp_b5_14_6_i,temp_b5_14_22_r,temp_b5_14_22_i,temp_b5_30_6_r,temp_b5_30_6_i,temp_b5_30_22_r,temp_b5_30_22_i);
MULT MULT1239 (clk,temp_b4_14_7_r,temp_b4_14_7_i,temp_b4_14_23_r,temp_b4_14_23_i,temp_b4_30_7_r,temp_b4_30_7_i,temp_b4_30_23_r,temp_b4_30_23_i,temp_m5_14_7_r,temp_m5_14_7_i,temp_m5_14_23_r,temp_m5_14_23_i,temp_m5_30_7_r,temp_m5_30_7_i,temp_m5_30_23_r,temp_m5_30_23_i,`W6_real,`W6_imag,`W13_real,`W13_imag,`W19_real,`W19_imag);
butterfly butterfly1239 (clk,temp_m5_14_7_r,temp_m5_14_7_i,temp_m5_14_23_r,temp_m5_14_23_i,temp_m5_30_7_r,temp_m5_30_7_i,temp_m5_30_23_r,temp_m5_30_23_i,temp_b5_14_7_r,temp_b5_14_7_i,temp_b5_14_23_r,temp_b5_14_23_i,temp_b5_30_7_r,temp_b5_30_7_i,temp_b5_30_23_r,temp_b5_30_23_i);
MULT MULT1240 (clk,temp_b4_14_8_r,temp_b4_14_8_i,temp_b4_14_24_r,temp_b4_14_24_i,temp_b4_30_8_r,temp_b4_30_8_i,temp_b4_30_24_r,temp_b4_30_24_i,temp_m5_14_8_r,temp_m5_14_8_i,temp_m5_14_24_r,temp_m5_14_24_i,temp_m5_30_8_r,temp_m5_30_8_i,temp_m5_30_24_r,temp_m5_30_24_i,`W7_real,`W7_imag,`W13_real,`W13_imag,`W20_real,`W20_imag);
butterfly butterfly1240 (clk,temp_m5_14_8_r,temp_m5_14_8_i,temp_m5_14_24_r,temp_m5_14_24_i,temp_m5_30_8_r,temp_m5_30_8_i,temp_m5_30_24_r,temp_m5_30_24_i,temp_b5_14_8_r,temp_b5_14_8_i,temp_b5_14_24_r,temp_b5_14_24_i,temp_b5_30_8_r,temp_b5_30_8_i,temp_b5_30_24_r,temp_b5_30_24_i);
MULT MULT1241 (clk,temp_b4_14_9_r,temp_b4_14_9_i,temp_b4_14_25_r,temp_b4_14_25_i,temp_b4_30_9_r,temp_b4_30_9_i,temp_b4_30_25_r,temp_b4_30_25_i,temp_m5_14_9_r,temp_m5_14_9_i,temp_m5_14_25_r,temp_m5_14_25_i,temp_m5_30_9_r,temp_m5_30_9_i,temp_m5_30_25_r,temp_m5_30_25_i,`W8_real,`W8_imag,`W13_real,`W13_imag,`W21_real,`W21_imag);
butterfly butterfly1241 (clk,temp_m5_14_9_r,temp_m5_14_9_i,temp_m5_14_25_r,temp_m5_14_25_i,temp_m5_30_9_r,temp_m5_30_9_i,temp_m5_30_25_r,temp_m5_30_25_i,temp_b5_14_9_r,temp_b5_14_9_i,temp_b5_14_25_r,temp_b5_14_25_i,temp_b5_30_9_r,temp_b5_30_9_i,temp_b5_30_25_r,temp_b5_30_25_i);
MULT MULT1242 (clk,temp_b4_14_10_r,temp_b4_14_10_i,temp_b4_14_26_r,temp_b4_14_26_i,temp_b4_30_10_r,temp_b4_30_10_i,temp_b4_30_26_r,temp_b4_30_26_i,temp_m5_14_10_r,temp_m5_14_10_i,temp_m5_14_26_r,temp_m5_14_26_i,temp_m5_30_10_r,temp_m5_30_10_i,temp_m5_30_26_r,temp_m5_30_26_i,`W9_real,`W9_imag,`W13_real,`W13_imag,`W22_real,`W22_imag);
butterfly butterfly1242 (clk,temp_m5_14_10_r,temp_m5_14_10_i,temp_m5_14_26_r,temp_m5_14_26_i,temp_m5_30_10_r,temp_m5_30_10_i,temp_m5_30_26_r,temp_m5_30_26_i,temp_b5_14_10_r,temp_b5_14_10_i,temp_b5_14_26_r,temp_b5_14_26_i,temp_b5_30_10_r,temp_b5_30_10_i,temp_b5_30_26_r,temp_b5_30_26_i);
MULT MULT1243 (clk,temp_b4_14_11_r,temp_b4_14_11_i,temp_b4_14_27_r,temp_b4_14_27_i,temp_b4_30_11_r,temp_b4_30_11_i,temp_b4_30_27_r,temp_b4_30_27_i,temp_m5_14_11_r,temp_m5_14_11_i,temp_m5_14_27_r,temp_m5_14_27_i,temp_m5_30_11_r,temp_m5_30_11_i,temp_m5_30_27_r,temp_m5_30_27_i,`W10_real,`W10_imag,`W13_real,`W13_imag,`W23_real,`W23_imag);
butterfly butterfly1243 (clk,temp_m5_14_11_r,temp_m5_14_11_i,temp_m5_14_27_r,temp_m5_14_27_i,temp_m5_30_11_r,temp_m5_30_11_i,temp_m5_30_27_r,temp_m5_30_27_i,temp_b5_14_11_r,temp_b5_14_11_i,temp_b5_14_27_r,temp_b5_14_27_i,temp_b5_30_11_r,temp_b5_30_11_i,temp_b5_30_27_r,temp_b5_30_27_i);
MULT MULT1244 (clk,temp_b4_14_12_r,temp_b4_14_12_i,temp_b4_14_28_r,temp_b4_14_28_i,temp_b4_30_12_r,temp_b4_30_12_i,temp_b4_30_28_r,temp_b4_30_28_i,temp_m5_14_12_r,temp_m5_14_12_i,temp_m5_14_28_r,temp_m5_14_28_i,temp_m5_30_12_r,temp_m5_30_12_i,temp_m5_30_28_r,temp_m5_30_28_i,`W11_real,`W11_imag,`W13_real,`W13_imag,`W24_real,`W24_imag);
butterfly butterfly1244 (clk,temp_m5_14_12_r,temp_m5_14_12_i,temp_m5_14_28_r,temp_m5_14_28_i,temp_m5_30_12_r,temp_m5_30_12_i,temp_m5_30_28_r,temp_m5_30_28_i,temp_b5_14_12_r,temp_b5_14_12_i,temp_b5_14_28_r,temp_b5_14_28_i,temp_b5_30_12_r,temp_b5_30_12_i,temp_b5_30_28_r,temp_b5_30_28_i);
MULT MULT1245 (clk,temp_b4_14_13_r,temp_b4_14_13_i,temp_b4_14_29_r,temp_b4_14_29_i,temp_b4_30_13_r,temp_b4_30_13_i,temp_b4_30_29_r,temp_b4_30_29_i,temp_m5_14_13_r,temp_m5_14_13_i,temp_m5_14_29_r,temp_m5_14_29_i,temp_m5_30_13_r,temp_m5_30_13_i,temp_m5_30_29_r,temp_m5_30_29_i,`W12_real,`W12_imag,`W13_real,`W13_imag,`W25_real,`W25_imag);
butterfly butterfly1245 (clk,temp_m5_14_13_r,temp_m5_14_13_i,temp_m5_14_29_r,temp_m5_14_29_i,temp_m5_30_13_r,temp_m5_30_13_i,temp_m5_30_29_r,temp_m5_30_29_i,temp_b5_14_13_r,temp_b5_14_13_i,temp_b5_14_29_r,temp_b5_14_29_i,temp_b5_30_13_r,temp_b5_30_13_i,temp_b5_30_29_r,temp_b5_30_29_i);
MULT MULT1246 (clk,temp_b4_14_14_r,temp_b4_14_14_i,temp_b4_14_30_r,temp_b4_14_30_i,temp_b4_30_14_r,temp_b4_30_14_i,temp_b4_30_30_r,temp_b4_30_30_i,temp_m5_14_14_r,temp_m5_14_14_i,temp_m5_14_30_r,temp_m5_14_30_i,temp_m5_30_14_r,temp_m5_30_14_i,temp_m5_30_30_r,temp_m5_30_30_i,`W13_real,`W13_imag,`W13_real,`W13_imag,`W26_real,`W26_imag);
butterfly butterfly1246 (clk,temp_m5_14_14_r,temp_m5_14_14_i,temp_m5_14_30_r,temp_m5_14_30_i,temp_m5_30_14_r,temp_m5_30_14_i,temp_m5_30_30_r,temp_m5_30_30_i,temp_b5_14_14_r,temp_b5_14_14_i,temp_b5_14_30_r,temp_b5_14_30_i,temp_b5_30_14_r,temp_b5_30_14_i,temp_b5_30_30_r,temp_b5_30_30_i);
MULT MULT1247 (clk,temp_b4_14_15_r,temp_b4_14_15_i,temp_b4_14_31_r,temp_b4_14_31_i,temp_b4_30_15_r,temp_b4_30_15_i,temp_b4_30_31_r,temp_b4_30_31_i,temp_m5_14_15_r,temp_m5_14_15_i,temp_m5_14_31_r,temp_m5_14_31_i,temp_m5_30_15_r,temp_m5_30_15_i,temp_m5_30_31_r,temp_m5_30_31_i,`W14_real,`W14_imag,`W13_real,`W13_imag,`W27_real,`W27_imag);
butterfly butterfly1247 (clk,temp_m5_14_15_r,temp_m5_14_15_i,temp_m5_14_31_r,temp_m5_14_31_i,temp_m5_30_15_r,temp_m5_30_15_i,temp_m5_30_31_r,temp_m5_30_31_i,temp_b5_14_15_r,temp_b5_14_15_i,temp_b5_14_31_r,temp_b5_14_31_i,temp_b5_30_15_r,temp_b5_30_15_i,temp_b5_30_31_r,temp_b5_30_31_i);
MULT MULT1248 (clk,temp_b4_14_16_r,temp_b4_14_16_i,temp_b4_14_32_r,temp_b4_14_32_i,temp_b4_30_16_r,temp_b4_30_16_i,temp_b4_30_32_r,temp_b4_30_32_i,temp_m5_14_16_r,temp_m5_14_16_i,temp_m5_14_32_r,temp_m5_14_32_i,temp_m5_30_16_r,temp_m5_30_16_i,temp_m5_30_32_r,temp_m5_30_32_i,`W15_real,`W15_imag,`W13_real,`W13_imag,`W28_real,`W28_imag);
butterfly butterfly1248 (clk,temp_m5_14_16_r,temp_m5_14_16_i,temp_m5_14_32_r,temp_m5_14_32_i,temp_m5_30_16_r,temp_m5_30_16_i,temp_m5_30_32_r,temp_m5_30_32_i,temp_b5_14_16_r,temp_b5_14_16_i,temp_b5_14_32_r,temp_b5_14_32_i,temp_b5_30_16_r,temp_b5_30_16_i,temp_b5_30_32_r,temp_b5_30_32_i);
MULT MULT1249 (clk,temp_b4_15_1_r,temp_b4_15_1_i,temp_b4_15_17_r,temp_b4_15_17_i,temp_b4_31_1_r,temp_b4_31_1_i,temp_b4_31_17_r,temp_b4_31_17_i,temp_m5_15_1_r,temp_m5_15_1_i,temp_m5_15_17_r,temp_m5_15_17_i,temp_m5_31_1_r,temp_m5_31_1_i,temp_m5_31_17_r,temp_m5_31_17_i,`W0_real,`W0_imag,`W14_real,`W14_imag,`W14_real,`W14_imag);
butterfly butterfly1249 (clk,temp_m5_15_1_r,temp_m5_15_1_i,temp_m5_15_17_r,temp_m5_15_17_i,temp_m5_31_1_r,temp_m5_31_1_i,temp_m5_31_17_r,temp_m5_31_17_i,temp_b5_15_1_r,temp_b5_15_1_i,temp_b5_15_17_r,temp_b5_15_17_i,temp_b5_31_1_r,temp_b5_31_1_i,temp_b5_31_17_r,temp_b5_31_17_i);
MULT MULT1250 (clk,temp_b4_15_2_r,temp_b4_15_2_i,temp_b4_15_18_r,temp_b4_15_18_i,temp_b4_31_2_r,temp_b4_31_2_i,temp_b4_31_18_r,temp_b4_31_18_i,temp_m5_15_2_r,temp_m5_15_2_i,temp_m5_15_18_r,temp_m5_15_18_i,temp_m5_31_2_r,temp_m5_31_2_i,temp_m5_31_18_r,temp_m5_31_18_i,`W1_real,`W1_imag,`W14_real,`W14_imag,`W15_real,`W15_imag);
butterfly butterfly1250 (clk,temp_m5_15_2_r,temp_m5_15_2_i,temp_m5_15_18_r,temp_m5_15_18_i,temp_m5_31_2_r,temp_m5_31_2_i,temp_m5_31_18_r,temp_m5_31_18_i,temp_b5_15_2_r,temp_b5_15_2_i,temp_b5_15_18_r,temp_b5_15_18_i,temp_b5_31_2_r,temp_b5_31_2_i,temp_b5_31_18_r,temp_b5_31_18_i);
MULT MULT1251 (clk,temp_b4_15_3_r,temp_b4_15_3_i,temp_b4_15_19_r,temp_b4_15_19_i,temp_b4_31_3_r,temp_b4_31_3_i,temp_b4_31_19_r,temp_b4_31_19_i,temp_m5_15_3_r,temp_m5_15_3_i,temp_m5_15_19_r,temp_m5_15_19_i,temp_m5_31_3_r,temp_m5_31_3_i,temp_m5_31_19_r,temp_m5_31_19_i,`W2_real,`W2_imag,`W14_real,`W14_imag,`W16_real,`W16_imag);
butterfly butterfly1251 (clk,temp_m5_15_3_r,temp_m5_15_3_i,temp_m5_15_19_r,temp_m5_15_19_i,temp_m5_31_3_r,temp_m5_31_3_i,temp_m5_31_19_r,temp_m5_31_19_i,temp_b5_15_3_r,temp_b5_15_3_i,temp_b5_15_19_r,temp_b5_15_19_i,temp_b5_31_3_r,temp_b5_31_3_i,temp_b5_31_19_r,temp_b5_31_19_i);
MULT MULT1252 (clk,temp_b4_15_4_r,temp_b4_15_4_i,temp_b4_15_20_r,temp_b4_15_20_i,temp_b4_31_4_r,temp_b4_31_4_i,temp_b4_31_20_r,temp_b4_31_20_i,temp_m5_15_4_r,temp_m5_15_4_i,temp_m5_15_20_r,temp_m5_15_20_i,temp_m5_31_4_r,temp_m5_31_4_i,temp_m5_31_20_r,temp_m5_31_20_i,`W3_real,`W3_imag,`W14_real,`W14_imag,`W17_real,`W17_imag);
butterfly butterfly1252 (clk,temp_m5_15_4_r,temp_m5_15_4_i,temp_m5_15_20_r,temp_m5_15_20_i,temp_m5_31_4_r,temp_m5_31_4_i,temp_m5_31_20_r,temp_m5_31_20_i,temp_b5_15_4_r,temp_b5_15_4_i,temp_b5_15_20_r,temp_b5_15_20_i,temp_b5_31_4_r,temp_b5_31_4_i,temp_b5_31_20_r,temp_b5_31_20_i);
MULT MULT1253 (clk,temp_b4_15_5_r,temp_b4_15_5_i,temp_b4_15_21_r,temp_b4_15_21_i,temp_b4_31_5_r,temp_b4_31_5_i,temp_b4_31_21_r,temp_b4_31_21_i,temp_m5_15_5_r,temp_m5_15_5_i,temp_m5_15_21_r,temp_m5_15_21_i,temp_m5_31_5_r,temp_m5_31_5_i,temp_m5_31_21_r,temp_m5_31_21_i,`W4_real,`W4_imag,`W14_real,`W14_imag,`W18_real,`W18_imag);
butterfly butterfly1253 (clk,temp_m5_15_5_r,temp_m5_15_5_i,temp_m5_15_21_r,temp_m5_15_21_i,temp_m5_31_5_r,temp_m5_31_5_i,temp_m5_31_21_r,temp_m5_31_21_i,temp_b5_15_5_r,temp_b5_15_5_i,temp_b5_15_21_r,temp_b5_15_21_i,temp_b5_31_5_r,temp_b5_31_5_i,temp_b5_31_21_r,temp_b5_31_21_i);
MULT MULT1254 (clk,temp_b4_15_6_r,temp_b4_15_6_i,temp_b4_15_22_r,temp_b4_15_22_i,temp_b4_31_6_r,temp_b4_31_6_i,temp_b4_31_22_r,temp_b4_31_22_i,temp_m5_15_6_r,temp_m5_15_6_i,temp_m5_15_22_r,temp_m5_15_22_i,temp_m5_31_6_r,temp_m5_31_6_i,temp_m5_31_22_r,temp_m5_31_22_i,`W5_real,`W5_imag,`W14_real,`W14_imag,`W19_real,`W19_imag);
butterfly butterfly1254 (clk,temp_m5_15_6_r,temp_m5_15_6_i,temp_m5_15_22_r,temp_m5_15_22_i,temp_m5_31_6_r,temp_m5_31_6_i,temp_m5_31_22_r,temp_m5_31_22_i,temp_b5_15_6_r,temp_b5_15_6_i,temp_b5_15_22_r,temp_b5_15_22_i,temp_b5_31_6_r,temp_b5_31_6_i,temp_b5_31_22_r,temp_b5_31_22_i);
MULT MULT1255 (clk,temp_b4_15_7_r,temp_b4_15_7_i,temp_b4_15_23_r,temp_b4_15_23_i,temp_b4_31_7_r,temp_b4_31_7_i,temp_b4_31_23_r,temp_b4_31_23_i,temp_m5_15_7_r,temp_m5_15_7_i,temp_m5_15_23_r,temp_m5_15_23_i,temp_m5_31_7_r,temp_m5_31_7_i,temp_m5_31_23_r,temp_m5_31_23_i,`W6_real,`W6_imag,`W14_real,`W14_imag,`W20_real,`W20_imag);
butterfly butterfly1255 (clk,temp_m5_15_7_r,temp_m5_15_7_i,temp_m5_15_23_r,temp_m5_15_23_i,temp_m5_31_7_r,temp_m5_31_7_i,temp_m5_31_23_r,temp_m5_31_23_i,temp_b5_15_7_r,temp_b5_15_7_i,temp_b5_15_23_r,temp_b5_15_23_i,temp_b5_31_7_r,temp_b5_31_7_i,temp_b5_31_23_r,temp_b5_31_23_i);
MULT MULT1256 (clk,temp_b4_15_8_r,temp_b4_15_8_i,temp_b4_15_24_r,temp_b4_15_24_i,temp_b4_31_8_r,temp_b4_31_8_i,temp_b4_31_24_r,temp_b4_31_24_i,temp_m5_15_8_r,temp_m5_15_8_i,temp_m5_15_24_r,temp_m5_15_24_i,temp_m5_31_8_r,temp_m5_31_8_i,temp_m5_31_24_r,temp_m5_31_24_i,`W7_real,`W7_imag,`W14_real,`W14_imag,`W21_real,`W21_imag);
butterfly butterfly1256 (clk,temp_m5_15_8_r,temp_m5_15_8_i,temp_m5_15_24_r,temp_m5_15_24_i,temp_m5_31_8_r,temp_m5_31_8_i,temp_m5_31_24_r,temp_m5_31_24_i,temp_b5_15_8_r,temp_b5_15_8_i,temp_b5_15_24_r,temp_b5_15_24_i,temp_b5_31_8_r,temp_b5_31_8_i,temp_b5_31_24_r,temp_b5_31_24_i);
MULT MULT1257 (clk,temp_b4_15_9_r,temp_b4_15_9_i,temp_b4_15_25_r,temp_b4_15_25_i,temp_b4_31_9_r,temp_b4_31_9_i,temp_b4_31_25_r,temp_b4_31_25_i,temp_m5_15_9_r,temp_m5_15_9_i,temp_m5_15_25_r,temp_m5_15_25_i,temp_m5_31_9_r,temp_m5_31_9_i,temp_m5_31_25_r,temp_m5_31_25_i,`W8_real,`W8_imag,`W14_real,`W14_imag,`W22_real,`W22_imag);
butterfly butterfly1257 (clk,temp_m5_15_9_r,temp_m5_15_9_i,temp_m5_15_25_r,temp_m5_15_25_i,temp_m5_31_9_r,temp_m5_31_9_i,temp_m5_31_25_r,temp_m5_31_25_i,temp_b5_15_9_r,temp_b5_15_9_i,temp_b5_15_25_r,temp_b5_15_25_i,temp_b5_31_9_r,temp_b5_31_9_i,temp_b5_31_25_r,temp_b5_31_25_i);
MULT MULT1258 (clk,temp_b4_15_10_r,temp_b4_15_10_i,temp_b4_15_26_r,temp_b4_15_26_i,temp_b4_31_10_r,temp_b4_31_10_i,temp_b4_31_26_r,temp_b4_31_26_i,temp_m5_15_10_r,temp_m5_15_10_i,temp_m5_15_26_r,temp_m5_15_26_i,temp_m5_31_10_r,temp_m5_31_10_i,temp_m5_31_26_r,temp_m5_31_26_i,`W9_real,`W9_imag,`W14_real,`W14_imag,`W23_real,`W23_imag);
butterfly butterfly1258 (clk,temp_m5_15_10_r,temp_m5_15_10_i,temp_m5_15_26_r,temp_m5_15_26_i,temp_m5_31_10_r,temp_m5_31_10_i,temp_m5_31_26_r,temp_m5_31_26_i,temp_b5_15_10_r,temp_b5_15_10_i,temp_b5_15_26_r,temp_b5_15_26_i,temp_b5_31_10_r,temp_b5_31_10_i,temp_b5_31_26_r,temp_b5_31_26_i);
MULT MULT1259 (clk,temp_b4_15_11_r,temp_b4_15_11_i,temp_b4_15_27_r,temp_b4_15_27_i,temp_b4_31_11_r,temp_b4_31_11_i,temp_b4_31_27_r,temp_b4_31_27_i,temp_m5_15_11_r,temp_m5_15_11_i,temp_m5_15_27_r,temp_m5_15_27_i,temp_m5_31_11_r,temp_m5_31_11_i,temp_m5_31_27_r,temp_m5_31_27_i,`W10_real,`W10_imag,`W14_real,`W14_imag,`W24_real,`W24_imag);
butterfly butterfly1259 (clk,temp_m5_15_11_r,temp_m5_15_11_i,temp_m5_15_27_r,temp_m5_15_27_i,temp_m5_31_11_r,temp_m5_31_11_i,temp_m5_31_27_r,temp_m5_31_27_i,temp_b5_15_11_r,temp_b5_15_11_i,temp_b5_15_27_r,temp_b5_15_27_i,temp_b5_31_11_r,temp_b5_31_11_i,temp_b5_31_27_r,temp_b5_31_27_i);
MULT MULT1260 (clk,temp_b4_15_12_r,temp_b4_15_12_i,temp_b4_15_28_r,temp_b4_15_28_i,temp_b4_31_12_r,temp_b4_31_12_i,temp_b4_31_28_r,temp_b4_31_28_i,temp_m5_15_12_r,temp_m5_15_12_i,temp_m5_15_28_r,temp_m5_15_28_i,temp_m5_31_12_r,temp_m5_31_12_i,temp_m5_31_28_r,temp_m5_31_28_i,`W11_real,`W11_imag,`W14_real,`W14_imag,`W25_real,`W25_imag);
butterfly butterfly1260 (clk,temp_m5_15_12_r,temp_m5_15_12_i,temp_m5_15_28_r,temp_m5_15_28_i,temp_m5_31_12_r,temp_m5_31_12_i,temp_m5_31_28_r,temp_m5_31_28_i,temp_b5_15_12_r,temp_b5_15_12_i,temp_b5_15_28_r,temp_b5_15_28_i,temp_b5_31_12_r,temp_b5_31_12_i,temp_b5_31_28_r,temp_b5_31_28_i);
MULT MULT1261 (clk,temp_b4_15_13_r,temp_b4_15_13_i,temp_b4_15_29_r,temp_b4_15_29_i,temp_b4_31_13_r,temp_b4_31_13_i,temp_b4_31_29_r,temp_b4_31_29_i,temp_m5_15_13_r,temp_m5_15_13_i,temp_m5_15_29_r,temp_m5_15_29_i,temp_m5_31_13_r,temp_m5_31_13_i,temp_m5_31_29_r,temp_m5_31_29_i,`W12_real,`W12_imag,`W14_real,`W14_imag,`W26_real,`W26_imag);
butterfly butterfly1261 (clk,temp_m5_15_13_r,temp_m5_15_13_i,temp_m5_15_29_r,temp_m5_15_29_i,temp_m5_31_13_r,temp_m5_31_13_i,temp_m5_31_29_r,temp_m5_31_29_i,temp_b5_15_13_r,temp_b5_15_13_i,temp_b5_15_29_r,temp_b5_15_29_i,temp_b5_31_13_r,temp_b5_31_13_i,temp_b5_31_29_r,temp_b5_31_29_i);
MULT MULT1262 (clk,temp_b4_15_14_r,temp_b4_15_14_i,temp_b4_15_30_r,temp_b4_15_30_i,temp_b4_31_14_r,temp_b4_31_14_i,temp_b4_31_30_r,temp_b4_31_30_i,temp_m5_15_14_r,temp_m5_15_14_i,temp_m5_15_30_r,temp_m5_15_30_i,temp_m5_31_14_r,temp_m5_31_14_i,temp_m5_31_30_r,temp_m5_31_30_i,`W13_real,`W13_imag,`W14_real,`W14_imag,`W27_real,`W27_imag);
butterfly butterfly1262 (clk,temp_m5_15_14_r,temp_m5_15_14_i,temp_m5_15_30_r,temp_m5_15_30_i,temp_m5_31_14_r,temp_m5_31_14_i,temp_m5_31_30_r,temp_m5_31_30_i,temp_b5_15_14_r,temp_b5_15_14_i,temp_b5_15_30_r,temp_b5_15_30_i,temp_b5_31_14_r,temp_b5_31_14_i,temp_b5_31_30_r,temp_b5_31_30_i);
MULT MULT1263 (clk,temp_b4_15_15_r,temp_b4_15_15_i,temp_b4_15_31_r,temp_b4_15_31_i,temp_b4_31_15_r,temp_b4_31_15_i,temp_b4_31_31_r,temp_b4_31_31_i,temp_m5_15_15_r,temp_m5_15_15_i,temp_m5_15_31_r,temp_m5_15_31_i,temp_m5_31_15_r,temp_m5_31_15_i,temp_m5_31_31_r,temp_m5_31_31_i,`W14_real,`W14_imag,`W14_real,`W14_imag,`W28_real,`W28_imag);
butterfly butterfly1263 (clk,temp_m5_15_15_r,temp_m5_15_15_i,temp_m5_15_31_r,temp_m5_15_31_i,temp_m5_31_15_r,temp_m5_31_15_i,temp_m5_31_31_r,temp_m5_31_31_i,temp_b5_15_15_r,temp_b5_15_15_i,temp_b5_15_31_r,temp_b5_15_31_i,temp_b5_31_15_r,temp_b5_31_15_i,temp_b5_31_31_r,temp_b5_31_31_i);
MULT MULT1264 (clk,temp_b4_15_16_r,temp_b4_15_16_i,temp_b4_15_32_r,temp_b4_15_32_i,temp_b4_31_16_r,temp_b4_31_16_i,temp_b4_31_32_r,temp_b4_31_32_i,temp_m5_15_16_r,temp_m5_15_16_i,temp_m5_15_32_r,temp_m5_15_32_i,temp_m5_31_16_r,temp_m5_31_16_i,temp_m5_31_32_r,temp_m5_31_32_i,`W15_real,`W15_imag,`W14_real,`W14_imag,`W29_real,`W29_imag);
butterfly butterfly1264 (clk,temp_m5_15_16_r,temp_m5_15_16_i,temp_m5_15_32_r,temp_m5_15_32_i,temp_m5_31_16_r,temp_m5_31_16_i,temp_m5_31_32_r,temp_m5_31_32_i,temp_b5_15_16_r,temp_b5_15_16_i,temp_b5_15_32_r,temp_b5_15_32_i,temp_b5_31_16_r,temp_b5_31_16_i,temp_b5_31_32_r,temp_b5_31_32_i);
MULT MULT1265 (clk,temp_b4_16_1_r,temp_b4_16_1_i,temp_b4_16_17_r,temp_b4_16_17_i,temp_b4_32_1_r,temp_b4_32_1_i,temp_b4_32_17_r,temp_b4_32_17_i,temp_m5_16_1_r,temp_m5_16_1_i,temp_m5_16_17_r,temp_m5_16_17_i,temp_m5_32_1_r,temp_m5_32_1_i,temp_m5_32_17_r,temp_m5_32_17_i,`W0_real,`W0_imag,`W15_real,`W15_imag,`W15_real,`W15_imag);
butterfly butterfly1265 (clk,temp_m5_16_1_r,temp_m5_16_1_i,temp_m5_16_17_r,temp_m5_16_17_i,temp_m5_32_1_r,temp_m5_32_1_i,temp_m5_32_17_r,temp_m5_32_17_i,temp_b5_16_1_r,temp_b5_16_1_i,temp_b5_16_17_r,temp_b5_16_17_i,temp_b5_32_1_r,temp_b5_32_1_i,temp_b5_32_17_r,temp_b5_32_17_i);
MULT MULT1266 (clk,temp_b4_16_2_r,temp_b4_16_2_i,temp_b4_16_18_r,temp_b4_16_18_i,temp_b4_32_2_r,temp_b4_32_2_i,temp_b4_32_18_r,temp_b4_32_18_i,temp_m5_16_2_r,temp_m5_16_2_i,temp_m5_16_18_r,temp_m5_16_18_i,temp_m5_32_2_r,temp_m5_32_2_i,temp_m5_32_18_r,temp_m5_32_18_i,`W1_real,`W1_imag,`W15_real,`W15_imag,`W16_real,`W16_imag);
butterfly butterfly1266 (clk,temp_m5_16_2_r,temp_m5_16_2_i,temp_m5_16_18_r,temp_m5_16_18_i,temp_m5_32_2_r,temp_m5_32_2_i,temp_m5_32_18_r,temp_m5_32_18_i,temp_b5_16_2_r,temp_b5_16_2_i,temp_b5_16_18_r,temp_b5_16_18_i,temp_b5_32_2_r,temp_b5_32_2_i,temp_b5_32_18_r,temp_b5_32_18_i);
MULT MULT1267 (clk,temp_b4_16_3_r,temp_b4_16_3_i,temp_b4_16_19_r,temp_b4_16_19_i,temp_b4_32_3_r,temp_b4_32_3_i,temp_b4_32_19_r,temp_b4_32_19_i,temp_m5_16_3_r,temp_m5_16_3_i,temp_m5_16_19_r,temp_m5_16_19_i,temp_m5_32_3_r,temp_m5_32_3_i,temp_m5_32_19_r,temp_m5_32_19_i,`W2_real,`W2_imag,`W15_real,`W15_imag,`W17_real,`W17_imag);
butterfly butterfly1267 (clk,temp_m5_16_3_r,temp_m5_16_3_i,temp_m5_16_19_r,temp_m5_16_19_i,temp_m5_32_3_r,temp_m5_32_3_i,temp_m5_32_19_r,temp_m5_32_19_i,temp_b5_16_3_r,temp_b5_16_3_i,temp_b5_16_19_r,temp_b5_16_19_i,temp_b5_32_3_r,temp_b5_32_3_i,temp_b5_32_19_r,temp_b5_32_19_i);
MULT MULT1268 (clk,temp_b4_16_4_r,temp_b4_16_4_i,temp_b4_16_20_r,temp_b4_16_20_i,temp_b4_32_4_r,temp_b4_32_4_i,temp_b4_32_20_r,temp_b4_32_20_i,temp_m5_16_4_r,temp_m5_16_4_i,temp_m5_16_20_r,temp_m5_16_20_i,temp_m5_32_4_r,temp_m5_32_4_i,temp_m5_32_20_r,temp_m5_32_20_i,`W3_real,`W3_imag,`W15_real,`W15_imag,`W18_real,`W18_imag);
butterfly butterfly1268 (clk,temp_m5_16_4_r,temp_m5_16_4_i,temp_m5_16_20_r,temp_m5_16_20_i,temp_m5_32_4_r,temp_m5_32_4_i,temp_m5_32_20_r,temp_m5_32_20_i,temp_b5_16_4_r,temp_b5_16_4_i,temp_b5_16_20_r,temp_b5_16_20_i,temp_b5_32_4_r,temp_b5_32_4_i,temp_b5_32_20_r,temp_b5_32_20_i);
MULT MULT1269 (clk,temp_b4_16_5_r,temp_b4_16_5_i,temp_b4_16_21_r,temp_b4_16_21_i,temp_b4_32_5_r,temp_b4_32_5_i,temp_b4_32_21_r,temp_b4_32_21_i,temp_m5_16_5_r,temp_m5_16_5_i,temp_m5_16_21_r,temp_m5_16_21_i,temp_m5_32_5_r,temp_m5_32_5_i,temp_m5_32_21_r,temp_m5_32_21_i,`W4_real,`W4_imag,`W15_real,`W15_imag,`W19_real,`W19_imag);
butterfly butterfly1269 (clk,temp_m5_16_5_r,temp_m5_16_5_i,temp_m5_16_21_r,temp_m5_16_21_i,temp_m5_32_5_r,temp_m5_32_5_i,temp_m5_32_21_r,temp_m5_32_21_i,temp_b5_16_5_r,temp_b5_16_5_i,temp_b5_16_21_r,temp_b5_16_21_i,temp_b5_32_5_r,temp_b5_32_5_i,temp_b5_32_21_r,temp_b5_32_21_i);
MULT MULT1270 (clk,temp_b4_16_6_r,temp_b4_16_6_i,temp_b4_16_22_r,temp_b4_16_22_i,temp_b4_32_6_r,temp_b4_32_6_i,temp_b4_32_22_r,temp_b4_32_22_i,temp_m5_16_6_r,temp_m5_16_6_i,temp_m5_16_22_r,temp_m5_16_22_i,temp_m5_32_6_r,temp_m5_32_6_i,temp_m5_32_22_r,temp_m5_32_22_i,`W5_real,`W5_imag,`W15_real,`W15_imag,`W20_real,`W20_imag);
butterfly butterfly1270 (clk,temp_m5_16_6_r,temp_m5_16_6_i,temp_m5_16_22_r,temp_m5_16_22_i,temp_m5_32_6_r,temp_m5_32_6_i,temp_m5_32_22_r,temp_m5_32_22_i,temp_b5_16_6_r,temp_b5_16_6_i,temp_b5_16_22_r,temp_b5_16_22_i,temp_b5_32_6_r,temp_b5_32_6_i,temp_b5_32_22_r,temp_b5_32_22_i);
MULT MULT1271 (clk,temp_b4_16_7_r,temp_b4_16_7_i,temp_b4_16_23_r,temp_b4_16_23_i,temp_b4_32_7_r,temp_b4_32_7_i,temp_b4_32_23_r,temp_b4_32_23_i,temp_m5_16_7_r,temp_m5_16_7_i,temp_m5_16_23_r,temp_m5_16_23_i,temp_m5_32_7_r,temp_m5_32_7_i,temp_m5_32_23_r,temp_m5_32_23_i,`W6_real,`W6_imag,`W15_real,`W15_imag,`W21_real,`W21_imag);
butterfly butterfly1271 (clk,temp_m5_16_7_r,temp_m5_16_7_i,temp_m5_16_23_r,temp_m5_16_23_i,temp_m5_32_7_r,temp_m5_32_7_i,temp_m5_32_23_r,temp_m5_32_23_i,temp_b5_16_7_r,temp_b5_16_7_i,temp_b5_16_23_r,temp_b5_16_23_i,temp_b5_32_7_r,temp_b5_32_7_i,temp_b5_32_23_r,temp_b5_32_23_i);
MULT MULT1272 (clk,temp_b4_16_8_r,temp_b4_16_8_i,temp_b4_16_24_r,temp_b4_16_24_i,temp_b4_32_8_r,temp_b4_32_8_i,temp_b4_32_24_r,temp_b4_32_24_i,temp_m5_16_8_r,temp_m5_16_8_i,temp_m5_16_24_r,temp_m5_16_24_i,temp_m5_32_8_r,temp_m5_32_8_i,temp_m5_32_24_r,temp_m5_32_24_i,`W7_real,`W7_imag,`W15_real,`W15_imag,`W22_real,`W22_imag);
butterfly butterfly1272 (clk,temp_m5_16_8_r,temp_m5_16_8_i,temp_m5_16_24_r,temp_m5_16_24_i,temp_m5_32_8_r,temp_m5_32_8_i,temp_m5_32_24_r,temp_m5_32_24_i,temp_b5_16_8_r,temp_b5_16_8_i,temp_b5_16_24_r,temp_b5_16_24_i,temp_b5_32_8_r,temp_b5_32_8_i,temp_b5_32_24_r,temp_b5_32_24_i);
MULT MULT1273 (clk,temp_b4_16_9_r,temp_b4_16_9_i,temp_b4_16_25_r,temp_b4_16_25_i,temp_b4_32_9_r,temp_b4_32_9_i,temp_b4_32_25_r,temp_b4_32_25_i,temp_m5_16_9_r,temp_m5_16_9_i,temp_m5_16_25_r,temp_m5_16_25_i,temp_m5_32_9_r,temp_m5_32_9_i,temp_m5_32_25_r,temp_m5_32_25_i,`W8_real,`W8_imag,`W15_real,`W15_imag,`W23_real,`W23_imag);
butterfly butterfly1273 (clk,temp_m5_16_9_r,temp_m5_16_9_i,temp_m5_16_25_r,temp_m5_16_25_i,temp_m5_32_9_r,temp_m5_32_9_i,temp_m5_32_25_r,temp_m5_32_25_i,temp_b5_16_9_r,temp_b5_16_9_i,temp_b5_16_25_r,temp_b5_16_25_i,temp_b5_32_9_r,temp_b5_32_9_i,temp_b5_32_25_r,temp_b5_32_25_i);
MULT MULT1274 (clk,temp_b4_16_10_r,temp_b4_16_10_i,temp_b4_16_26_r,temp_b4_16_26_i,temp_b4_32_10_r,temp_b4_32_10_i,temp_b4_32_26_r,temp_b4_32_26_i,temp_m5_16_10_r,temp_m5_16_10_i,temp_m5_16_26_r,temp_m5_16_26_i,temp_m5_32_10_r,temp_m5_32_10_i,temp_m5_32_26_r,temp_m5_32_26_i,`W9_real,`W9_imag,`W15_real,`W15_imag,`W24_real,`W24_imag);
butterfly butterfly1274 (clk,temp_m5_16_10_r,temp_m5_16_10_i,temp_m5_16_26_r,temp_m5_16_26_i,temp_m5_32_10_r,temp_m5_32_10_i,temp_m5_32_26_r,temp_m5_32_26_i,temp_b5_16_10_r,temp_b5_16_10_i,temp_b5_16_26_r,temp_b5_16_26_i,temp_b5_32_10_r,temp_b5_32_10_i,temp_b5_32_26_r,temp_b5_32_26_i);
MULT MULT1275 (clk,temp_b4_16_11_r,temp_b4_16_11_i,temp_b4_16_27_r,temp_b4_16_27_i,temp_b4_32_11_r,temp_b4_32_11_i,temp_b4_32_27_r,temp_b4_32_27_i,temp_m5_16_11_r,temp_m5_16_11_i,temp_m5_16_27_r,temp_m5_16_27_i,temp_m5_32_11_r,temp_m5_32_11_i,temp_m5_32_27_r,temp_m5_32_27_i,`W10_real,`W10_imag,`W15_real,`W15_imag,`W25_real,`W25_imag);
butterfly butterfly1275 (clk,temp_m5_16_11_r,temp_m5_16_11_i,temp_m5_16_27_r,temp_m5_16_27_i,temp_m5_32_11_r,temp_m5_32_11_i,temp_m5_32_27_r,temp_m5_32_27_i,temp_b5_16_11_r,temp_b5_16_11_i,temp_b5_16_27_r,temp_b5_16_27_i,temp_b5_32_11_r,temp_b5_32_11_i,temp_b5_32_27_r,temp_b5_32_27_i);
MULT MULT1276 (clk,temp_b4_16_12_r,temp_b4_16_12_i,temp_b4_16_28_r,temp_b4_16_28_i,temp_b4_32_12_r,temp_b4_32_12_i,temp_b4_32_28_r,temp_b4_32_28_i,temp_m5_16_12_r,temp_m5_16_12_i,temp_m5_16_28_r,temp_m5_16_28_i,temp_m5_32_12_r,temp_m5_32_12_i,temp_m5_32_28_r,temp_m5_32_28_i,`W11_real,`W11_imag,`W15_real,`W15_imag,`W26_real,`W26_imag);
butterfly butterfly1276 (clk,temp_m5_16_12_r,temp_m5_16_12_i,temp_m5_16_28_r,temp_m5_16_28_i,temp_m5_32_12_r,temp_m5_32_12_i,temp_m5_32_28_r,temp_m5_32_28_i,temp_b5_16_12_r,temp_b5_16_12_i,temp_b5_16_28_r,temp_b5_16_28_i,temp_b5_32_12_r,temp_b5_32_12_i,temp_b5_32_28_r,temp_b5_32_28_i);
MULT MULT1277 (clk,temp_b4_16_13_r,temp_b4_16_13_i,temp_b4_16_29_r,temp_b4_16_29_i,temp_b4_32_13_r,temp_b4_32_13_i,temp_b4_32_29_r,temp_b4_32_29_i,temp_m5_16_13_r,temp_m5_16_13_i,temp_m5_16_29_r,temp_m5_16_29_i,temp_m5_32_13_r,temp_m5_32_13_i,temp_m5_32_29_r,temp_m5_32_29_i,`W12_real,`W12_imag,`W15_real,`W15_imag,`W27_real,`W27_imag);
butterfly butterfly1277 (clk,temp_m5_16_13_r,temp_m5_16_13_i,temp_m5_16_29_r,temp_m5_16_29_i,temp_m5_32_13_r,temp_m5_32_13_i,temp_m5_32_29_r,temp_m5_32_29_i,temp_b5_16_13_r,temp_b5_16_13_i,temp_b5_16_29_r,temp_b5_16_29_i,temp_b5_32_13_r,temp_b5_32_13_i,temp_b5_32_29_r,temp_b5_32_29_i);
MULT MULT1278 (clk,temp_b4_16_14_r,temp_b4_16_14_i,temp_b4_16_30_r,temp_b4_16_30_i,temp_b4_32_14_r,temp_b4_32_14_i,temp_b4_32_30_r,temp_b4_32_30_i,temp_m5_16_14_r,temp_m5_16_14_i,temp_m5_16_30_r,temp_m5_16_30_i,temp_m5_32_14_r,temp_m5_32_14_i,temp_m5_32_30_r,temp_m5_32_30_i,`W13_real,`W13_imag,`W15_real,`W15_imag,`W28_real,`W28_imag);
butterfly butterfly1278 (clk,temp_m5_16_14_r,temp_m5_16_14_i,temp_m5_16_30_r,temp_m5_16_30_i,temp_m5_32_14_r,temp_m5_32_14_i,temp_m5_32_30_r,temp_m5_32_30_i,temp_b5_16_14_r,temp_b5_16_14_i,temp_b5_16_30_r,temp_b5_16_30_i,temp_b5_32_14_r,temp_b5_32_14_i,temp_b5_32_30_r,temp_b5_32_30_i);
MULT MULT1279 (clk,temp_b4_16_15_r,temp_b4_16_15_i,temp_b4_16_31_r,temp_b4_16_31_i,temp_b4_32_15_r,temp_b4_32_15_i,temp_b4_32_31_r,temp_b4_32_31_i,temp_m5_16_15_r,temp_m5_16_15_i,temp_m5_16_31_r,temp_m5_16_31_i,temp_m5_32_15_r,temp_m5_32_15_i,temp_m5_32_31_r,temp_m5_32_31_i,`W14_real,`W14_imag,`W15_real,`W15_imag,`W29_real,`W29_imag);
butterfly butterfly1279 (clk,temp_m5_16_15_r,temp_m5_16_15_i,temp_m5_16_31_r,temp_m5_16_31_i,temp_m5_32_15_r,temp_m5_32_15_i,temp_m5_32_31_r,temp_m5_32_31_i,temp_b5_16_15_r,temp_b5_16_15_i,temp_b5_16_31_r,temp_b5_16_31_i,temp_b5_32_15_r,temp_b5_32_15_i,temp_b5_32_31_r,temp_b5_32_31_i);
MULT MULT1280 (clk,temp_b4_16_16_r,temp_b4_16_16_i,temp_b4_16_32_r,temp_b4_16_32_i,temp_b4_32_16_r,temp_b4_32_16_i,temp_b4_32_32_r,temp_b4_32_32_i,temp_m5_16_16_r,temp_m5_16_16_i,temp_m5_16_32_r,temp_m5_16_32_i,temp_m5_32_16_r,temp_m5_32_16_i,temp_m5_32_32_r,temp_m5_32_32_i,`W15_real,`W15_imag,`W15_real,`W15_imag,`W30_real,`W30_imag);
butterfly butterfly1280 (clk,temp_m5_16_16_r,temp_m5_16_16_i,temp_m5_16_32_r,temp_m5_16_32_i,temp_m5_32_16_r,temp_m5_32_16_i,temp_m5_32_32_r,temp_m5_32_32_i,temp_b5_16_16_r,temp_b5_16_16_i,temp_b5_16_32_r,temp_b5_16_32_i,temp_b5_32_16_r,temp_b5_32_16_i,temp_b5_32_32_r,temp_b5_32_32_i);

/******************in out assgin*******************/

assign in_1_1_r = in_r;
assign in_1_1_i = in_i;
assign in_1_2_r = in_r;
assign in_1_2_i = in_i;
assign in_1_3_r = in_r;
assign in_1_3_i = in_i;
assign in_1_4_r = in_r;
assign in_1_4_i = in_i;
assign in_1_5_r = in_r;
assign in_1_5_i = in_i;
assign in_1_6_r = in_r;
assign in_1_6_i = in_i;
assign in_1_7_r = in_r;
assign in_1_7_i = in_i;
assign in_1_8_r = in_r;
assign in_1_8_i = in_i;
assign in_1_9_r = in_r;
assign in_1_9_i = in_i;
assign in_1_10_r = in_r;
assign in_1_10_i = in_i;
assign in_1_11_r = in_r;
assign in_1_11_i = in_i;
assign in_1_12_r = in_r;
assign in_1_12_i = in_i;
assign in_1_13_r = in_r;
assign in_1_13_i = in_i;
assign in_1_14_r = in_r;
assign in_1_14_i = in_i;
assign in_1_15_r = in_r;
assign in_1_15_i = in_i;
assign in_1_16_r = in_r;
assign in_1_16_i = in_i;
assign in_1_17_r = in_r;
assign in_1_17_i = in_i;
assign in_1_18_r = in_r;
assign in_1_18_i = in_i;
assign in_1_19_r = in_r;
assign in_1_19_i = in_i;
assign in_1_20_r = in_r;
assign in_1_20_i = in_i;
assign in_1_21_r = in_r;
assign in_1_21_i = in_i;
assign in_1_22_r = in_r;
assign in_1_22_i = in_i;
assign in_1_23_r = in_r;
assign in_1_23_i = in_i;
assign in_1_24_r = in_r;
assign in_1_24_i = in_i;
assign in_1_25_r = in_r;
assign in_1_25_i = in_i;
assign in_1_26_r = in_r;
assign in_1_26_i = in_i;
assign in_1_27_r = in_r;
assign in_1_27_i = in_i;
assign in_1_28_r = in_r;
assign in_1_28_i = in_i;
assign in_1_29_r = in_r;
assign in_1_29_i = in_i;
assign in_1_30_r = in_r;
assign in_1_30_i = in_i;
assign in_1_31_r = in_r;
assign in_1_31_i = in_i;
assign in_1_32_r = in_r;
assign in_1_32_i = in_i;
assign in_2_1_r = in_r;
assign in_2_1_i = in_i;
assign in_2_2_r = in_r;
assign in_2_2_i = in_i;
assign in_2_3_r = in_r;
assign in_2_3_i = in_i;
assign in_2_4_r = in_r;
assign in_2_4_i = in_i;
assign in_2_5_r = in_r;
assign in_2_5_i = in_i;
assign in_2_6_r = in_r;
assign in_2_6_i = in_i;
assign in_2_7_r = in_r;
assign in_2_7_i = in_i;
assign in_2_8_r = in_r;
assign in_2_8_i = in_i;
assign in_2_9_r = in_r;
assign in_2_9_i = in_i;
assign in_2_10_r = in_r;
assign in_2_10_i = in_i;
assign in_2_11_r = in_r;
assign in_2_11_i = in_i;
assign in_2_12_r = in_r;
assign in_2_12_i = in_i;
assign in_2_13_r = in_r;
assign in_2_13_i = in_i;
assign in_2_14_r = in_r;
assign in_2_14_i = in_i;
assign in_2_15_r = in_r;
assign in_2_15_i = in_i;
assign in_2_16_r = in_r;
assign in_2_16_i = in_i;
assign in_2_17_r = in_r;
assign in_2_17_i = in_i;
assign in_2_18_r = in_r;
assign in_2_18_i = in_i;
assign in_2_19_r = in_r;
assign in_2_19_i = in_i;
assign in_2_20_r = in_r;
assign in_2_20_i = in_i;
assign in_2_21_r = in_r;
assign in_2_21_i = in_i;
assign in_2_22_r = in_r;
assign in_2_22_i = in_i;
assign in_2_23_r = in_r;
assign in_2_23_i = in_i;
assign in_2_24_r = in_r;
assign in_2_24_i = in_i;
assign in_2_25_r = in_r;
assign in_2_25_i = in_i;
assign in_2_26_r = in_r;
assign in_2_26_i = in_i;
assign in_2_27_r = in_r;
assign in_2_27_i = in_i;
assign in_2_28_r = in_r;
assign in_2_28_i = in_i;
assign in_2_29_r = in_r;
assign in_2_29_i = in_i;
assign in_2_30_r = in_r;
assign in_2_30_i = in_i;
assign in_2_31_r = in_r;
assign in_2_31_i = in_i;
assign in_2_32_r = in_r;
assign in_2_32_i = in_i;
assign in_3_1_r = in_r;
assign in_3_1_i = in_i;
assign in_3_2_r = in_r;
assign in_3_2_i = in_i;
assign in_3_3_r = in_r;
assign in_3_3_i = in_i;
assign in_3_4_r = in_r;
assign in_3_4_i = in_i;
assign in_3_5_r = in_r;
assign in_3_5_i = in_i;
assign in_3_6_r = in_r;
assign in_3_6_i = in_i;
assign in_3_7_r = in_r;
assign in_3_7_i = in_i;
assign in_3_8_r = in_r;
assign in_3_8_i = in_i;
assign in_3_9_r = in_r;
assign in_3_9_i = in_i;
assign in_3_10_r = in_r;
assign in_3_10_i = in_i;
assign in_3_11_r = in_r;
assign in_3_11_i = in_i;
assign in_3_12_r = in_r;
assign in_3_12_i = in_i;
assign in_3_13_r = in_r;
assign in_3_13_i = in_i;
assign in_3_14_r = in_r;
assign in_3_14_i = in_i;
assign in_3_15_r = in_r;
assign in_3_15_i = in_i;
assign in_3_16_r = in_r;
assign in_3_16_i = in_i;
assign in_3_17_r = in_r;
assign in_3_17_i = in_i;
assign in_3_18_r = in_r;
assign in_3_18_i = in_i;
assign in_3_19_r = in_r;
assign in_3_19_i = in_i;
assign in_3_20_r = in_r;
assign in_3_20_i = in_i;
assign in_3_21_r = in_r;
assign in_3_21_i = in_i;
assign in_3_22_r = in_r;
assign in_3_22_i = in_i;
assign in_3_23_r = in_r;
assign in_3_23_i = in_i;
assign in_3_24_r = in_r;
assign in_3_24_i = in_i;
assign in_3_25_r = in_r;
assign in_3_25_i = in_i;
assign in_3_26_r = in_r;
assign in_3_26_i = in_i;
assign in_3_27_r = in_r;
assign in_3_27_i = in_i;
assign in_3_28_r = in_r;
assign in_3_28_i = in_i;
assign in_3_29_r = in_r;
assign in_3_29_i = in_i;
assign in_3_30_r = in_r;
assign in_3_30_i = in_i;
assign in_3_31_r = in_r;
assign in_3_31_i = in_i;
assign in_3_32_r = in_r;
assign in_3_32_i = in_i;
assign in_4_1_r = in_r;
assign in_4_1_i = in_i;
assign in_4_2_r = in_r;
assign in_4_2_i = in_i;
assign in_4_3_r = in_r;
assign in_4_3_i = in_i;
assign in_4_4_r = in_r;
assign in_4_4_i = in_i;
assign in_4_5_r = in_r;
assign in_4_5_i = in_i;
assign in_4_6_r = in_r;
assign in_4_6_i = in_i;
assign in_4_7_r = in_r;
assign in_4_7_i = in_i;
assign in_4_8_r = in_r;
assign in_4_8_i = in_i;
assign in_4_9_r = in_r;
assign in_4_9_i = in_i;
assign in_4_10_r = in_r;
assign in_4_10_i = in_i;
assign in_4_11_r = in_r;
assign in_4_11_i = in_i;
assign in_4_12_r = in_r;
assign in_4_12_i = in_i;
assign in_4_13_r = in_r;
assign in_4_13_i = in_i;
assign in_4_14_r = in_r;
assign in_4_14_i = in_i;
assign in_4_15_r = in_r;
assign in_4_15_i = in_i;
assign in_4_16_r = in_r;
assign in_4_16_i = in_i;
assign in_4_17_r = in_r;
assign in_4_17_i = in_i;
assign in_4_18_r = in_r;
assign in_4_18_i = in_i;
assign in_4_19_r = in_r;
assign in_4_19_i = in_i;
assign in_4_20_r = in_r;
assign in_4_20_i = in_i;
assign in_4_21_r = in_r;
assign in_4_21_i = in_i;
assign in_4_22_r = in_r;
assign in_4_22_i = in_i;
assign in_4_23_r = in_r;
assign in_4_23_i = in_i;
assign in_4_24_r = in_r;
assign in_4_24_i = in_i;
assign in_4_25_r = in_r;
assign in_4_25_i = in_i;
assign in_4_26_r = in_r;
assign in_4_26_i = in_i;
assign in_4_27_r = in_r;
assign in_4_27_i = in_i;
assign in_4_28_r = in_r;
assign in_4_28_i = in_i;
assign in_4_29_r = in_r;
assign in_4_29_i = in_i;
assign in_4_30_r = in_r;
assign in_4_30_i = in_i;
assign in_4_31_r = in_r;
assign in_4_31_i = in_i;
assign in_4_32_r = in_r;
assign in_4_32_i = in_i;
assign in_5_1_r = in_r;
assign in_5_1_i = in_i;
assign in_5_2_r = in_r;
assign in_5_2_i = in_i;
assign in_5_3_r = in_r;
assign in_5_3_i = in_i;
assign in_5_4_r = in_r;
assign in_5_4_i = in_i;
assign in_5_5_r = in_r;
assign in_5_5_i = in_i;
assign in_5_6_r = in_r;
assign in_5_6_i = in_i;
assign in_5_7_r = in_r;
assign in_5_7_i = in_i;
assign in_5_8_r = in_r;
assign in_5_8_i = in_i;
assign in_5_9_r = in_r;
assign in_5_9_i = in_i;
assign in_5_10_r = in_r;
assign in_5_10_i = in_i;
assign in_5_11_r = in_r;
assign in_5_11_i = in_i;
assign in_5_12_r = in_r;
assign in_5_12_i = in_i;
assign in_5_13_r = in_r;
assign in_5_13_i = in_i;
assign in_5_14_r = in_r;
assign in_5_14_i = in_i;
assign in_5_15_r = in_r;
assign in_5_15_i = in_i;
assign in_5_16_r = in_r;
assign in_5_16_i = in_i;
assign in_5_17_r = in_r;
assign in_5_17_i = in_i;
assign in_5_18_r = in_r;
assign in_5_18_i = in_i;
assign in_5_19_r = in_r;
assign in_5_19_i = in_i;
assign in_5_20_r = in_r;
assign in_5_20_i = in_i;
assign in_5_21_r = in_r;
assign in_5_21_i = in_i;
assign in_5_22_r = in_r;
assign in_5_22_i = in_i;
assign in_5_23_r = in_r;
assign in_5_23_i = in_i;
assign in_5_24_r = in_r;
assign in_5_24_i = in_i;
assign in_5_25_r = in_r;
assign in_5_25_i = in_i;
assign in_5_26_r = in_r;
assign in_5_26_i = in_i;
assign in_5_27_r = in_r;
assign in_5_27_i = in_i;
assign in_5_28_r = in_r;
assign in_5_28_i = in_i;
assign in_5_29_r = in_r;
assign in_5_29_i = in_i;
assign in_5_30_r = in_r;
assign in_5_30_i = in_i;
assign in_5_31_r = in_r;
assign in_5_31_i = in_i;
assign in_5_32_r = in_r;
assign in_5_32_i = in_i;
assign in_6_1_r = in_r;
assign in_6_1_i = in_i;
assign in_6_2_r = in_r;
assign in_6_2_i = in_i;
assign in_6_3_r = in_r;
assign in_6_3_i = in_i;
assign in_6_4_r = in_r;
assign in_6_4_i = in_i;
assign in_6_5_r = in_r;
assign in_6_5_i = in_i;
assign in_6_6_r = in_r;
assign in_6_6_i = in_i;
assign in_6_7_r = in_r;
assign in_6_7_i = in_i;
assign in_6_8_r = in_r;
assign in_6_8_i = in_i;
assign in_6_9_r = in_r;
assign in_6_9_i = in_i;
assign in_6_10_r = in_r;
assign in_6_10_i = in_i;
assign in_6_11_r = in_r;
assign in_6_11_i = in_i;
assign in_6_12_r = in_r;
assign in_6_12_i = in_i;
assign in_6_13_r = in_r;
assign in_6_13_i = in_i;
assign in_6_14_r = in_r;
assign in_6_14_i = in_i;
assign in_6_15_r = in_r;
assign in_6_15_i = in_i;
assign in_6_16_r = in_r;
assign in_6_16_i = in_i;
assign in_6_17_r = in_r;
assign in_6_17_i = in_i;
assign in_6_18_r = in_r;
assign in_6_18_i = in_i;
assign in_6_19_r = in_r;
assign in_6_19_i = in_i;
assign in_6_20_r = in_r;
assign in_6_20_i = in_i;
assign in_6_21_r = in_r;
assign in_6_21_i = in_i;
assign in_6_22_r = in_r;
assign in_6_22_i = in_i;
assign in_6_23_r = in_r;
assign in_6_23_i = in_i;
assign in_6_24_r = in_r;
assign in_6_24_i = in_i;
assign in_6_25_r = in_r;
assign in_6_25_i = in_i;
assign in_6_26_r = in_r;
assign in_6_26_i = in_i;
assign in_6_27_r = in_r;
assign in_6_27_i = in_i;
assign in_6_28_r = in_r;
assign in_6_28_i = in_i;
assign in_6_29_r = in_r;
assign in_6_29_i = in_i;
assign in_6_30_r = in_r;
assign in_6_30_i = in_i;
assign in_6_31_r = in_r;
assign in_6_31_i = in_i;
assign in_6_32_r = in_r;
assign in_6_32_i = in_i;
assign in_7_1_r = in_r;
assign in_7_1_i = in_i;
assign in_7_2_r = in_r;
assign in_7_2_i = in_i;
assign in_7_3_r = in_r;
assign in_7_3_i = in_i;
assign in_7_4_r = in_r;
assign in_7_4_i = in_i;
assign in_7_5_r = in_r;
assign in_7_5_i = in_i;
assign in_7_6_r = in_r;
assign in_7_6_i = in_i;
assign in_7_7_r = in_r;
assign in_7_7_i = in_i;
assign in_7_8_r = in_r;
assign in_7_8_i = in_i;
assign in_7_9_r = in_r;
assign in_7_9_i = in_i;
assign in_7_10_r = in_r;
assign in_7_10_i = in_i;
assign in_7_11_r = in_r;
assign in_7_11_i = in_i;
assign in_7_12_r = in_r;
assign in_7_12_i = in_i;
assign in_7_13_r = in_r;
assign in_7_13_i = in_i;
assign in_7_14_r = in_r;
assign in_7_14_i = in_i;
assign in_7_15_r = in_r;
assign in_7_15_i = in_i;
assign in_7_16_r = in_r;
assign in_7_16_i = in_i;
assign in_7_17_r = in_r;
assign in_7_17_i = in_i;
assign in_7_18_r = in_r;
assign in_7_18_i = in_i;
assign in_7_19_r = in_r;
assign in_7_19_i = in_i;
assign in_7_20_r = in_r;
assign in_7_20_i = in_i;
assign in_7_21_r = in_r;
assign in_7_21_i = in_i;
assign in_7_22_r = in_r;
assign in_7_22_i = in_i;
assign in_7_23_r = in_r;
assign in_7_23_i = in_i;
assign in_7_24_r = in_r;
assign in_7_24_i = in_i;
assign in_7_25_r = in_r;
assign in_7_25_i = in_i;
assign in_7_26_r = in_r;
assign in_7_26_i = in_i;
assign in_7_27_r = in_r;
assign in_7_27_i = in_i;
assign in_7_28_r = in_r;
assign in_7_28_i = in_i;
assign in_7_29_r = in_r;
assign in_7_29_i = in_i;
assign in_7_30_r = in_r;
assign in_7_30_i = in_i;
assign in_7_31_r = in_r;
assign in_7_31_i = in_i;
assign in_7_32_r = in_r;
assign in_7_32_i = in_i;
assign in_8_1_r = in_r;
assign in_8_1_i = in_i;
assign in_8_2_r = in_r;
assign in_8_2_i = in_i;
assign in_8_3_r = in_r;
assign in_8_3_i = in_i;
assign in_8_4_r = in_r;
assign in_8_4_i = in_i;
assign in_8_5_r = in_r;
assign in_8_5_i = in_i;
assign in_8_6_r = in_r;
assign in_8_6_i = in_i;
assign in_8_7_r = in_r;
assign in_8_7_i = in_i;
assign in_8_8_r = in_r;
assign in_8_8_i = in_i;
assign in_8_9_r = in_r;
assign in_8_9_i = in_i;
assign in_8_10_r = in_r;
assign in_8_10_i = in_i;
assign in_8_11_r = in_r;
assign in_8_11_i = in_i;
assign in_8_12_r = in_r;
assign in_8_12_i = in_i;
assign in_8_13_r = in_r;
assign in_8_13_i = in_i;
assign in_8_14_r = in_r;
assign in_8_14_i = in_i;
assign in_8_15_r = in_r;
assign in_8_15_i = in_i;
assign in_8_16_r = in_r;
assign in_8_16_i = in_i;
assign in_8_17_r = in_r;
assign in_8_17_i = in_i;
assign in_8_18_r = in_r;
assign in_8_18_i = in_i;
assign in_8_19_r = in_r;
assign in_8_19_i = in_i;
assign in_8_20_r = in_r;
assign in_8_20_i = in_i;
assign in_8_21_r = in_r;
assign in_8_21_i = in_i;
assign in_8_22_r = in_r;
assign in_8_22_i = in_i;
assign in_8_23_r = in_r;
assign in_8_23_i = in_i;
assign in_8_24_r = in_r;
assign in_8_24_i = in_i;
assign in_8_25_r = in_r;
assign in_8_25_i = in_i;
assign in_8_26_r = in_r;
assign in_8_26_i = in_i;
assign in_8_27_r = in_r;
assign in_8_27_i = in_i;
assign in_8_28_r = in_r;
assign in_8_28_i = in_i;
assign in_8_29_r = in_r;
assign in_8_29_i = in_i;
assign in_8_30_r = in_r;
assign in_8_30_i = in_i;
assign in_8_31_r = in_r;
assign in_8_31_i = in_i;
assign in_8_32_r = in_r;
assign in_8_32_i = in_i;
assign in_9_1_r = in_r;
assign in_9_1_i = in_i;
assign in_9_2_r = in_r;
assign in_9_2_i = in_i;
assign in_9_3_r = in_r;
assign in_9_3_i = in_i;
assign in_9_4_r = in_r;
assign in_9_4_i = in_i;
assign in_9_5_r = in_r;
assign in_9_5_i = in_i;
assign in_9_6_r = in_r;
assign in_9_6_i = in_i;
assign in_9_7_r = in_r;
assign in_9_7_i = in_i;
assign in_9_8_r = in_r;
assign in_9_8_i = in_i;
assign in_9_9_r = in_r;
assign in_9_9_i = in_i;
assign in_9_10_r = in_r;
assign in_9_10_i = in_i;
assign in_9_11_r = in_r;
assign in_9_11_i = in_i;
assign in_9_12_r = in_r;
assign in_9_12_i = in_i;
assign in_9_13_r = in_r;
assign in_9_13_i = in_i;
assign in_9_14_r = in_r;
assign in_9_14_i = in_i;
assign in_9_15_r = in_r;
assign in_9_15_i = in_i;
assign in_9_16_r = in_r;
assign in_9_16_i = in_i;
assign in_9_17_r = in_r;
assign in_9_17_i = in_i;
assign in_9_18_r = in_r;
assign in_9_18_i = in_i;
assign in_9_19_r = in_r;
assign in_9_19_i = in_i;
assign in_9_20_r = in_r;
assign in_9_20_i = in_i;
assign in_9_21_r = in_r;
assign in_9_21_i = in_i;
assign in_9_22_r = in_r;
assign in_9_22_i = in_i;
assign in_9_23_r = in_r;
assign in_9_23_i = in_i;
assign in_9_24_r = in_r;
assign in_9_24_i = in_i;
assign in_9_25_r = in_r;
assign in_9_25_i = in_i;
assign in_9_26_r = in_r;
assign in_9_26_i = in_i;
assign in_9_27_r = in_r;
assign in_9_27_i = in_i;
assign in_9_28_r = in_r;
assign in_9_28_i = in_i;
assign in_9_29_r = in_r;
assign in_9_29_i = in_i;
assign in_9_30_r = in_r;
assign in_9_30_i = in_i;
assign in_9_31_r = in_r;
assign in_9_31_i = in_i;
assign in_9_32_r = in_r;
assign in_9_32_i = in_i;
assign in_10_1_r = in_r;
assign in_10_1_i = in_i;
assign in_10_2_r = in_r;
assign in_10_2_i = in_i;
assign in_10_3_r = in_r;
assign in_10_3_i = in_i;
assign in_10_4_r = in_r;
assign in_10_4_i = in_i;
assign in_10_5_r = in_r;
assign in_10_5_i = in_i;
assign in_10_6_r = in_r;
assign in_10_6_i = in_i;
assign in_10_7_r = in_r;
assign in_10_7_i = in_i;
assign in_10_8_r = in_r;
assign in_10_8_i = in_i;
assign in_10_9_r = in_r;
assign in_10_9_i = in_i;
assign in_10_10_r = in_r;
assign in_10_10_i = in_i;
assign in_10_11_r = in_r;
assign in_10_11_i = in_i;
assign in_10_12_r = in_r;
assign in_10_12_i = in_i;
assign in_10_13_r = in_r;
assign in_10_13_i = in_i;
assign in_10_14_r = in_r;
assign in_10_14_i = in_i;
assign in_10_15_r = in_r;
assign in_10_15_i = in_i;
assign in_10_16_r = in_r;
assign in_10_16_i = in_i;
assign in_10_17_r = in_r;
assign in_10_17_i = in_i;
assign in_10_18_r = in_r;
assign in_10_18_i = in_i;
assign in_10_19_r = in_r;
assign in_10_19_i = in_i;
assign in_10_20_r = in_r;
assign in_10_20_i = in_i;
assign in_10_21_r = in_r;
assign in_10_21_i = in_i;
assign in_10_22_r = in_r;
assign in_10_22_i = in_i;
assign in_10_23_r = in_r;
assign in_10_23_i = in_i;
assign in_10_24_r = in_r;
assign in_10_24_i = in_i;
assign in_10_25_r = in_r;
assign in_10_25_i = in_i;
assign in_10_26_r = in_r;
assign in_10_26_i = in_i;
assign in_10_27_r = in_r;
assign in_10_27_i = in_i;
assign in_10_28_r = in_r;
assign in_10_28_i = in_i;
assign in_10_29_r = in_r;
assign in_10_29_i = in_i;
assign in_10_30_r = in_r;
assign in_10_30_i = in_i;
assign in_10_31_r = in_r;
assign in_10_31_i = in_i;
assign in_10_32_r = in_r;
assign in_10_32_i = in_i;
assign in_11_1_r = in_r;
assign in_11_1_i = in_i;
assign in_11_2_r = in_r;
assign in_11_2_i = in_i;
assign in_11_3_r = in_r;
assign in_11_3_i = in_i;
assign in_11_4_r = in_r;
assign in_11_4_i = in_i;
assign in_11_5_r = in_r;
assign in_11_5_i = in_i;
assign in_11_6_r = in_r;
assign in_11_6_i = in_i;
assign in_11_7_r = in_r;
assign in_11_7_i = in_i;
assign in_11_8_r = in_r;
assign in_11_8_i = in_i;
assign in_11_9_r = in_r;
assign in_11_9_i = in_i;
assign in_11_10_r = in_r;
assign in_11_10_i = in_i;
assign in_11_11_r = in_r;
assign in_11_11_i = in_i;
assign in_11_12_r = in_r;
assign in_11_12_i = in_i;
assign in_11_13_r = in_r;
assign in_11_13_i = in_i;
assign in_11_14_r = in_r;
assign in_11_14_i = in_i;
assign in_11_15_r = in_r;
assign in_11_15_i = in_i;
assign in_11_16_r = in_r;
assign in_11_16_i = in_i;
assign in_11_17_r = in_r;
assign in_11_17_i = in_i;
assign in_11_18_r = in_r;
assign in_11_18_i = in_i;
assign in_11_19_r = in_r;
assign in_11_19_i = in_i;
assign in_11_20_r = in_r;
assign in_11_20_i = in_i;
assign in_11_21_r = in_r;
assign in_11_21_i = in_i;
assign in_11_22_r = in_r;
assign in_11_22_i = in_i;
assign in_11_23_r = in_r;
assign in_11_23_i = in_i;
assign in_11_24_r = in_r;
assign in_11_24_i = in_i;
assign in_11_25_r = in_r;
assign in_11_25_i = in_i;
assign in_11_26_r = in_r;
assign in_11_26_i = in_i;
assign in_11_27_r = in_r;
assign in_11_27_i = in_i;
assign in_11_28_r = in_r;
assign in_11_28_i = in_i;
assign in_11_29_r = in_r;
assign in_11_29_i = in_i;
assign in_11_30_r = in_r;
assign in_11_30_i = in_i;
assign in_11_31_r = in_r;
assign in_11_31_i = in_i;
assign in_11_32_r = in_r;
assign in_11_32_i = in_i;
assign in_12_1_r = in_r;
assign in_12_1_i = in_i;
assign in_12_2_r = in_r;
assign in_12_2_i = in_i;
assign in_12_3_r = in_r;
assign in_12_3_i = in_i;
assign in_12_4_r = in_r;
assign in_12_4_i = in_i;
assign in_12_5_r = in_r;
assign in_12_5_i = in_i;
assign in_12_6_r = in_r;
assign in_12_6_i = in_i;
assign in_12_7_r = in_r;
assign in_12_7_i = in_i;
assign in_12_8_r = in_r;
assign in_12_8_i = in_i;
assign in_12_9_r = in_r;
assign in_12_9_i = in_i;
assign in_12_10_r = in_r;
assign in_12_10_i = in_i;
assign in_12_11_r = in_r;
assign in_12_11_i = in_i;
assign in_12_12_r = in_r;
assign in_12_12_i = in_i;
assign in_12_13_r = in_r;
assign in_12_13_i = in_i;
assign in_12_14_r = in_r;
assign in_12_14_i = in_i;
assign in_12_15_r = in_r;
assign in_12_15_i = in_i;
assign in_12_16_r = in_r;
assign in_12_16_i = in_i;
assign in_12_17_r = in_r;
assign in_12_17_i = in_i;
assign in_12_18_r = in_r;
assign in_12_18_i = in_i;
assign in_12_19_r = in_r;
assign in_12_19_i = in_i;
assign in_12_20_r = in_r;
assign in_12_20_i = in_i;
assign in_12_21_r = in_r;
assign in_12_21_i = in_i;
assign in_12_22_r = in_r;
assign in_12_22_i = in_i;
assign in_12_23_r = in_r;
assign in_12_23_i = in_i;
assign in_12_24_r = in_r;
assign in_12_24_i = in_i;
assign in_12_25_r = in_r;
assign in_12_25_i = in_i;
assign in_12_26_r = in_r;
assign in_12_26_i = in_i;
assign in_12_27_r = in_r;
assign in_12_27_i = in_i;
assign in_12_28_r = in_r;
assign in_12_28_i = in_i;
assign in_12_29_r = in_r;
assign in_12_29_i = in_i;
assign in_12_30_r = in_r;
assign in_12_30_i = in_i;
assign in_12_31_r = in_r;
assign in_12_31_i = in_i;
assign in_12_32_r = in_r;
assign in_12_32_i = in_i;
assign in_13_1_r = in_r;
assign in_13_1_i = in_i;
assign in_13_2_r = in_r;
assign in_13_2_i = in_i;
assign in_13_3_r = in_r;
assign in_13_3_i = in_i;
assign in_13_4_r = in_r;
assign in_13_4_i = in_i;
assign in_13_5_r = in_r;
assign in_13_5_i = in_i;
assign in_13_6_r = in_r;
assign in_13_6_i = in_i;
assign in_13_7_r = in_r;
assign in_13_7_i = in_i;
assign in_13_8_r = in_r;
assign in_13_8_i = in_i;
assign in_13_9_r = in_r;
assign in_13_9_i = in_i;
assign in_13_10_r = in_r;
assign in_13_10_i = in_i;
assign in_13_11_r = in_r;
assign in_13_11_i = in_i;
assign in_13_12_r = in_r;
assign in_13_12_i = in_i;
assign in_13_13_r = in_r;
assign in_13_13_i = in_i;
assign in_13_14_r = in_r;
assign in_13_14_i = in_i;
assign in_13_15_r = in_r;
assign in_13_15_i = in_i;
assign in_13_16_r = in_r;
assign in_13_16_i = in_i;
assign in_13_17_r = in_r;
assign in_13_17_i = in_i;
assign in_13_18_r = in_r;
assign in_13_18_i = in_i;
assign in_13_19_r = in_r;
assign in_13_19_i = in_i;
assign in_13_20_r = in_r;
assign in_13_20_i = in_i;
assign in_13_21_r = in_r;
assign in_13_21_i = in_i;
assign in_13_22_r = in_r;
assign in_13_22_i = in_i;
assign in_13_23_r = in_r;
assign in_13_23_i = in_i;
assign in_13_24_r = in_r;
assign in_13_24_i = in_i;
assign in_13_25_r = in_r;
assign in_13_25_i = in_i;
assign in_13_26_r = in_r;
assign in_13_26_i = in_i;
assign in_13_27_r = in_r;
assign in_13_27_i = in_i;
assign in_13_28_r = in_r;
assign in_13_28_i = in_i;
assign in_13_29_r = in_r;
assign in_13_29_i = in_i;
assign in_13_30_r = in_r;
assign in_13_30_i = in_i;
assign in_13_31_r = in_r;
assign in_13_31_i = in_i;
assign in_13_32_r = in_r;
assign in_13_32_i = in_i;
assign in_14_1_r = in_r;
assign in_14_1_i = in_i;
assign in_14_2_r = in_r;
assign in_14_2_i = in_i;
assign in_14_3_r = in_r;
assign in_14_3_i = in_i;
assign in_14_4_r = in_r;
assign in_14_4_i = in_i;
assign in_14_5_r = in_r;
assign in_14_5_i = in_i;
assign in_14_6_r = in_r;
assign in_14_6_i = in_i;
assign in_14_7_r = in_r;
assign in_14_7_i = in_i;
assign in_14_8_r = in_r;
assign in_14_8_i = in_i;
assign in_14_9_r = in_r;
assign in_14_9_i = in_i;
assign in_14_10_r = in_r;
assign in_14_10_i = in_i;
assign in_14_11_r = in_r;
assign in_14_11_i = in_i;
assign in_14_12_r = in_r;
assign in_14_12_i = in_i;
assign in_14_13_r = in_r;
assign in_14_13_i = in_i;
assign in_14_14_r = in_r;
assign in_14_14_i = in_i;
assign in_14_15_r = in_r;
assign in_14_15_i = in_i;
assign in_14_16_r = in_r;
assign in_14_16_i = in_i;
assign in_14_17_r = in_r;
assign in_14_17_i = in_i;
assign in_14_18_r = in_r;
assign in_14_18_i = in_i;
assign in_14_19_r = in_r;
assign in_14_19_i = in_i;
assign in_14_20_r = in_r;
assign in_14_20_i = in_i;
assign in_14_21_r = in_r;
assign in_14_21_i = in_i;
assign in_14_22_r = in_r;
assign in_14_22_i = in_i;
assign in_14_23_r = in_r;
assign in_14_23_i = in_i;
assign in_14_24_r = in_r;
assign in_14_24_i = in_i;
assign in_14_25_r = in_r;
assign in_14_25_i = in_i;
assign in_14_26_r = in_r;
assign in_14_26_i = in_i;
assign in_14_27_r = in_r;
assign in_14_27_i = in_i;
assign in_14_28_r = in_r;
assign in_14_28_i = in_i;
assign in_14_29_r = in_r;
assign in_14_29_i = in_i;
assign in_14_30_r = in_r;
assign in_14_30_i = in_i;
assign in_14_31_r = in_r;
assign in_14_31_i = in_i;
assign in_14_32_r = in_r;
assign in_14_32_i = in_i;
assign in_15_1_r = in_r;
assign in_15_1_i = in_i;
assign in_15_2_r = in_r;
assign in_15_2_i = in_i;
assign in_15_3_r = in_r;
assign in_15_3_i = in_i;
assign in_15_4_r = in_r;
assign in_15_4_i = in_i;
assign in_15_5_r = in_r;
assign in_15_5_i = in_i;
assign in_15_6_r = in_r;
assign in_15_6_i = in_i;
assign in_15_7_r = in_r;
assign in_15_7_i = in_i;
assign in_15_8_r = in_r;
assign in_15_8_i = in_i;
assign in_15_9_r = in_r;
assign in_15_9_i = in_i;
assign in_15_10_r = in_r;
assign in_15_10_i = in_i;
assign in_15_11_r = in_r;
assign in_15_11_i = in_i;
assign in_15_12_r = in_r;
assign in_15_12_i = in_i;
assign in_15_13_r = in_r;
assign in_15_13_i = in_i;
assign in_15_14_r = in_r;
assign in_15_14_i = in_i;
assign in_15_15_r = in_r;
assign in_15_15_i = in_i;
assign in_15_16_r = in_r;
assign in_15_16_i = in_i;
assign in_15_17_r = in_r;
assign in_15_17_i = in_i;
assign in_15_18_r = in_r;
assign in_15_18_i = in_i;
assign in_15_19_r = in_r;
assign in_15_19_i = in_i;
assign in_15_20_r = in_r;
assign in_15_20_i = in_i;
assign in_15_21_r = in_r;
assign in_15_21_i = in_i;
assign in_15_22_r = in_r;
assign in_15_22_i = in_i;
assign in_15_23_r = in_r;
assign in_15_23_i = in_i;
assign in_15_24_r = in_r;
assign in_15_24_i = in_i;
assign in_15_25_r = in_r;
assign in_15_25_i = in_i;
assign in_15_26_r = in_r;
assign in_15_26_i = in_i;
assign in_15_27_r = in_r;
assign in_15_27_i = in_i;
assign in_15_28_r = in_r;
assign in_15_28_i = in_i;
assign in_15_29_r = in_r;
assign in_15_29_i = in_i;
assign in_15_30_r = in_r;
assign in_15_30_i = in_i;
assign in_15_31_r = in_r;
assign in_15_31_i = in_i;
assign in_15_32_r = in_r;
assign in_15_32_i = in_i;
assign in_16_1_r = in_r;
assign in_16_1_i = in_i;
assign in_16_2_r = in_r;
assign in_16_2_i = in_i;
assign in_16_3_r = in_r;
assign in_16_3_i = in_i;
assign in_16_4_r = in_r;
assign in_16_4_i = in_i;
assign in_16_5_r = in_r;
assign in_16_5_i = in_i;
assign in_16_6_r = in_r;
assign in_16_6_i = in_i;
assign in_16_7_r = in_r;
assign in_16_7_i = in_i;
assign in_16_8_r = in_r;
assign in_16_8_i = in_i;
assign in_16_9_r = in_r;
assign in_16_9_i = in_i;
assign in_16_10_r = in_r;
assign in_16_10_i = in_i;
assign in_16_11_r = in_r;
assign in_16_11_i = in_i;
assign in_16_12_r = in_r;
assign in_16_12_i = in_i;
assign in_16_13_r = in_r;
assign in_16_13_i = in_i;
assign in_16_14_r = in_r;
assign in_16_14_i = in_i;
assign in_16_15_r = in_r;
assign in_16_15_i = in_i;
assign in_16_16_r = in_r;
assign in_16_16_i = in_i;
assign in_16_17_r = in_r;
assign in_16_17_i = in_i;
assign in_16_18_r = in_r;
assign in_16_18_i = in_i;
assign in_16_19_r = in_r;
assign in_16_19_i = in_i;
assign in_16_20_r = in_r;
assign in_16_20_i = in_i;
assign in_16_21_r = in_r;
assign in_16_21_i = in_i;
assign in_16_22_r = in_r;
assign in_16_22_i = in_i;
assign in_16_23_r = in_r;
assign in_16_23_i = in_i;
assign in_16_24_r = in_r;
assign in_16_24_i = in_i;
assign in_16_25_r = in_r;
assign in_16_25_i = in_i;
assign in_16_26_r = in_r;
assign in_16_26_i = in_i;
assign in_16_27_r = in_r;
assign in_16_27_i = in_i;
assign in_16_28_r = in_r;
assign in_16_28_i = in_i;
assign in_16_29_r = in_r;
assign in_16_29_i = in_i;
assign in_16_30_r = in_r;
assign in_16_30_i = in_i;
assign in_16_31_r = in_r;
assign in_16_31_i = in_i;
assign in_16_32_r = in_r;
assign in_16_32_i = in_i;
assign in_17_1_r = in_r;
assign in_17_1_i = in_i;
assign in_17_2_r = in_r;
assign in_17_2_i = in_i;
assign in_17_3_r = in_r;
assign in_17_3_i = in_i;
assign in_17_4_r = in_r;
assign in_17_4_i = in_i;
assign in_17_5_r = in_r;
assign in_17_5_i = in_i;
assign in_17_6_r = in_r;
assign in_17_6_i = in_i;
assign in_17_7_r = in_r;
assign in_17_7_i = in_i;
assign in_17_8_r = in_r;
assign in_17_8_i = in_i;
assign in_17_9_r = in_r;
assign in_17_9_i = in_i;
assign in_17_10_r = in_r;
assign in_17_10_i = in_i;
assign in_17_11_r = in_r;
assign in_17_11_i = in_i;
assign in_17_12_r = in_r;
assign in_17_12_i = in_i;
assign in_17_13_r = in_r;
assign in_17_13_i = in_i;
assign in_17_14_r = in_r;
assign in_17_14_i = in_i;
assign in_17_15_r = in_r;
assign in_17_15_i = in_i;
assign in_17_16_r = in_r;
assign in_17_16_i = in_i;
assign in_17_17_r = in_r;
assign in_17_17_i = in_i;
assign in_17_18_r = in_r;
assign in_17_18_i = in_i;
assign in_17_19_r = in_r;
assign in_17_19_i = in_i;
assign in_17_20_r = in_r;
assign in_17_20_i = in_i;
assign in_17_21_r = in_r;
assign in_17_21_i = in_i;
assign in_17_22_r = in_r;
assign in_17_22_i = in_i;
assign in_17_23_r = in_r;
assign in_17_23_i = in_i;
assign in_17_24_r = in_r;
assign in_17_24_i = in_i;
assign in_17_25_r = in_r;
assign in_17_25_i = in_i;
assign in_17_26_r = in_r;
assign in_17_26_i = in_i;
assign in_17_27_r = in_r;
assign in_17_27_i = in_i;
assign in_17_28_r = in_r;
assign in_17_28_i = in_i;
assign in_17_29_r = in_r;
assign in_17_29_i = in_i;
assign in_17_30_r = in_r;
assign in_17_30_i = in_i;
assign in_17_31_r = in_r;
assign in_17_31_i = in_i;
assign in_17_32_r = in_r;
assign in_17_32_i = in_i;
assign in_18_1_r = in_r;
assign in_18_1_i = in_i;
assign in_18_2_r = in_r;
assign in_18_2_i = in_i;
assign in_18_3_r = in_r;
assign in_18_3_i = in_i;
assign in_18_4_r = in_r;
assign in_18_4_i = in_i;
assign in_18_5_r = in_r;
assign in_18_5_i = in_i;
assign in_18_6_r = in_r;
assign in_18_6_i = in_i;
assign in_18_7_r = in_r;
assign in_18_7_i = in_i;
assign in_18_8_r = in_r;
assign in_18_8_i = in_i;
assign in_18_9_r = in_r;
assign in_18_9_i = in_i;
assign in_18_10_r = in_r;
assign in_18_10_i = in_i;
assign in_18_11_r = in_r;
assign in_18_11_i = in_i;
assign in_18_12_r = in_r;
assign in_18_12_i = in_i;
assign in_18_13_r = in_r;
assign in_18_13_i = in_i;
assign in_18_14_r = in_r;
assign in_18_14_i = in_i;
assign in_18_15_r = in_r;
assign in_18_15_i = in_i;
assign in_18_16_r = in_r;
assign in_18_16_i = in_i;
assign in_18_17_r = in_r;
assign in_18_17_i = in_i;
assign in_18_18_r = in_r;
assign in_18_18_i = in_i;
assign in_18_19_r = in_r;
assign in_18_19_i = in_i;
assign in_18_20_r = in_r;
assign in_18_20_i = in_i;
assign in_18_21_r = in_r;
assign in_18_21_i = in_i;
assign in_18_22_r = in_r;
assign in_18_22_i = in_i;
assign in_18_23_r = in_r;
assign in_18_23_i = in_i;
assign in_18_24_r = in_r;
assign in_18_24_i = in_i;
assign in_18_25_r = in_r;
assign in_18_25_i = in_i;
assign in_18_26_r = in_r;
assign in_18_26_i = in_i;
assign in_18_27_r = in_r;
assign in_18_27_i = in_i;
assign in_18_28_r = in_r;
assign in_18_28_i = in_i;
assign in_18_29_r = in_r;
assign in_18_29_i = in_i;
assign in_18_30_r = in_r;
assign in_18_30_i = in_i;
assign in_18_31_r = in_r;
assign in_18_31_i = in_i;
assign in_18_32_r = in_r;
assign in_18_32_i = in_i;
assign in_19_1_r = in_r;
assign in_19_1_i = in_i;
assign in_19_2_r = in_r;
assign in_19_2_i = in_i;
assign in_19_3_r = in_r;
assign in_19_3_i = in_i;
assign in_19_4_r = in_r;
assign in_19_4_i = in_i;
assign in_19_5_r = in_r;
assign in_19_5_i = in_i;
assign in_19_6_r = in_r;
assign in_19_6_i = in_i;
assign in_19_7_r = in_r;
assign in_19_7_i = in_i;
assign in_19_8_r = in_r;
assign in_19_8_i = in_i;
assign in_19_9_r = in_r;
assign in_19_9_i = in_i;
assign in_19_10_r = in_r;
assign in_19_10_i = in_i;
assign in_19_11_r = in_r;
assign in_19_11_i = in_i;
assign in_19_12_r = in_r;
assign in_19_12_i = in_i;
assign in_19_13_r = in_r;
assign in_19_13_i = in_i;
assign in_19_14_r = in_r;
assign in_19_14_i = in_i;
assign in_19_15_r = in_r;
assign in_19_15_i = in_i;
assign in_19_16_r = in_r;
assign in_19_16_i = in_i;
assign in_19_17_r = in_r;
assign in_19_17_i = in_i;
assign in_19_18_r = in_r;
assign in_19_18_i = in_i;
assign in_19_19_r = in_r;
assign in_19_19_i = in_i;
assign in_19_20_r = in_r;
assign in_19_20_i = in_i;
assign in_19_21_r = in_r;
assign in_19_21_i = in_i;
assign in_19_22_r = in_r;
assign in_19_22_i = in_i;
assign in_19_23_r = in_r;
assign in_19_23_i = in_i;
assign in_19_24_r = in_r;
assign in_19_24_i = in_i;
assign in_19_25_r = in_r;
assign in_19_25_i = in_i;
assign in_19_26_r = in_r;
assign in_19_26_i = in_i;
assign in_19_27_r = in_r;
assign in_19_27_i = in_i;
assign in_19_28_r = in_r;
assign in_19_28_i = in_i;
assign in_19_29_r = in_r;
assign in_19_29_i = in_i;
assign in_19_30_r = in_r;
assign in_19_30_i = in_i;
assign in_19_31_r = in_r;
assign in_19_31_i = in_i;
assign in_19_32_r = in_r;
assign in_19_32_i = in_i;
assign in_20_1_r = in_r;
assign in_20_1_i = in_i;
assign in_20_2_r = in_r;
assign in_20_2_i = in_i;
assign in_20_3_r = in_r;
assign in_20_3_i = in_i;
assign in_20_4_r = in_r;
assign in_20_4_i = in_i;
assign in_20_5_r = in_r;
assign in_20_5_i = in_i;
assign in_20_6_r = in_r;
assign in_20_6_i = in_i;
assign in_20_7_r = in_r;
assign in_20_7_i = in_i;
assign in_20_8_r = in_r;
assign in_20_8_i = in_i;
assign in_20_9_r = in_r;
assign in_20_9_i = in_i;
assign in_20_10_r = in_r;
assign in_20_10_i = in_i;
assign in_20_11_r = in_r;
assign in_20_11_i = in_i;
assign in_20_12_r = in_r;
assign in_20_12_i = in_i;
assign in_20_13_r = in_r;
assign in_20_13_i = in_i;
assign in_20_14_r = in_r;
assign in_20_14_i = in_i;
assign in_20_15_r = in_r;
assign in_20_15_i = in_i;
assign in_20_16_r = in_r;
assign in_20_16_i = in_i;
assign in_20_17_r = in_r;
assign in_20_17_i = in_i;
assign in_20_18_r = in_r;
assign in_20_18_i = in_i;
assign in_20_19_r = in_r;
assign in_20_19_i = in_i;
assign in_20_20_r = in_r;
assign in_20_20_i = in_i;
assign in_20_21_r = in_r;
assign in_20_21_i = in_i;
assign in_20_22_r = in_r;
assign in_20_22_i = in_i;
assign in_20_23_r = in_r;
assign in_20_23_i = in_i;
assign in_20_24_r = in_r;
assign in_20_24_i = in_i;
assign in_20_25_r = in_r;
assign in_20_25_i = in_i;
assign in_20_26_r = in_r;
assign in_20_26_i = in_i;
assign in_20_27_r = in_r;
assign in_20_27_i = in_i;
assign in_20_28_r = in_r;
assign in_20_28_i = in_i;
assign in_20_29_r = in_r;
assign in_20_29_i = in_i;
assign in_20_30_r = in_r;
assign in_20_30_i = in_i;
assign in_20_31_r = in_r;
assign in_20_31_i = in_i;
assign in_20_32_r = in_r;
assign in_20_32_i = in_i;
assign in_21_1_r = in_r;
assign in_21_1_i = in_i;
assign in_21_2_r = in_r;
assign in_21_2_i = in_i;
assign in_21_3_r = in_r;
assign in_21_3_i = in_i;
assign in_21_4_r = in_r;
assign in_21_4_i = in_i;
assign in_21_5_r = in_r;
assign in_21_5_i = in_i;
assign in_21_6_r = in_r;
assign in_21_6_i = in_i;
assign in_21_7_r = in_r;
assign in_21_7_i = in_i;
assign in_21_8_r = in_r;
assign in_21_8_i = in_i;
assign in_21_9_r = in_r;
assign in_21_9_i = in_i;
assign in_21_10_r = in_r;
assign in_21_10_i = in_i;
assign in_21_11_r = in_r;
assign in_21_11_i = in_i;
assign in_21_12_r = in_r;
assign in_21_12_i = in_i;
assign in_21_13_r = in_r;
assign in_21_13_i = in_i;
assign in_21_14_r = in_r;
assign in_21_14_i = in_i;
assign in_21_15_r = in_r;
assign in_21_15_i = in_i;
assign in_21_16_r = in_r;
assign in_21_16_i = in_i;
assign in_21_17_r = in_r;
assign in_21_17_i = in_i;
assign in_21_18_r = in_r;
assign in_21_18_i = in_i;
assign in_21_19_r = in_r;
assign in_21_19_i = in_i;
assign in_21_20_r = in_r;
assign in_21_20_i = in_i;
assign in_21_21_r = in_r;
assign in_21_21_i = in_i;
assign in_21_22_r = in_r;
assign in_21_22_i = in_i;
assign in_21_23_r = in_r;
assign in_21_23_i = in_i;
assign in_21_24_r = in_r;
assign in_21_24_i = in_i;
assign in_21_25_r = in_r;
assign in_21_25_i = in_i;
assign in_21_26_r = in_r;
assign in_21_26_i = in_i;
assign in_21_27_r = in_r;
assign in_21_27_i = in_i;
assign in_21_28_r = in_r;
assign in_21_28_i = in_i;
assign in_21_29_r = in_r;
assign in_21_29_i = in_i;
assign in_21_30_r = in_r;
assign in_21_30_i = in_i;
assign in_21_31_r = in_r;
assign in_21_31_i = in_i;
assign in_21_32_r = in_r;
assign in_21_32_i = in_i;
assign in_22_1_r = in_r;
assign in_22_1_i = in_i;
assign in_22_2_r = in_r;
assign in_22_2_i = in_i;
assign in_22_3_r = in_r;
assign in_22_3_i = in_i;
assign in_22_4_r = in_r;
assign in_22_4_i = in_i;
assign in_22_5_r = in_r;
assign in_22_5_i = in_i;
assign in_22_6_r = in_r;
assign in_22_6_i = in_i;
assign in_22_7_r = in_r;
assign in_22_7_i = in_i;
assign in_22_8_r = in_r;
assign in_22_8_i = in_i;
assign in_22_9_r = in_r;
assign in_22_9_i = in_i;
assign in_22_10_r = in_r;
assign in_22_10_i = in_i;
assign in_22_11_r = in_r;
assign in_22_11_i = in_i;
assign in_22_12_r = in_r;
assign in_22_12_i = in_i;
assign in_22_13_r = in_r;
assign in_22_13_i = in_i;
assign in_22_14_r = in_r;
assign in_22_14_i = in_i;
assign in_22_15_r = in_r;
assign in_22_15_i = in_i;
assign in_22_16_r = in_r;
assign in_22_16_i = in_i;
assign in_22_17_r = in_r;
assign in_22_17_i = in_i;
assign in_22_18_r = in_r;
assign in_22_18_i = in_i;
assign in_22_19_r = in_r;
assign in_22_19_i = in_i;
assign in_22_20_r = in_r;
assign in_22_20_i = in_i;
assign in_22_21_r = in_r;
assign in_22_21_i = in_i;
assign in_22_22_r = in_r;
assign in_22_22_i = in_i;
assign in_22_23_r = in_r;
assign in_22_23_i = in_i;
assign in_22_24_r = in_r;
assign in_22_24_i = in_i;
assign in_22_25_r = in_r;
assign in_22_25_i = in_i;
assign in_22_26_r = in_r;
assign in_22_26_i = in_i;
assign in_22_27_r = in_r;
assign in_22_27_i = in_i;
assign in_22_28_r = in_r;
assign in_22_28_i = in_i;
assign in_22_29_r = in_r;
assign in_22_29_i = in_i;
assign in_22_30_r = in_r;
assign in_22_30_i = in_i;
assign in_22_31_r = in_r;
assign in_22_31_i = in_i;
assign in_22_32_r = in_r;
assign in_22_32_i = in_i;
assign in_23_1_r = in_r;
assign in_23_1_i = in_i;
assign in_23_2_r = in_r;
assign in_23_2_i = in_i;
assign in_23_3_r = in_r;
assign in_23_3_i = in_i;
assign in_23_4_r = in_r;
assign in_23_4_i = in_i;
assign in_23_5_r = in_r;
assign in_23_5_i = in_i;
assign in_23_6_r = in_r;
assign in_23_6_i = in_i;
assign in_23_7_r = in_r;
assign in_23_7_i = in_i;
assign in_23_8_r = in_r;
assign in_23_8_i = in_i;
assign in_23_9_r = in_r;
assign in_23_9_i = in_i;
assign in_23_10_r = in_r;
assign in_23_10_i = in_i;
assign in_23_11_r = in_r;
assign in_23_11_i = in_i;
assign in_23_12_r = in_r;
assign in_23_12_i = in_i;
assign in_23_13_r = in_r;
assign in_23_13_i = in_i;
assign in_23_14_r = in_r;
assign in_23_14_i = in_i;
assign in_23_15_r = in_r;
assign in_23_15_i = in_i;
assign in_23_16_r = in_r;
assign in_23_16_i = in_i;
assign in_23_17_r = in_r;
assign in_23_17_i = in_i;
assign in_23_18_r = in_r;
assign in_23_18_i = in_i;
assign in_23_19_r = in_r;
assign in_23_19_i = in_i;
assign in_23_20_r = in_r;
assign in_23_20_i = in_i;
assign in_23_21_r = in_r;
assign in_23_21_i = in_i;
assign in_23_22_r = in_r;
assign in_23_22_i = in_i;
assign in_23_23_r = in_r;
assign in_23_23_i = in_i;
assign in_23_24_r = in_r;
assign in_23_24_i = in_i;
assign in_23_25_r = in_r;
assign in_23_25_i = in_i;
assign in_23_26_r = in_r;
assign in_23_26_i = in_i;
assign in_23_27_r = in_r;
assign in_23_27_i = in_i;
assign in_23_28_r = in_r;
assign in_23_28_i = in_i;
assign in_23_29_r = in_r;
assign in_23_29_i = in_i;
assign in_23_30_r = in_r;
assign in_23_30_i = in_i;
assign in_23_31_r = in_r;
assign in_23_31_i = in_i;
assign in_23_32_r = in_r;
assign in_23_32_i = in_i;
assign in_24_1_r = in_r;
assign in_24_1_i = in_i;
assign in_24_2_r = in_r;
assign in_24_2_i = in_i;
assign in_24_3_r = in_r;
assign in_24_3_i = in_i;
assign in_24_4_r = in_r;
assign in_24_4_i = in_i;
assign in_24_5_r = in_r;
assign in_24_5_i = in_i;
assign in_24_6_r = in_r;
assign in_24_6_i = in_i;
assign in_24_7_r = in_r;
assign in_24_7_i = in_i;
assign in_24_8_r = in_r;
assign in_24_8_i = in_i;
assign in_24_9_r = in_r;
assign in_24_9_i = in_i;
assign in_24_10_r = in_r;
assign in_24_10_i = in_i;
assign in_24_11_r = in_r;
assign in_24_11_i = in_i;
assign in_24_12_r = in_r;
assign in_24_12_i = in_i;
assign in_24_13_r = in_r;
assign in_24_13_i = in_i;
assign in_24_14_r = in_r;
assign in_24_14_i = in_i;
assign in_24_15_r = in_r;
assign in_24_15_i = in_i;
assign in_24_16_r = in_r;
assign in_24_16_i = in_i;
assign in_24_17_r = in_r;
assign in_24_17_i = in_i;
assign in_24_18_r = in_r;
assign in_24_18_i = in_i;
assign in_24_19_r = in_r;
assign in_24_19_i = in_i;
assign in_24_20_r = in_r;
assign in_24_20_i = in_i;
assign in_24_21_r = in_r;
assign in_24_21_i = in_i;
assign in_24_22_r = in_r;
assign in_24_22_i = in_i;
assign in_24_23_r = in_r;
assign in_24_23_i = in_i;
assign in_24_24_r = in_r;
assign in_24_24_i = in_i;
assign in_24_25_r = in_r;
assign in_24_25_i = in_i;
assign in_24_26_r = in_r;
assign in_24_26_i = in_i;
assign in_24_27_r = in_r;
assign in_24_27_i = in_i;
assign in_24_28_r = in_r;
assign in_24_28_i = in_i;
assign in_24_29_r = in_r;
assign in_24_29_i = in_i;
assign in_24_30_r = in_r;
assign in_24_30_i = in_i;
assign in_24_31_r = in_r;
assign in_24_31_i = in_i;
assign in_24_32_r = in_r;
assign in_24_32_i = in_i;
assign in_25_1_r = in_r;
assign in_25_1_i = in_i;
assign in_25_2_r = in_r;
assign in_25_2_i = in_i;
assign in_25_3_r = in_r;
assign in_25_3_i = in_i;
assign in_25_4_r = in_r;
assign in_25_4_i = in_i;
assign in_25_5_r = in_r;
assign in_25_5_i = in_i;
assign in_25_6_r = in_r;
assign in_25_6_i = in_i;
assign in_25_7_r = in_r;
assign in_25_7_i = in_i;
assign in_25_8_r = in_r;
assign in_25_8_i = in_i;
assign in_25_9_r = in_r;
assign in_25_9_i = in_i;
assign in_25_10_r = in_r;
assign in_25_10_i = in_i;
assign in_25_11_r = in_r;
assign in_25_11_i = in_i;
assign in_25_12_r = in_r;
assign in_25_12_i = in_i;
assign in_25_13_r = in_r;
assign in_25_13_i = in_i;
assign in_25_14_r = in_r;
assign in_25_14_i = in_i;
assign in_25_15_r = in_r;
assign in_25_15_i = in_i;
assign in_25_16_r = in_r;
assign in_25_16_i = in_i;
assign in_25_17_r = in_r;
assign in_25_17_i = in_i;
assign in_25_18_r = in_r;
assign in_25_18_i = in_i;
assign in_25_19_r = in_r;
assign in_25_19_i = in_i;
assign in_25_20_r = in_r;
assign in_25_20_i = in_i;
assign in_25_21_r = in_r;
assign in_25_21_i = in_i;
assign in_25_22_r = in_r;
assign in_25_22_i = in_i;
assign in_25_23_r = in_r;
assign in_25_23_i = in_i;
assign in_25_24_r = in_r;
assign in_25_24_i = in_i;
assign in_25_25_r = in_r;
assign in_25_25_i = in_i;
assign in_25_26_r = in_r;
assign in_25_26_i = in_i;
assign in_25_27_r = in_r;
assign in_25_27_i = in_i;
assign in_25_28_r = in_r;
assign in_25_28_i = in_i;
assign in_25_29_r = in_r;
assign in_25_29_i = in_i;
assign in_25_30_r = in_r;
assign in_25_30_i = in_i;
assign in_25_31_r = in_r;
assign in_25_31_i = in_i;
assign in_25_32_r = in_r;
assign in_25_32_i = in_i;
assign in_26_1_r = in_r;
assign in_26_1_i = in_i;
assign in_26_2_r = in_r;
assign in_26_2_i = in_i;
assign in_26_3_r = in_r;
assign in_26_3_i = in_i;
assign in_26_4_r = in_r;
assign in_26_4_i = in_i;
assign in_26_5_r = in_r;
assign in_26_5_i = in_i;
assign in_26_6_r = in_r;
assign in_26_6_i = in_i;
assign in_26_7_r = in_r;
assign in_26_7_i = in_i;
assign in_26_8_r = in_r;
assign in_26_8_i = in_i;
assign in_26_9_r = in_r;
assign in_26_9_i = in_i;
assign in_26_10_r = in_r;
assign in_26_10_i = in_i;
assign in_26_11_r = in_r;
assign in_26_11_i = in_i;
assign in_26_12_r = in_r;
assign in_26_12_i = in_i;
assign in_26_13_r = in_r;
assign in_26_13_i = in_i;
assign in_26_14_r = in_r;
assign in_26_14_i = in_i;
assign in_26_15_r = in_r;
assign in_26_15_i = in_i;
assign in_26_16_r = in_r;
assign in_26_16_i = in_i;
assign in_26_17_r = in_r;
assign in_26_17_i = in_i;
assign in_26_18_r = in_r;
assign in_26_18_i = in_i;
assign in_26_19_r = in_r;
assign in_26_19_i = in_i;
assign in_26_20_r = in_r;
assign in_26_20_i = in_i;
assign in_26_21_r = in_r;
assign in_26_21_i = in_i;
assign in_26_22_r = in_r;
assign in_26_22_i = in_i;
assign in_26_23_r = in_r;
assign in_26_23_i = in_i;
assign in_26_24_r = in_r;
assign in_26_24_i = in_i;
assign in_26_25_r = in_r;
assign in_26_25_i = in_i;
assign in_26_26_r = in_r;
assign in_26_26_i = in_i;
assign in_26_27_r = in_r;
assign in_26_27_i = in_i;
assign in_26_28_r = in_r;
assign in_26_28_i = in_i;
assign in_26_29_r = in_r;
assign in_26_29_i = in_i;
assign in_26_30_r = in_r;
assign in_26_30_i = in_i;
assign in_26_31_r = in_r;
assign in_26_31_i = in_i;
assign in_26_32_r = in_r;
assign in_26_32_i = in_i;
assign in_27_1_r = in_r;
assign in_27_1_i = in_i;
assign in_27_2_r = in_r;
assign in_27_2_i = in_i;
assign in_27_3_r = in_r;
assign in_27_3_i = in_i;
assign in_27_4_r = in_r;
assign in_27_4_i = in_i;
assign in_27_5_r = in_r;
assign in_27_5_i = in_i;
assign in_27_6_r = in_r;
assign in_27_6_i = in_i;
assign in_27_7_r = in_r;
assign in_27_7_i = in_i;
assign in_27_8_r = in_r;
assign in_27_8_i = in_i;
assign in_27_9_r = in_r;
assign in_27_9_i = in_i;
assign in_27_10_r = in_r;
assign in_27_10_i = in_i;
assign in_27_11_r = in_r;
assign in_27_11_i = in_i;
assign in_27_12_r = in_r;
assign in_27_12_i = in_i;
assign in_27_13_r = in_r;
assign in_27_13_i = in_i;
assign in_27_14_r = in_r;
assign in_27_14_i = in_i;
assign in_27_15_r = in_r;
assign in_27_15_i = in_i;
assign in_27_16_r = in_r;
assign in_27_16_i = in_i;
assign in_27_17_r = in_r;
assign in_27_17_i = in_i;
assign in_27_18_r = in_r;
assign in_27_18_i = in_i;
assign in_27_19_r = in_r;
assign in_27_19_i = in_i;
assign in_27_20_r = in_r;
assign in_27_20_i = in_i;
assign in_27_21_r = in_r;
assign in_27_21_i = in_i;
assign in_27_22_r = in_r;
assign in_27_22_i = in_i;
assign in_27_23_r = in_r;
assign in_27_23_i = in_i;
assign in_27_24_r = in_r;
assign in_27_24_i = in_i;
assign in_27_25_r = in_r;
assign in_27_25_i = in_i;
assign in_27_26_r = in_r;
assign in_27_26_i = in_i;
assign in_27_27_r = in_r;
assign in_27_27_i = in_i;
assign in_27_28_r = in_r;
assign in_27_28_i = in_i;
assign in_27_29_r = in_r;
assign in_27_29_i = in_i;
assign in_27_30_r = in_r;
assign in_27_30_i = in_i;
assign in_27_31_r = in_r;
assign in_27_31_i = in_i;
assign in_27_32_r = in_r;
assign in_27_32_i = in_i;
assign in_28_1_r = in_r;
assign in_28_1_i = in_i;
assign in_28_2_r = in_r;
assign in_28_2_i = in_i;
assign in_28_3_r = in_r;
assign in_28_3_i = in_i;
assign in_28_4_r = in_r;
assign in_28_4_i = in_i;
assign in_28_5_r = in_r;
assign in_28_5_i = in_i;
assign in_28_6_r = in_r;
assign in_28_6_i = in_i;
assign in_28_7_r = in_r;
assign in_28_7_i = in_i;
assign in_28_8_r = in_r;
assign in_28_8_i = in_i;
assign in_28_9_r = in_r;
assign in_28_9_i = in_i;
assign in_28_10_r = in_r;
assign in_28_10_i = in_i;
assign in_28_11_r = in_r;
assign in_28_11_i = in_i;
assign in_28_12_r = in_r;
assign in_28_12_i = in_i;
assign in_28_13_r = in_r;
assign in_28_13_i = in_i;
assign in_28_14_r = in_r;
assign in_28_14_i = in_i;
assign in_28_15_r = in_r;
assign in_28_15_i = in_i;
assign in_28_16_r = in_r;
assign in_28_16_i = in_i;
assign in_28_17_r = in_r;
assign in_28_17_i = in_i;
assign in_28_18_r = in_r;
assign in_28_18_i = in_i;
assign in_28_19_r = in_r;
assign in_28_19_i = in_i;
assign in_28_20_r = in_r;
assign in_28_20_i = in_i;
assign in_28_21_r = in_r;
assign in_28_21_i = in_i;
assign in_28_22_r = in_r;
assign in_28_22_i = in_i;
assign in_28_23_r = in_r;
assign in_28_23_i = in_i;
assign in_28_24_r = in_r;
assign in_28_24_i = in_i;
assign in_28_25_r = in_r;
assign in_28_25_i = in_i;
assign in_28_26_r = in_r;
assign in_28_26_i = in_i;
assign in_28_27_r = in_r;
assign in_28_27_i = in_i;
assign in_28_28_r = in_r;
assign in_28_28_i = in_i;
assign in_28_29_r = in_r;
assign in_28_29_i = in_i;
assign in_28_30_r = in_r;
assign in_28_30_i = in_i;
assign in_28_31_r = in_r;
assign in_28_31_i = in_i;
assign in_28_32_r = in_r;
assign in_28_32_i = in_i;
assign in_29_1_r = in_r;
assign in_29_1_i = in_i;
assign in_29_2_r = in_r;
assign in_29_2_i = in_i;
assign in_29_3_r = in_r;
assign in_29_3_i = in_i;
assign in_29_4_r = in_r;
assign in_29_4_i = in_i;
assign in_29_5_r = in_r;
assign in_29_5_i = in_i;
assign in_29_6_r = in_r;
assign in_29_6_i = in_i;
assign in_29_7_r = in_r;
assign in_29_7_i = in_i;
assign in_29_8_r = in_r;
assign in_29_8_i = in_i;
assign in_29_9_r = in_r;
assign in_29_9_i = in_i;
assign in_29_10_r = in_r;
assign in_29_10_i = in_i;
assign in_29_11_r = in_r;
assign in_29_11_i = in_i;
assign in_29_12_r = in_r;
assign in_29_12_i = in_i;
assign in_29_13_r = in_r;
assign in_29_13_i = in_i;
assign in_29_14_r = in_r;
assign in_29_14_i = in_i;
assign in_29_15_r = in_r;
assign in_29_15_i = in_i;
assign in_29_16_r = in_r;
assign in_29_16_i = in_i;
assign in_29_17_r = in_r;
assign in_29_17_i = in_i;
assign in_29_18_r = in_r;
assign in_29_18_i = in_i;
assign in_29_19_r = in_r;
assign in_29_19_i = in_i;
assign in_29_20_r = in_r;
assign in_29_20_i = in_i;
assign in_29_21_r = in_r;
assign in_29_21_i = in_i;
assign in_29_22_r = in_r;
assign in_29_22_i = in_i;
assign in_29_23_r = in_r;
assign in_29_23_i = in_i;
assign in_29_24_r = in_r;
assign in_29_24_i = in_i;
assign in_29_25_r = in_r;
assign in_29_25_i = in_i;
assign in_29_26_r = in_r;
assign in_29_26_i = in_i;
assign in_29_27_r = in_r;
assign in_29_27_i = in_i;
assign in_29_28_r = in_r;
assign in_29_28_i = in_i;
assign in_29_29_r = in_r;
assign in_29_29_i = in_i;
assign in_29_30_r = in_r;
assign in_29_30_i = in_i;
assign in_29_31_r = in_r;
assign in_29_31_i = in_i;
assign in_29_32_r = in_r;
assign in_29_32_i = in_i;
assign in_30_1_r = in_r;
assign in_30_1_i = in_i;
assign in_30_2_r = in_r;
assign in_30_2_i = in_i;
assign in_30_3_r = in_r;
assign in_30_3_i = in_i;
assign in_30_4_r = in_r;
assign in_30_4_i = in_i;
assign in_30_5_r = in_r;
assign in_30_5_i = in_i;
assign in_30_6_r = in_r;
assign in_30_6_i = in_i;
assign in_30_7_r = in_r;
assign in_30_7_i = in_i;
assign in_30_8_r = in_r;
assign in_30_8_i = in_i;
assign in_30_9_r = in_r;
assign in_30_9_i = in_i;
assign in_30_10_r = in_r;
assign in_30_10_i = in_i;
assign in_30_11_r = in_r;
assign in_30_11_i = in_i;
assign in_30_12_r = in_r;
assign in_30_12_i = in_i;
assign in_30_13_r = in_r;
assign in_30_13_i = in_i;
assign in_30_14_r = in_r;
assign in_30_14_i = in_i;
assign in_30_15_r = in_r;
assign in_30_15_i = in_i;
assign in_30_16_r = in_r;
assign in_30_16_i = in_i;
assign in_30_17_r = in_r;
assign in_30_17_i = in_i;
assign in_30_18_r = in_r;
assign in_30_18_i = in_i;
assign in_30_19_r = in_r;
assign in_30_19_i = in_i;
assign in_30_20_r = in_r;
assign in_30_20_i = in_i;
assign in_30_21_r = in_r;
assign in_30_21_i = in_i;
assign in_30_22_r = in_r;
assign in_30_22_i = in_i;
assign in_30_23_r = in_r;
assign in_30_23_i = in_i;
assign in_30_24_r = in_r;
assign in_30_24_i = in_i;
assign in_30_25_r = in_r;
assign in_30_25_i = in_i;
assign in_30_26_r = in_r;
assign in_30_26_i = in_i;
assign in_30_27_r = in_r;
assign in_30_27_i = in_i;
assign in_30_28_r = in_r;
assign in_30_28_i = in_i;
assign in_30_29_r = in_r;
assign in_30_29_i = in_i;
assign in_30_30_r = in_r;
assign in_30_30_i = in_i;
assign in_30_31_r = in_r;
assign in_30_31_i = in_i;
assign in_30_32_r = in_r;
assign in_30_32_i = in_i;
assign in_31_1_r = in_r;
assign in_31_1_i = in_i;
assign in_31_2_r = in_r;
assign in_31_2_i = in_i;
assign in_31_3_r = in_r;
assign in_31_3_i = in_i;
assign in_31_4_r = in_r;
assign in_31_4_i = in_i;
assign in_31_5_r = in_r;
assign in_31_5_i = in_i;
assign in_31_6_r = in_r;
assign in_31_6_i = in_i;
assign in_31_7_r = in_r;
assign in_31_7_i = in_i;
assign in_31_8_r = in_r;
assign in_31_8_i = in_i;
assign in_31_9_r = in_r;
assign in_31_9_i = in_i;
assign in_31_10_r = in_r;
assign in_31_10_i = in_i;
assign in_31_11_r = in_r;
assign in_31_11_i = in_i;
assign in_31_12_r = in_r;
assign in_31_12_i = in_i;
assign in_31_13_r = in_r;
assign in_31_13_i = in_i;
assign in_31_14_r = in_r;
assign in_31_14_i = in_i;
assign in_31_15_r = in_r;
assign in_31_15_i = in_i;
assign in_31_16_r = in_r;
assign in_31_16_i = in_i;
assign in_31_17_r = in_r;
assign in_31_17_i = in_i;
assign in_31_18_r = in_r;
assign in_31_18_i = in_i;
assign in_31_19_r = in_r;
assign in_31_19_i = in_i;
assign in_31_20_r = in_r;
assign in_31_20_i = in_i;
assign in_31_21_r = in_r;
assign in_31_21_i = in_i;
assign in_31_22_r = in_r;
assign in_31_22_i = in_i;
assign in_31_23_r = in_r;
assign in_31_23_i = in_i;
assign in_31_24_r = in_r;
assign in_31_24_i = in_i;
assign in_31_25_r = in_r;
assign in_31_25_i = in_i;
assign in_31_26_r = in_r;
assign in_31_26_i = in_i;
assign in_31_27_r = in_r;
assign in_31_27_i = in_i;
assign in_31_28_r = in_r;
assign in_31_28_i = in_i;
assign in_31_29_r = in_r;
assign in_31_29_i = in_i;
assign in_31_30_r = in_r;
assign in_31_30_i = in_i;
assign in_31_31_r = in_r;
assign in_31_31_i = in_i;
assign in_31_32_r = in_r;
assign in_31_32_i = in_i;
assign in_32_1_r = in_r;
assign in_32_1_i = in_i;
assign in_32_2_r = in_r;
assign in_32_2_i = in_i;
assign in_32_3_r = in_r;
assign in_32_3_i = in_i;
assign in_32_4_r = in_r;
assign in_32_4_i = in_i;
assign in_32_5_r = in_r;
assign in_32_5_i = in_i;
assign in_32_6_r = in_r;
assign in_32_6_i = in_i;
assign in_32_7_r = in_r;
assign in_32_7_i = in_i;
assign in_32_8_r = in_r;
assign in_32_8_i = in_i;
assign in_32_9_r = in_r;
assign in_32_9_i = in_i;
assign in_32_10_r = in_r;
assign in_32_10_i = in_i;
assign in_32_11_r = in_r;
assign in_32_11_i = in_i;
assign in_32_12_r = in_r;
assign in_32_12_i = in_i;
assign in_32_13_r = in_r;
assign in_32_13_i = in_i;
assign in_32_14_r = in_r;
assign in_32_14_i = in_i;
assign in_32_15_r = in_r;
assign in_32_15_i = in_i;
assign in_32_16_r = in_r;
assign in_32_16_i = in_i;
assign in_32_17_r = in_r;
assign in_32_17_i = in_i;
assign in_32_18_r = in_r;
assign in_32_18_i = in_i;
assign in_32_19_r = in_r;
assign in_32_19_i = in_i;
assign in_32_20_r = in_r;
assign in_32_20_i = in_i;
assign in_32_21_r = in_r;
assign in_32_21_i = in_i;
assign in_32_22_r = in_r;
assign in_32_22_i = in_i;
assign in_32_23_r = in_r;
assign in_32_23_i = in_i;
assign in_32_24_r = in_r;
assign in_32_24_i = in_i;
assign in_32_25_r = in_r;
assign in_32_25_i = in_i;
assign in_32_26_r = in_r;
assign in_32_26_i = in_i;
assign in_32_27_r = in_r;
assign in_32_27_i = in_i;
assign in_32_28_r = in_r;
assign in_32_28_i = in_i;
assign in_32_29_r = in_r;
assign in_32_29_i = in_i;
assign in_32_30_r = in_r;
assign in_32_30_i = in_i;
assign in_32_31_r = in_r;
assign in_32_31_i = in_i;
assign in_32_32_r = in_r;
assign in_32_32_i = in_i;

assign out_1_1_r = temp_b5_1_1_r;
assign out_1_1_i = temp_b5_1_1_i;
assign out_1_2_r = temp_b5_1_2_r;
assign out_1_2_i = temp_b5_1_2_i;
assign out_1_3_r = temp_b5_1_3_r;
assign out_1_3_i = temp_b5_1_3_i;
assign out_1_4_r = temp_b5_1_4_r;
assign out_1_4_i = temp_b5_1_4_i;
assign out_1_5_r = temp_b5_1_5_r;
assign out_1_5_i = temp_b5_1_5_i;
assign out_1_6_r = temp_b5_1_6_r;
assign out_1_6_i = temp_b5_1_6_i;
assign out_1_7_r = temp_b5_1_7_r;
assign out_1_7_i = temp_b5_1_7_i;
assign out_1_8_r = temp_b5_1_8_r;
assign out_1_8_i = temp_b5_1_8_i;
assign out_1_9_r = temp_b5_1_9_r;
assign out_1_9_i = temp_b5_1_9_i;
assign out_1_10_r = temp_b5_1_10_r;
assign out_1_10_i = temp_b5_1_10_i;
assign out_1_11_r = temp_b5_1_11_r;
assign out_1_11_i = temp_b5_1_11_i;
assign out_1_12_r = temp_b5_1_12_r;
assign out_1_12_i = temp_b5_1_12_i;
assign out_1_13_r = temp_b5_1_13_r;
assign out_1_13_i = temp_b5_1_13_i;
assign out_1_14_r = temp_b5_1_14_r;
assign out_1_14_i = temp_b5_1_14_i;
assign out_1_15_r = temp_b5_1_15_r;
assign out_1_15_i = temp_b5_1_15_i;
assign out_1_16_r = temp_b5_1_16_r;
assign out_1_16_i = temp_b5_1_16_i;
assign out_1_17_r = temp_b5_1_17_r;
assign out_1_17_i = temp_b5_1_17_i;
assign out_1_18_r = temp_b5_1_18_r;
assign out_1_18_i = temp_b5_1_18_i;
assign out_1_19_r = temp_b5_1_19_r;
assign out_1_19_i = temp_b5_1_19_i;
assign out_1_20_r = temp_b5_1_20_r;
assign out_1_20_i = temp_b5_1_20_i;
assign out_1_21_r = temp_b5_1_21_r;
assign out_1_21_i = temp_b5_1_21_i;
assign out_1_22_r = temp_b5_1_22_r;
assign out_1_22_i = temp_b5_1_22_i;
assign out_1_23_r = temp_b5_1_23_r;
assign out_1_23_i = temp_b5_1_23_i;
assign out_1_24_r = temp_b5_1_24_r;
assign out_1_24_i = temp_b5_1_24_i;
assign out_1_25_r = temp_b5_1_25_r;
assign out_1_25_i = temp_b5_1_25_i;
assign out_1_26_r = temp_b5_1_26_r;
assign out_1_26_i = temp_b5_1_26_i;
assign out_1_27_r = temp_b5_1_27_r;
assign out_1_27_i = temp_b5_1_27_i;
assign out_1_28_r = temp_b5_1_28_r;
assign out_1_28_i = temp_b5_1_28_i;
assign out_1_29_r = temp_b5_1_29_r;
assign out_1_29_i = temp_b5_1_29_i;
assign out_1_30_r = temp_b5_1_30_r;
assign out_1_30_i = temp_b5_1_30_i;
assign out_1_31_r = temp_b5_1_31_r;
assign out_1_31_i = temp_b5_1_31_i;
assign out_1_32_r = temp_b5_1_32_r;
assign out_1_32_i = temp_b5_1_32_i;
assign out_2_1_r = temp_b5_2_1_r;
assign out_2_1_i = temp_b5_2_1_i;
assign out_2_2_r = temp_b5_2_2_r;
assign out_2_2_i = temp_b5_2_2_i;
assign out_2_3_r = temp_b5_2_3_r;
assign out_2_3_i = temp_b5_2_3_i;
assign out_2_4_r = temp_b5_2_4_r;
assign out_2_4_i = temp_b5_2_4_i;
assign out_2_5_r = temp_b5_2_5_r;
assign out_2_5_i = temp_b5_2_5_i;
assign out_2_6_r = temp_b5_2_6_r;
assign out_2_6_i = temp_b5_2_6_i;
assign out_2_7_r = temp_b5_2_7_r;
assign out_2_7_i = temp_b5_2_7_i;
assign out_2_8_r = temp_b5_2_8_r;
assign out_2_8_i = temp_b5_2_8_i;
assign out_2_9_r = temp_b5_2_9_r;
assign out_2_9_i = temp_b5_2_9_i;
assign out_2_10_r = temp_b5_2_10_r;
assign out_2_10_i = temp_b5_2_10_i;
assign out_2_11_r = temp_b5_2_11_r;
assign out_2_11_i = temp_b5_2_11_i;
assign out_2_12_r = temp_b5_2_12_r;
assign out_2_12_i = temp_b5_2_12_i;
assign out_2_13_r = temp_b5_2_13_r;
assign out_2_13_i = temp_b5_2_13_i;
assign out_2_14_r = temp_b5_2_14_r;
assign out_2_14_i = temp_b5_2_14_i;
assign out_2_15_r = temp_b5_2_15_r;
assign out_2_15_i = temp_b5_2_15_i;
assign out_2_16_r = temp_b5_2_16_r;
assign out_2_16_i = temp_b5_2_16_i;
assign out_2_17_r = temp_b5_2_17_r;
assign out_2_17_i = temp_b5_2_17_i;
assign out_2_18_r = temp_b5_2_18_r;
assign out_2_18_i = temp_b5_2_18_i;
assign out_2_19_r = temp_b5_2_19_r;
assign out_2_19_i = temp_b5_2_19_i;
assign out_2_20_r = temp_b5_2_20_r;
assign out_2_20_i = temp_b5_2_20_i;
assign out_2_21_r = temp_b5_2_21_r;
assign out_2_21_i = temp_b5_2_21_i;
assign out_2_22_r = temp_b5_2_22_r;
assign out_2_22_i = temp_b5_2_22_i;
assign out_2_23_r = temp_b5_2_23_r;
assign out_2_23_i = temp_b5_2_23_i;
assign out_2_24_r = temp_b5_2_24_r;
assign out_2_24_i = temp_b5_2_24_i;
assign out_2_25_r = temp_b5_2_25_r;
assign out_2_25_i = temp_b5_2_25_i;
assign out_2_26_r = temp_b5_2_26_r;
assign out_2_26_i = temp_b5_2_26_i;
assign out_2_27_r = temp_b5_2_27_r;
assign out_2_27_i = temp_b5_2_27_i;
assign out_2_28_r = temp_b5_2_28_r;
assign out_2_28_i = temp_b5_2_28_i;
assign out_2_29_r = temp_b5_2_29_r;
assign out_2_29_i = temp_b5_2_29_i;
assign out_2_30_r = temp_b5_2_30_r;
assign out_2_30_i = temp_b5_2_30_i;
assign out_2_31_r = temp_b5_2_31_r;
assign out_2_31_i = temp_b5_2_31_i;
assign out_2_32_r = temp_b5_2_32_r;
assign out_2_32_i = temp_b5_2_32_i;
assign out_3_1_r = temp_b5_3_1_r;
assign out_3_1_i = temp_b5_3_1_i;
assign out_3_2_r = temp_b5_3_2_r;
assign out_3_2_i = temp_b5_3_2_i;
assign out_3_3_r = temp_b5_3_3_r;
assign out_3_3_i = temp_b5_3_3_i;
assign out_3_4_r = temp_b5_3_4_r;
assign out_3_4_i = temp_b5_3_4_i;
assign out_3_5_r = temp_b5_3_5_r;
assign out_3_5_i = temp_b5_3_5_i;
assign out_3_6_r = temp_b5_3_6_r;
assign out_3_6_i = temp_b5_3_6_i;
assign out_3_7_r = temp_b5_3_7_r;
assign out_3_7_i = temp_b5_3_7_i;
assign out_3_8_r = temp_b5_3_8_r;
assign out_3_8_i = temp_b5_3_8_i;
assign out_3_9_r = temp_b5_3_9_r;
assign out_3_9_i = temp_b5_3_9_i;
assign out_3_10_r = temp_b5_3_10_r;
assign out_3_10_i = temp_b5_3_10_i;
assign out_3_11_r = temp_b5_3_11_r;
assign out_3_11_i = temp_b5_3_11_i;
assign out_3_12_r = temp_b5_3_12_r;
assign out_3_12_i = temp_b5_3_12_i;
assign out_3_13_r = temp_b5_3_13_r;
assign out_3_13_i = temp_b5_3_13_i;
assign out_3_14_r = temp_b5_3_14_r;
assign out_3_14_i = temp_b5_3_14_i;
assign out_3_15_r = temp_b5_3_15_r;
assign out_3_15_i = temp_b5_3_15_i;
assign out_3_16_r = temp_b5_3_16_r;
assign out_3_16_i = temp_b5_3_16_i;
assign out_3_17_r = temp_b5_3_17_r;
assign out_3_17_i = temp_b5_3_17_i;
assign out_3_18_r = temp_b5_3_18_r;
assign out_3_18_i = temp_b5_3_18_i;
assign out_3_19_r = temp_b5_3_19_r;
assign out_3_19_i = temp_b5_3_19_i;
assign out_3_20_r = temp_b5_3_20_r;
assign out_3_20_i = temp_b5_3_20_i;
assign out_3_21_r = temp_b5_3_21_r;
assign out_3_21_i = temp_b5_3_21_i;
assign out_3_22_r = temp_b5_3_22_r;
assign out_3_22_i = temp_b5_3_22_i;
assign out_3_23_r = temp_b5_3_23_r;
assign out_3_23_i = temp_b5_3_23_i;
assign out_3_24_r = temp_b5_3_24_r;
assign out_3_24_i = temp_b5_3_24_i;
assign out_3_25_r = temp_b5_3_25_r;
assign out_3_25_i = temp_b5_3_25_i;
assign out_3_26_r = temp_b5_3_26_r;
assign out_3_26_i = temp_b5_3_26_i;
assign out_3_27_r = temp_b5_3_27_r;
assign out_3_27_i = temp_b5_3_27_i;
assign out_3_28_r = temp_b5_3_28_r;
assign out_3_28_i = temp_b5_3_28_i;
assign out_3_29_r = temp_b5_3_29_r;
assign out_3_29_i = temp_b5_3_29_i;
assign out_3_30_r = temp_b5_3_30_r;
assign out_3_30_i = temp_b5_3_30_i;
assign out_3_31_r = temp_b5_3_31_r;
assign out_3_31_i = temp_b5_3_31_i;
assign out_3_32_r = temp_b5_3_32_r;
assign out_3_32_i = temp_b5_3_32_i;
assign out_4_1_r = temp_b5_4_1_r;
assign out_4_1_i = temp_b5_4_1_i;
assign out_4_2_r = temp_b5_4_2_r;
assign out_4_2_i = temp_b5_4_2_i;
assign out_4_3_r = temp_b5_4_3_r;
assign out_4_3_i = temp_b5_4_3_i;
assign out_4_4_r = temp_b5_4_4_r;
assign out_4_4_i = temp_b5_4_4_i;
assign out_4_5_r = temp_b5_4_5_r;
assign out_4_5_i = temp_b5_4_5_i;
assign out_4_6_r = temp_b5_4_6_r;
assign out_4_6_i = temp_b5_4_6_i;
assign out_4_7_r = temp_b5_4_7_r;
assign out_4_7_i = temp_b5_4_7_i;
assign out_4_8_r = temp_b5_4_8_r;
assign out_4_8_i = temp_b5_4_8_i;
assign out_4_9_r = temp_b5_4_9_r;
assign out_4_9_i = temp_b5_4_9_i;
assign out_4_10_r = temp_b5_4_10_r;
assign out_4_10_i = temp_b5_4_10_i;
assign out_4_11_r = temp_b5_4_11_r;
assign out_4_11_i = temp_b5_4_11_i;
assign out_4_12_r = temp_b5_4_12_r;
assign out_4_12_i = temp_b5_4_12_i;
assign out_4_13_r = temp_b5_4_13_r;
assign out_4_13_i = temp_b5_4_13_i;
assign out_4_14_r = temp_b5_4_14_r;
assign out_4_14_i = temp_b5_4_14_i;
assign out_4_15_r = temp_b5_4_15_r;
assign out_4_15_i = temp_b5_4_15_i;
assign out_4_16_r = temp_b5_4_16_r;
assign out_4_16_i = temp_b5_4_16_i;
assign out_4_17_r = temp_b5_4_17_r;
assign out_4_17_i = temp_b5_4_17_i;
assign out_4_18_r = temp_b5_4_18_r;
assign out_4_18_i = temp_b5_4_18_i;
assign out_4_19_r = temp_b5_4_19_r;
assign out_4_19_i = temp_b5_4_19_i;
assign out_4_20_r = temp_b5_4_20_r;
assign out_4_20_i = temp_b5_4_20_i;
assign out_4_21_r = temp_b5_4_21_r;
assign out_4_21_i = temp_b5_4_21_i;
assign out_4_22_r = temp_b5_4_22_r;
assign out_4_22_i = temp_b5_4_22_i;
assign out_4_23_r = temp_b5_4_23_r;
assign out_4_23_i = temp_b5_4_23_i;
assign out_4_24_r = temp_b5_4_24_r;
assign out_4_24_i = temp_b5_4_24_i;
assign out_4_25_r = temp_b5_4_25_r;
assign out_4_25_i = temp_b5_4_25_i;
assign out_4_26_r = temp_b5_4_26_r;
assign out_4_26_i = temp_b5_4_26_i;
assign out_4_27_r = temp_b5_4_27_r;
assign out_4_27_i = temp_b5_4_27_i;
assign out_4_28_r = temp_b5_4_28_r;
assign out_4_28_i = temp_b5_4_28_i;
assign out_4_29_r = temp_b5_4_29_r;
assign out_4_29_i = temp_b5_4_29_i;
assign out_4_30_r = temp_b5_4_30_r;
assign out_4_30_i = temp_b5_4_30_i;
assign out_4_31_r = temp_b5_4_31_r;
assign out_4_31_i = temp_b5_4_31_i;
assign out_4_32_r = temp_b5_4_32_r;
assign out_4_32_i = temp_b5_4_32_i;
assign out_5_1_r = temp_b5_5_1_r;
assign out_5_1_i = temp_b5_5_1_i;
assign out_5_2_r = temp_b5_5_2_r;
assign out_5_2_i = temp_b5_5_2_i;
assign out_5_3_r = temp_b5_5_3_r;
assign out_5_3_i = temp_b5_5_3_i;
assign out_5_4_r = temp_b5_5_4_r;
assign out_5_4_i = temp_b5_5_4_i;
assign out_5_5_r = temp_b5_5_5_r;
assign out_5_5_i = temp_b5_5_5_i;
assign out_5_6_r = temp_b5_5_6_r;
assign out_5_6_i = temp_b5_5_6_i;
assign out_5_7_r = temp_b5_5_7_r;
assign out_5_7_i = temp_b5_5_7_i;
assign out_5_8_r = temp_b5_5_8_r;
assign out_5_8_i = temp_b5_5_8_i;
assign out_5_9_r = temp_b5_5_9_r;
assign out_5_9_i = temp_b5_5_9_i;
assign out_5_10_r = temp_b5_5_10_r;
assign out_5_10_i = temp_b5_5_10_i;
assign out_5_11_r = temp_b5_5_11_r;
assign out_5_11_i = temp_b5_5_11_i;
assign out_5_12_r = temp_b5_5_12_r;
assign out_5_12_i = temp_b5_5_12_i;
assign out_5_13_r = temp_b5_5_13_r;
assign out_5_13_i = temp_b5_5_13_i;
assign out_5_14_r = temp_b5_5_14_r;
assign out_5_14_i = temp_b5_5_14_i;
assign out_5_15_r = temp_b5_5_15_r;
assign out_5_15_i = temp_b5_5_15_i;
assign out_5_16_r = temp_b5_5_16_r;
assign out_5_16_i = temp_b5_5_16_i;
assign out_5_17_r = temp_b5_5_17_r;
assign out_5_17_i = temp_b5_5_17_i;
assign out_5_18_r = temp_b5_5_18_r;
assign out_5_18_i = temp_b5_5_18_i;
assign out_5_19_r = temp_b5_5_19_r;
assign out_5_19_i = temp_b5_5_19_i;
assign out_5_20_r = temp_b5_5_20_r;
assign out_5_20_i = temp_b5_5_20_i;
assign out_5_21_r = temp_b5_5_21_r;
assign out_5_21_i = temp_b5_5_21_i;
assign out_5_22_r = temp_b5_5_22_r;
assign out_5_22_i = temp_b5_5_22_i;
assign out_5_23_r = temp_b5_5_23_r;
assign out_5_23_i = temp_b5_5_23_i;
assign out_5_24_r = temp_b5_5_24_r;
assign out_5_24_i = temp_b5_5_24_i;
assign out_5_25_r = temp_b5_5_25_r;
assign out_5_25_i = temp_b5_5_25_i;
assign out_5_26_r = temp_b5_5_26_r;
assign out_5_26_i = temp_b5_5_26_i;
assign out_5_27_r = temp_b5_5_27_r;
assign out_5_27_i = temp_b5_5_27_i;
assign out_5_28_r = temp_b5_5_28_r;
assign out_5_28_i = temp_b5_5_28_i;
assign out_5_29_r = temp_b5_5_29_r;
assign out_5_29_i = temp_b5_5_29_i;
assign out_5_30_r = temp_b5_5_30_r;
assign out_5_30_i = temp_b5_5_30_i;
assign out_5_31_r = temp_b5_5_31_r;
assign out_5_31_i = temp_b5_5_31_i;
assign out_5_32_r = temp_b5_5_32_r;
assign out_5_32_i = temp_b5_5_32_i;
assign out_6_1_r = temp_b5_6_1_r;
assign out_6_1_i = temp_b5_6_1_i;
assign out_6_2_r = temp_b5_6_2_r;
assign out_6_2_i = temp_b5_6_2_i;
assign out_6_3_r = temp_b5_6_3_r;
assign out_6_3_i = temp_b5_6_3_i;
assign out_6_4_r = temp_b5_6_4_r;
assign out_6_4_i = temp_b5_6_4_i;
assign out_6_5_r = temp_b5_6_5_r;
assign out_6_5_i = temp_b5_6_5_i;
assign out_6_6_r = temp_b5_6_6_r;
assign out_6_6_i = temp_b5_6_6_i;
assign out_6_7_r = temp_b5_6_7_r;
assign out_6_7_i = temp_b5_6_7_i;
assign out_6_8_r = temp_b5_6_8_r;
assign out_6_8_i = temp_b5_6_8_i;
assign out_6_9_r = temp_b5_6_9_r;
assign out_6_9_i = temp_b5_6_9_i;
assign out_6_10_r = temp_b5_6_10_r;
assign out_6_10_i = temp_b5_6_10_i;
assign out_6_11_r = temp_b5_6_11_r;
assign out_6_11_i = temp_b5_6_11_i;
assign out_6_12_r = temp_b5_6_12_r;
assign out_6_12_i = temp_b5_6_12_i;
assign out_6_13_r = temp_b5_6_13_r;
assign out_6_13_i = temp_b5_6_13_i;
assign out_6_14_r = temp_b5_6_14_r;
assign out_6_14_i = temp_b5_6_14_i;
assign out_6_15_r = temp_b5_6_15_r;
assign out_6_15_i = temp_b5_6_15_i;
assign out_6_16_r = temp_b5_6_16_r;
assign out_6_16_i = temp_b5_6_16_i;
assign out_6_17_r = temp_b5_6_17_r;
assign out_6_17_i = temp_b5_6_17_i;
assign out_6_18_r = temp_b5_6_18_r;
assign out_6_18_i = temp_b5_6_18_i;
assign out_6_19_r = temp_b5_6_19_r;
assign out_6_19_i = temp_b5_6_19_i;
assign out_6_20_r = temp_b5_6_20_r;
assign out_6_20_i = temp_b5_6_20_i;
assign out_6_21_r = temp_b5_6_21_r;
assign out_6_21_i = temp_b5_6_21_i;
assign out_6_22_r = temp_b5_6_22_r;
assign out_6_22_i = temp_b5_6_22_i;
assign out_6_23_r = temp_b5_6_23_r;
assign out_6_23_i = temp_b5_6_23_i;
assign out_6_24_r = temp_b5_6_24_r;
assign out_6_24_i = temp_b5_6_24_i;
assign out_6_25_r = temp_b5_6_25_r;
assign out_6_25_i = temp_b5_6_25_i;
assign out_6_26_r = temp_b5_6_26_r;
assign out_6_26_i = temp_b5_6_26_i;
assign out_6_27_r = temp_b5_6_27_r;
assign out_6_27_i = temp_b5_6_27_i;
assign out_6_28_r = temp_b5_6_28_r;
assign out_6_28_i = temp_b5_6_28_i;
assign out_6_29_r = temp_b5_6_29_r;
assign out_6_29_i = temp_b5_6_29_i;
assign out_6_30_r = temp_b5_6_30_r;
assign out_6_30_i = temp_b5_6_30_i;
assign out_6_31_r = temp_b5_6_31_r;
assign out_6_31_i = temp_b5_6_31_i;
assign out_6_32_r = temp_b5_6_32_r;
assign out_6_32_i = temp_b5_6_32_i;
assign out_7_1_r = temp_b5_7_1_r;
assign out_7_1_i = temp_b5_7_1_i;
assign out_7_2_r = temp_b5_7_2_r;
assign out_7_2_i = temp_b5_7_2_i;
assign out_7_3_r = temp_b5_7_3_r;
assign out_7_3_i = temp_b5_7_3_i;
assign out_7_4_r = temp_b5_7_4_r;
assign out_7_4_i = temp_b5_7_4_i;
assign out_7_5_r = temp_b5_7_5_r;
assign out_7_5_i = temp_b5_7_5_i;
assign out_7_6_r = temp_b5_7_6_r;
assign out_7_6_i = temp_b5_7_6_i;
assign out_7_7_r = temp_b5_7_7_r;
assign out_7_7_i = temp_b5_7_7_i;
assign out_7_8_r = temp_b5_7_8_r;
assign out_7_8_i = temp_b5_7_8_i;
assign out_7_9_r = temp_b5_7_9_r;
assign out_7_9_i = temp_b5_7_9_i;
assign out_7_10_r = temp_b5_7_10_r;
assign out_7_10_i = temp_b5_7_10_i;
assign out_7_11_r = temp_b5_7_11_r;
assign out_7_11_i = temp_b5_7_11_i;
assign out_7_12_r = temp_b5_7_12_r;
assign out_7_12_i = temp_b5_7_12_i;
assign out_7_13_r = temp_b5_7_13_r;
assign out_7_13_i = temp_b5_7_13_i;
assign out_7_14_r = temp_b5_7_14_r;
assign out_7_14_i = temp_b5_7_14_i;
assign out_7_15_r = temp_b5_7_15_r;
assign out_7_15_i = temp_b5_7_15_i;
assign out_7_16_r = temp_b5_7_16_r;
assign out_7_16_i = temp_b5_7_16_i;
assign out_7_17_r = temp_b5_7_17_r;
assign out_7_17_i = temp_b5_7_17_i;
assign out_7_18_r = temp_b5_7_18_r;
assign out_7_18_i = temp_b5_7_18_i;
assign out_7_19_r = temp_b5_7_19_r;
assign out_7_19_i = temp_b5_7_19_i;
assign out_7_20_r = temp_b5_7_20_r;
assign out_7_20_i = temp_b5_7_20_i;
assign out_7_21_r = temp_b5_7_21_r;
assign out_7_21_i = temp_b5_7_21_i;
assign out_7_22_r = temp_b5_7_22_r;
assign out_7_22_i = temp_b5_7_22_i;
assign out_7_23_r = temp_b5_7_23_r;
assign out_7_23_i = temp_b5_7_23_i;
assign out_7_24_r = temp_b5_7_24_r;
assign out_7_24_i = temp_b5_7_24_i;
assign out_7_25_r = temp_b5_7_25_r;
assign out_7_25_i = temp_b5_7_25_i;
assign out_7_26_r = temp_b5_7_26_r;
assign out_7_26_i = temp_b5_7_26_i;
assign out_7_27_r = temp_b5_7_27_r;
assign out_7_27_i = temp_b5_7_27_i;
assign out_7_28_r = temp_b5_7_28_r;
assign out_7_28_i = temp_b5_7_28_i;
assign out_7_29_r = temp_b5_7_29_r;
assign out_7_29_i = temp_b5_7_29_i;
assign out_7_30_r = temp_b5_7_30_r;
assign out_7_30_i = temp_b5_7_30_i;
assign out_7_31_r = temp_b5_7_31_r;
assign out_7_31_i = temp_b5_7_31_i;
assign out_7_32_r = temp_b5_7_32_r;
assign out_7_32_i = temp_b5_7_32_i;
assign out_8_1_r = temp_b5_8_1_r;
assign out_8_1_i = temp_b5_8_1_i;
assign out_8_2_r = temp_b5_8_2_r;
assign out_8_2_i = temp_b5_8_2_i;
assign out_8_3_r = temp_b5_8_3_r;
assign out_8_3_i = temp_b5_8_3_i;
assign out_8_4_r = temp_b5_8_4_r;
assign out_8_4_i = temp_b5_8_4_i;
assign out_8_5_r = temp_b5_8_5_r;
assign out_8_5_i = temp_b5_8_5_i;
assign out_8_6_r = temp_b5_8_6_r;
assign out_8_6_i = temp_b5_8_6_i;
assign out_8_7_r = temp_b5_8_7_r;
assign out_8_7_i = temp_b5_8_7_i;
assign out_8_8_r = temp_b5_8_8_r;
assign out_8_8_i = temp_b5_8_8_i;
assign out_8_9_r = temp_b5_8_9_r;
assign out_8_9_i = temp_b5_8_9_i;
assign out_8_10_r = temp_b5_8_10_r;
assign out_8_10_i = temp_b5_8_10_i;
assign out_8_11_r = temp_b5_8_11_r;
assign out_8_11_i = temp_b5_8_11_i;
assign out_8_12_r = temp_b5_8_12_r;
assign out_8_12_i = temp_b5_8_12_i;
assign out_8_13_r = temp_b5_8_13_r;
assign out_8_13_i = temp_b5_8_13_i;
assign out_8_14_r = temp_b5_8_14_r;
assign out_8_14_i = temp_b5_8_14_i;
assign out_8_15_r = temp_b5_8_15_r;
assign out_8_15_i = temp_b5_8_15_i;
assign out_8_16_r = temp_b5_8_16_r;
assign out_8_16_i = temp_b5_8_16_i;
assign out_8_17_r = temp_b5_8_17_r;
assign out_8_17_i = temp_b5_8_17_i;
assign out_8_18_r = temp_b5_8_18_r;
assign out_8_18_i = temp_b5_8_18_i;
assign out_8_19_r = temp_b5_8_19_r;
assign out_8_19_i = temp_b5_8_19_i;
assign out_8_20_r = temp_b5_8_20_r;
assign out_8_20_i = temp_b5_8_20_i;
assign out_8_21_r = temp_b5_8_21_r;
assign out_8_21_i = temp_b5_8_21_i;
assign out_8_22_r = temp_b5_8_22_r;
assign out_8_22_i = temp_b5_8_22_i;
assign out_8_23_r = temp_b5_8_23_r;
assign out_8_23_i = temp_b5_8_23_i;
assign out_8_24_r = temp_b5_8_24_r;
assign out_8_24_i = temp_b5_8_24_i;
assign out_8_25_r = temp_b5_8_25_r;
assign out_8_25_i = temp_b5_8_25_i;
assign out_8_26_r = temp_b5_8_26_r;
assign out_8_26_i = temp_b5_8_26_i;
assign out_8_27_r = temp_b5_8_27_r;
assign out_8_27_i = temp_b5_8_27_i;
assign out_8_28_r = temp_b5_8_28_r;
assign out_8_28_i = temp_b5_8_28_i;
assign out_8_29_r = temp_b5_8_29_r;
assign out_8_29_i = temp_b5_8_29_i;
assign out_8_30_r = temp_b5_8_30_r;
assign out_8_30_i = temp_b5_8_30_i;
assign out_8_31_r = temp_b5_8_31_r;
assign out_8_31_i = temp_b5_8_31_i;
assign out_8_32_r = temp_b5_8_32_r;
assign out_8_32_i = temp_b5_8_32_i;
assign out_9_1_r = temp_b5_9_1_r;
assign out_9_1_i = temp_b5_9_1_i;
assign out_9_2_r = temp_b5_9_2_r;
assign out_9_2_i = temp_b5_9_2_i;
assign out_9_3_r = temp_b5_9_3_r;
assign out_9_3_i = temp_b5_9_3_i;
assign out_9_4_r = temp_b5_9_4_r;
assign out_9_4_i = temp_b5_9_4_i;
assign out_9_5_r = temp_b5_9_5_r;
assign out_9_5_i = temp_b5_9_5_i;
assign out_9_6_r = temp_b5_9_6_r;
assign out_9_6_i = temp_b5_9_6_i;
assign out_9_7_r = temp_b5_9_7_r;
assign out_9_7_i = temp_b5_9_7_i;
assign out_9_8_r = temp_b5_9_8_r;
assign out_9_8_i = temp_b5_9_8_i;
assign out_9_9_r = temp_b5_9_9_r;
assign out_9_9_i = temp_b5_9_9_i;
assign out_9_10_r = temp_b5_9_10_r;
assign out_9_10_i = temp_b5_9_10_i;
assign out_9_11_r = temp_b5_9_11_r;
assign out_9_11_i = temp_b5_9_11_i;
assign out_9_12_r = temp_b5_9_12_r;
assign out_9_12_i = temp_b5_9_12_i;
assign out_9_13_r = temp_b5_9_13_r;
assign out_9_13_i = temp_b5_9_13_i;
assign out_9_14_r = temp_b5_9_14_r;
assign out_9_14_i = temp_b5_9_14_i;
assign out_9_15_r = temp_b5_9_15_r;
assign out_9_15_i = temp_b5_9_15_i;
assign out_9_16_r = temp_b5_9_16_r;
assign out_9_16_i = temp_b5_9_16_i;
assign out_9_17_r = temp_b5_9_17_r;
assign out_9_17_i = temp_b5_9_17_i;
assign out_9_18_r = temp_b5_9_18_r;
assign out_9_18_i = temp_b5_9_18_i;
assign out_9_19_r = temp_b5_9_19_r;
assign out_9_19_i = temp_b5_9_19_i;
assign out_9_20_r = temp_b5_9_20_r;
assign out_9_20_i = temp_b5_9_20_i;
assign out_9_21_r = temp_b5_9_21_r;
assign out_9_21_i = temp_b5_9_21_i;
assign out_9_22_r = temp_b5_9_22_r;
assign out_9_22_i = temp_b5_9_22_i;
assign out_9_23_r = temp_b5_9_23_r;
assign out_9_23_i = temp_b5_9_23_i;
assign out_9_24_r = temp_b5_9_24_r;
assign out_9_24_i = temp_b5_9_24_i;
assign out_9_25_r = temp_b5_9_25_r;
assign out_9_25_i = temp_b5_9_25_i;
assign out_9_26_r = temp_b5_9_26_r;
assign out_9_26_i = temp_b5_9_26_i;
assign out_9_27_r = temp_b5_9_27_r;
assign out_9_27_i = temp_b5_9_27_i;
assign out_9_28_r = temp_b5_9_28_r;
assign out_9_28_i = temp_b5_9_28_i;
assign out_9_29_r = temp_b5_9_29_r;
assign out_9_29_i = temp_b5_9_29_i;
assign out_9_30_r = temp_b5_9_30_r;
assign out_9_30_i = temp_b5_9_30_i;
assign out_9_31_r = temp_b5_9_31_r;
assign out_9_31_i = temp_b5_9_31_i;
assign out_9_32_r = temp_b5_9_32_r;
assign out_9_32_i = temp_b5_9_32_i;
assign out_10_1_r = temp_b5_10_1_r;
assign out_10_1_i = temp_b5_10_1_i;
assign out_10_2_r = temp_b5_10_2_r;
assign out_10_2_i = temp_b5_10_2_i;
assign out_10_3_r = temp_b5_10_3_r;
assign out_10_3_i = temp_b5_10_3_i;
assign out_10_4_r = temp_b5_10_4_r;
assign out_10_4_i = temp_b5_10_4_i;
assign out_10_5_r = temp_b5_10_5_r;
assign out_10_5_i = temp_b5_10_5_i;
assign out_10_6_r = temp_b5_10_6_r;
assign out_10_6_i = temp_b5_10_6_i;
assign out_10_7_r = temp_b5_10_7_r;
assign out_10_7_i = temp_b5_10_7_i;
assign out_10_8_r = temp_b5_10_8_r;
assign out_10_8_i = temp_b5_10_8_i;
assign out_10_9_r = temp_b5_10_9_r;
assign out_10_9_i = temp_b5_10_9_i;
assign out_10_10_r = temp_b5_10_10_r;
assign out_10_10_i = temp_b5_10_10_i;
assign out_10_11_r = temp_b5_10_11_r;
assign out_10_11_i = temp_b5_10_11_i;
assign out_10_12_r = temp_b5_10_12_r;
assign out_10_12_i = temp_b5_10_12_i;
assign out_10_13_r = temp_b5_10_13_r;
assign out_10_13_i = temp_b5_10_13_i;
assign out_10_14_r = temp_b5_10_14_r;
assign out_10_14_i = temp_b5_10_14_i;
assign out_10_15_r = temp_b5_10_15_r;
assign out_10_15_i = temp_b5_10_15_i;
assign out_10_16_r = temp_b5_10_16_r;
assign out_10_16_i = temp_b5_10_16_i;
assign out_10_17_r = temp_b5_10_17_r;
assign out_10_17_i = temp_b5_10_17_i;
assign out_10_18_r = temp_b5_10_18_r;
assign out_10_18_i = temp_b5_10_18_i;
assign out_10_19_r = temp_b5_10_19_r;
assign out_10_19_i = temp_b5_10_19_i;
assign out_10_20_r = temp_b5_10_20_r;
assign out_10_20_i = temp_b5_10_20_i;
assign out_10_21_r = temp_b5_10_21_r;
assign out_10_21_i = temp_b5_10_21_i;
assign out_10_22_r = temp_b5_10_22_r;
assign out_10_22_i = temp_b5_10_22_i;
assign out_10_23_r = temp_b5_10_23_r;
assign out_10_23_i = temp_b5_10_23_i;
assign out_10_24_r = temp_b5_10_24_r;
assign out_10_24_i = temp_b5_10_24_i;
assign out_10_25_r = temp_b5_10_25_r;
assign out_10_25_i = temp_b5_10_25_i;
assign out_10_26_r = temp_b5_10_26_r;
assign out_10_26_i = temp_b5_10_26_i;
assign out_10_27_r = temp_b5_10_27_r;
assign out_10_27_i = temp_b5_10_27_i;
assign out_10_28_r = temp_b5_10_28_r;
assign out_10_28_i = temp_b5_10_28_i;
assign out_10_29_r = temp_b5_10_29_r;
assign out_10_29_i = temp_b5_10_29_i;
assign out_10_30_r = temp_b5_10_30_r;
assign out_10_30_i = temp_b5_10_30_i;
assign out_10_31_r = temp_b5_10_31_r;
assign out_10_31_i = temp_b5_10_31_i;
assign out_10_32_r = temp_b5_10_32_r;
assign out_10_32_i = temp_b5_10_32_i;
assign out_11_1_r = temp_b5_11_1_r;
assign out_11_1_i = temp_b5_11_1_i;
assign out_11_2_r = temp_b5_11_2_r;
assign out_11_2_i = temp_b5_11_2_i;
assign out_11_3_r = temp_b5_11_3_r;
assign out_11_3_i = temp_b5_11_3_i;
assign out_11_4_r = temp_b5_11_4_r;
assign out_11_4_i = temp_b5_11_4_i;
assign out_11_5_r = temp_b5_11_5_r;
assign out_11_5_i = temp_b5_11_5_i;
assign out_11_6_r = temp_b5_11_6_r;
assign out_11_6_i = temp_b5_11_6_i;
assign out_11_7_r = temp_b5_11_7_r;
assign out_11_7_i = temp_b5_11_7_i;
assign out_11_8_r = temp_b5_11_8_r;
assign out_11_8_i = temp_b5_11_8_i;
assign out_11_9_r = temp_b5_11_9_r;
assign out_11_9_i = temp_b5_11_9_i;
assign out_11_10_r = temp_b5_11_10_r;
assign out_11_10_i = temp_b5_11_10_i;
assign out_11_11_r = temp_b5_11_11_r;
assign out_11_11_i = temp_b5_11_11_i;
assign out_11_12_r = temp_b5_11_12_r;
assign out_11_12_i = temp_b5_11_12_i;
assign out_11_13_r = temp_b5_11_13_r;
assign out_11_13_i = temp_b5_11_13_i;
assign out_11_14_r = temp_b5_11_14_r;
assign out_11_14_i = temp_b5_11_14_i;
assign out_11_15_r = temp_b5_11_15_r;
assign out_11_15_i = temp_b5_11_15_i;
assign out_11_16_r = temp_b5_11_16_r;
assign out_11_16_i = temp_b5_11_16_i;
assign out_11_17_r = temp_b5_11_17_r;
assign out_11_17_i = temp_b5_11_17_i;
assign out_11_18_r = temp_b5_11_18_r;
assign out_11_18_i = temp_b5_11_18_i;
assign out_11_19_r = temp_b5_11_19_r;
assign out_11_19_i = temp_b5_11_19_i;
assign out_11_20_r = temp_b5_11_20_r;
assign out_11_20_i = temp_b5_11_20_i;
assign out_11_21_r = temp_b5_11_21_r;
assign out_11_21_i = temp_b5_11_21_i;
assign out_11_22_r = temp_b5_11_22_r;
assign out_11_22_i = temp_b5_11_22_i;
assign out_11_23_r = temp_b5_11_23_r;
assign out_11_23_i = temp_b5_11_23_i;
assign out_11_24_r = temp_b5_11_24_r;
assign out_11_24_i = temp_b5_11_24_i;
assign out_11_25_r = temp_b5_11_25_r;
assign out_11_25_i = temp_b5_11_25_i;
assign out_11_26_r = temp_b5_11_26_r;
assign out_11_26_i = temp_b5_11_26_i;
assign out_11_27_r = temp_b5_11_27_r;
assign out_11_27_i = temp_b5_11_27_i;
assign out_11_28_r = temp_b5_11_28_r;
assign out_11_28_i = temp_b5_11_28_i;
assign out_11_29_r = temp_b5_11_29_r;
assign out_11_29_i = temp_b5_11_29_i;
assign out_11_30_r = temp_b5_11_30_r;
assign out_11_30_i = temp_b5_11_30_i;
assign out_11_31_r = temp_b5_11_31_r;
assign out_11_31_i = temp_b5_11_31_i;
assign out_11_32_r = temp_b5_11_32_r;
assign out_11_32_i = temp_b5_11_32_i;
assign out_12_1_r = temp_b5_12_1_r;
assign out_12_1_i = temp_b5_12_1_i;
assign out_12_2_r = temp_b5_12_2_r;
assign out_12_2_i = temp_b5_12_2_i;
assign out_12_3_r = temp_b5_12_3_r;
assign out_12_3_i = temp_b5_12_3_i;
assign out_12_4_r = temp_b5_12_4_r;
assign out_12_4_i = temp_b5_12_4_i;
assign out_12_5_r = temp_b5_12_5_r;
assign out_12_5_i = temp_b5_12_5_i;
assign out_12_6_r = temp_b5_12_6_r;
assign out_12_6_i = temp_b5_12_6_i;
assign out_12_7_r = temp_b5_12_7_r;
assign out_12_7_i = temp_b5_12_7_i;
assign out_12_8_r = temp_b5_12_8_r;
assign out_12_8_i = temp_b5_12_8_i;
assign out_12_9_r = temp_b5_12_9_r;
assign out_12_9_i = temp_b5_12_9_i;
assign out_12_10_r = temp_b5_12_10_r;
assign out_12_10_i = temp_b5_12_10_i;
assign out_12_11_r = temp_b5_12_11_r;
assign out_12_11_i = temp_b5_12_11_i;
assign out_12_12_r = temp_b5_12_12_r;
assign out_12_12_i = temp_b5_12_12_i;
assign out_12_13_r = temp_b5_12_13_r;
assign out_12_13_i = temp_b5_12_13_i;
assign out_12_14_r = temp_b5_12_14_r;
assign out_12_14_i = temp_b5_12_14_i;
assign out_12_15_r = temp_b5_12_15_r;
assign out_12_15_i = temp_b5_12_15_i;
assign out_12_16_r = temp_b5_12_16_r;
assign out_12_16_i = temp_b5_12_16_i;
assign out_12_17_r = temp_b5_12_17_r;
assign out_12_17_i = temp_b5_12_17_i;
assign out_12_18_r = temp_b5_12_18_r;
assign out_12_18_i = temp_b5_12_18_i;
assign out_12_19_r = temp_b5_12_19_r;
assign out_12_19_i = temp_b5_12_19_i;
assign out_12_20_r = temp_b5_12_20_r;
assign out_12_20_i = temp_b5_12_20_i;
assign out_12_21_r = temp_b5_12_21_r;
assign out_12_21_i = temp_b5_12_21_i;
assign out_12_22_r = temp_b5_12_22_r;
assign out_12_22_i = temp_b5_12_22_i;
assign out_12_23_r = temp_b5_12_23_r;
assign out_12_23_i = temp_b5_12_23_i;
assign out_12_24_r = temp_b5_12_24_r;
assign out_12_24_i = temp_b5_12_24_i;
assign out_12_25_r = temp_b5_12_25_r;
assign out_12_25_i = temp_b5_12_25_i;
assign out_12_26_r = temp_b5_12_26_r;
assign out_12_26_i = temp_b5_12_26_i;
assign out_12_27_r = temp_b5_12_27_r;
assign out_12_27_i = temp_b5_12_27_i;
assign out_12_28_r = temp_b5_12_28_r;
assign out_12_28_i = temp_b5_12_28_i;
assign out_12_29_r = temp_b5_12_29_r;
assign out_12_29_i = temp_b5_12_29_i;
assign out_12_30_r = temp_b5_12_30_r;
assign out_12_30_i = temp_b5_12_30_i;
assign out_12_31_r = temp_b5_12_31_r;
assign out_12_31_i = temp_b5_12_31_i;
assign out_12_32_r = temp_b5_12_32_r;
assign out_12_32_i = temp_b5_12_32_i;
assign out_13_1_r = temp_b5_13_1_r;
assign out_13_1_i = temp_b5_13_1_i;
assign out_13_2_r = temp_b5_13_2_r;
assign out_13_2_i = temp_b5_13_2_i;
assign out_13_3_r = temp_b5_13_3_r;
assign out_13_3_i = temp_b5_13_3_i;
assign out_13_4_r = temp_b5_13_4_r;
assign out_13_4_i = temp_b5_13_4_i;
assign out_13_5_r = temp_b5_13_5_r;
assign out_13_5_i = temp_b5_13_5_i;
assign out_13_6_r = temp_b5_13_6_r;
assign out_13_6_i = temp_b5_13_6_i;
assign out_13_7_r = temp_b5_13_7_r;
assign out_13_7_i = temp_b5_13_7_i;
assign out_13_8_r = temp_b5_13_8_r;
assign out_13_8_i = temp_b5_13_8_i;
assign out_13_9_r = temp_b5_13_9_r;
assign out_13_9_i = temp_b5_13_9_i;
assign out_13_10_r = temp_b5_13_10_r;
assign out_13_10_i = temp_b5_13_10_i;
assign out_13_11_r = temp_b5_13_11_r;
assign out_13_11_i = temp_b5_13_11_i;
assign out_13_12_r = temp_b5_13_12_r;
assign out_13_12_i = temp_b5_13_12_i;
assign out_13_13_r = temp_b5_13_13_r;
assign out_13_13_i = temp_b5_13_13_i;
assign out_13_14_r = temp_b5_13_14_r;
assign out_13_14_i = temp_b5_13_14_i;
assign out_13_15_r = temp_b5_13_15_r;
assign out_13_15_i = temp_b5_13_15_i;
assign out_13_16_r = temp_b5_13_16_r;
assign out_13_16_i = temp_b5_13_16_i;
assign out_13_17_r = temp_b5_13_17_r;
assign out_13_17_i = temp_b5_13_17_i;
assign out_13_18_r = temp_b5_13_18_r;
assign out_13_18_i = temp_b5_13_18_i;
assign out_13_19_r = temp_b5_13_19_r;
assign out_13_19_i = temp_b5_13_19_i;
assign out_13_20_r = temp_b5_13_20_r;
assign out_13_20_i = temp_b5_13_20_i;
assign out_13_21_r = temp_b5_13_21_r;
assign out_13_21_i = temp_b5_13_21_i;
assign out_13_22_r = temp_b5_13_22_r;
assign out_13_22_i = temp_b5_13_22_i;
assign out_13_23_r = temp_b5_13_23_r;
assign out_13_23_i = temp_b5_13_23_i;
assign out_13_24_r = temp_b5_13_24_r;
assign out_13_24_i = temp_b5_13_24_i;
assign out_13_25_r = temp_b5_13_25_r;
assign out_13_25_i = temp_b5_13_25_i;
assign out_13_26_r = temp_b5_13_26_r;
assign out_13_26_i = temp_b5_13_26_i;
assign out_13_27_r = temp_b5_13_27_r;
assign out_13_27_i = temp_b5_13_27_i;
assign out_13_28_r = temp_b5_13_28_r;
assign out_13_28_i = temp_b5_13_28_i;
assign out_13_29_r = temp_b5_13_29_r;
assign out_13_29_i = temp_b5_13_29_i;
assign out_13_30_r = temp_b5_13_30_r;
assign out_13_30_i = temp_b5_13_30_i;
assign out_13_31_r = temp_b5_13_31_r;
assign out_13_31_i = temp_b5_13_31_i;
assign out_13_32_r = temp_b5_13_32_r;
assign out_13_32_i = temp_b5_13_32_i;
assign out_14_1_r = temp_b5_14_1_r;
assign out_14_1_i = temp_b5_14_1_i;
assign out_14_2_r = temp_b5_14_2_r;
assign out_14_2_i = temp_b5_14_2_i;
assign out_14_3_r = temp_b5_14_3_r;
assign out_14_3_i = temp_b5_14_3_i;
assign out_14_4_r = temp_b5_14_4_r;
assign out_14_4_i = temp_b5_14_4_i;
assign out_14_5_r = temp_b5_14_5_r;
assign out_14_5_i = temp_b5_14_5_i;
assign out_14_6_r = temp_b5_14_6_r;
assign out_14_6_i = temp_b5_14_6_i;
assign out_14_7_r = temp_b5_14_7_r;
assign out_14_7_i = temp_b5_14_7_i;
assign out_14_8_r = temp_b5_14_8_r;
assign out_14_8_i = temp_b5_14_8_i;
assign out_14_9_r = temp_b5_14_9_r;
assign out_14_9_i = temp_b5_14_9_i;
assign out_14_10_r = temp_b5_14_10_r;
assign out_14_10_i = temp_b5_14_10_i;
assign out_14_11_r = temp_b5_14_11_r;
assign out_14_11_i = temp_b5_14_11_i;
assign out_14_12_r = temp_b5_14_12_r;
assign out_14_12_i = temp_b5_14_12_i;
assign out_14_13_r = temp_b5_14_13_r;
assign out_14_13_i = temp_b5_14_13_i;
assign out_14_14_r = temp_b5_14_14_r;
assign out_14_14_i = temp_b5_14_14_i;
assign out_14_15_r = temp_b5_14_15_r;
assign out_14_15_i = temp_b5_14_15_i;
assign out_14_16_r = temp_b5_14_16_r;
assign out_14_16_i = temp_b5_14_16_i;
assign out_14_17_r = temp_b5_14_17_r;
assign out_14_17_i = temp_b5_14_17_i;
assign out_14_18_r = temp_b5_14_18_r;
assign out_14_18_i = temp_b5_14_18_i;
assign out_14_19_r = temp_b5_14_19_r;
assign out_14_19_i = temp_b5_14_19_i;
assign out_14_20_r = temp_b5_14_20_r;
assign out_14_20_i = temp_b5_14_20_i;
assign out_14_21_r = temp_b5_14_21_r;
assign out_14_21_i = temp_b5_14_21_i;
assign out_14_22_r = temp_b5_14_22_r;
assign out_14_22_i = temp_b5_14_22_i;
assign out_14_23_r = temp_b5_14_23_r;
assign out_14_23_i = temp_b5_14_23_i;
assign out_14_24_r = temp_b5_14_24_r;
assign out_14_24_i = temp_b5_14_24_i;
assign out_14_25_r = temp_b5_14_25_r;
assign out_14_25_i = temp_b5_14_25_i;
assign out_14_26_r = temp_b5_14_26_r;
assign out_14_26_i = temp_b5_14_26_i;
assign out_14_27_r = temp_b5_14_27_r;
assign out_14_27_i = temp_b5_14_27_i;
assign out_14_28_r = temp_b5_14_28_r;
assign out_14_28_i = temp_b5_14_28_i;
assign out_14_29_r = temp_b5_14_29_r;
assign out_14_29_i = temp_b5_14_29_i;
assign out_14_30_r = temp_b5_14_30_r;
assign out_14_30_i = temp_b5_14_30_i;
assign out_14_31_r = temp_b5_14_31_r;
assign out_14_31_i = temp_b5_14_31_i;
assign out_14_32_r = temp_b5_14_32_r;
assign out_14_32_i = temp_b5_14_32_i;
assign out_15_1_r = temp_b5_15_1_r;
assign out_15_1_i = temp_b5_15_1_i;
assign out_15_2_r = temp_b5_15_2_r;
assign out_15_2_i = temp_b5_15_2_i;
assign out_15_3_r = temp_b5_15_3_r;
assign out_15_3_i = temp_b5_15_3_i;
assign out_15_4_r = temp_b5_15_4_r;
assign out_15_4_i = temp_b5_15_4_i;
assign out_15_5_r = temp_b5_15_5_r;
assign out_15_5_i = temp_b5_15_5_i;
assign out_15_6_r = temp_b5_15_6_r;
assign out_15_6_i = temp_b5_15_6_i;
assign out_15_7_r = temp_b5_15_7_r;
assign out_15_7_i = temp_b5_15_7_i;
assign out_15_8_r = temp_b5_15_8_r;
assign out_15_8_i = temp_b5_15_8_i;
assign out_15_9_r = temp_b5_15_9_r;
assign out_15_9_i = temp_b5_15_9_i;
assign out_15_10_r = temp_b5_15_10_r;
assign out_15_10_i = temp_b5_15_10_i;
assign out_15_11_r = temp_b5_15_11_r;
assign out_15_11_i = temp_b5_15_11_i;
assign out_15_12_r = temp_b5_15_12_r;
assign out_15_12_i = temp_b5_15_12_i;
assign out_15_13_r = temp_b5_15_13_r;
assign out_15_13_i = temp_b5_15_13_i;
assign out_15_14_r = temp_b5_15_14_r;
assign out_15_14_i = temp_b5_15_14_i;
assign out_15_15_r = temp_b5_15_15_r;
assign out_15_15_i = temp_b5_15_15_i;
assign out_15_16_r = temp_b5_15_16_r;
assign out_15_16_i = temp_b5_15_16_i;
assign out_15_17_r = temp_b5_15_17_r;
assign out_15_17_i = temp_b5_15_17_i;
assign out_15_18_r = temp_b5_15_18_r;
assign out_15_18_i = temp_b5_15_18_i;
assign out_15_19_r = temp_b5_15_19_r;
assign out_15_19_i = temp_b5_15_19_i;
assign out_15_20_r = temp_b5_15_20_r;
assign out_15_20_i = temp_b5_15_20_i;
assign out_15_21_r = temp_b5_15_21_r;
assign out_15_21_i = temp_b5_15_21_i;
assign out_15_22_r = temp_b5_15_22_r;
assign out_15_22_i = temp_b5_15_22_i;
assign out_15_23_r = temp_b5_15_23_r;
assign out_15_23_i = temp_b5_15_23_i;
assign out_15_24_r = temp_b5_15_24_r;
assign out_15_24_i = temp_b5_15_24_i;
assign out_15_25_r = temp_b5_15_25_r;
assign out_15_25_i = temp_b5_15_25_i;
assign out_15_26_r = temp_b5_15_26_r;
assign out_15_26_i = temp_b5_15_26_i;
assign out_15_27_r = temp_b5_15_27_r;
assign out_15_27_i = temp_b5_15_27_i;
assign out_15_28_r = temp_b5_15_28_r;
assign out_15_28_i = temp_b5_15_28_i;
assign out_15_29_r = temp_b5_15_29_r;
assign out_15_29_i = temp_b5_15_29_i;
assign out_15_30_r = temp_b5_15_30_r;
assign out_15_30_i = temp_b5_15_30_i;
assign out_15_31_r = temp_b5_15_31_r;
assign out_15_31_i = temp_b5_15_31_i;
assign out_15_32_r = temp_b5_15_32_r;
assign out_15_32_i = temp_b5_15_32_i;
assign out_16_1_r = temp_b5_16_1_r;
assign out_16_1_i = temp_b5_16_1_i;
assign out_16_2_r = temp_b5_16_2_r;
assign out_16_2_i = temp_b5_16_2_i;
assign out_16_3_r = temp_b5_16_3_r;
assign out_16_3_i = temp_b5_16_3_i;
assign out_16_4_r = temp_b5_16_4_r;
assign out_16_4_i = temp_b5_16_4_i;
assign out_16_5_r = temp_b5_16_5_r;
assign out_16_5_i = temp_b5_16_5_i;
assign out_16_6_r = temp_b5_16_6_r;
assign out_16_6_i = temp_b5_16_6_i;
assign out_16_7_r = temp_b5_16_7_r;
assign out_16_7_i = temp_b5_16_7_i;
assign out_16_8_r = temp_b5_16_8_r;
assign out_16_8_i = temp_b5_16_8_i;
assign out_16_9_r = temp_b5_16_9_r;
assign out_16_9_i = temp_b5_16_9_i;
assign out_16_10_r = temp_b5_16_10_r;
assign out_16_10_i = temp_b5_16_10_i;
assign out_16_11_r = temp_b5_16_11_r;
assign out_16_11_i = temp_b5_16_11_i;
assign out_16_12_r = temp_b5_16_12_r;
assign out_16_12_i = temp_b5_16_12_i;
assign out_16_13_r = temp_b5_16_13_r;
assign out_16_13_i = temp_b5_16_13_i;
assign out_16_14_r = temp_b5_16_14_r;
assign out_16_14_i = temp_b5_16_14_i;
assign out_16_15_r = temp_b5_16_15_r;
assign out_16_15_i = temp_b5_16_15_i;
assign out_16_16_r = temp_b5_16_16_r;
assign out_16_16_i = temp_b5_16_16_i;
assign out_16_17_r = temp_b5_16_17_r;
assign out_16_17_i = temp_b5_16_17_i;
assign out_16_18_r = temp_b5_16_18_r;
assign out_16_18_i = temp_b5_16_18_i;
assign out_16_19_r = temp_b5_16_19_r;
assign out_16_19_i = temp_b5_16_19_i;
assign out_16_20_r = temp_b5_16_20_r;
assign out_16_20_i = temp_b5_16_20_i;
assign out_16_21_r = temp_b5_16_21_r;
assign out_16_21_i = temp_b5_16_21_i;
assign out_16_22_r = temp_b5_16_22_r;
assign out_16_22_i = temp_b5_16_22_i;
assign out_16_23_r = temp_b5_16_23_r;
assign out_16_23_i = temp_b5_16_23_i;
assign out_16_24_r = temp_b5_16_24_r;
assign out_16_24_i = temp_b5_16_24_i;
assign out_16_25_r = temp_b5_16_25_r;
assign out_16_25_i = temp_b5_16_25_i;
assign out_16_26_r = temp_b5_16_26_r;
assign out_16_26_i = temp_b5_16_26_i;
assign out_16_27_r = temp_b5_16_27_r;
assign out_16_27_i = temp_b5_16_27_i;
assign out_16_28_r = temp_b5_16_28_r;
assign out_16_28_i = temp_b5_16_28_i;
assign out_16_29_r = temp_b5_16_29_r;
assign out_16_29_i = temp_b5_16_29_i;
assign out_16_30_r = temp_b5_16_30_r;
assign out_16_30_i = temp_b5_16_30_i;
assign out_16_31_r = temp_b5_16_31_r;
assign out_16_31_i = temp_b5_16_31_i;
assign out_16_32_r = temp_b5_16_32_r;
assign out_16_32_i = temp_b5_16_32_i;
assign out_17_1_r = temp_b5_17_1_r;
assign out_17_1_i = temp_b5_17_1_i;
assign out_17_2_r = temp_b5_17_2_r;
assign out_17_2_i = temp_b5_17_2_i;
assign out_17_3_r = temp_b5_17_3_r;
assign out_17_3_i = temp_b5_17_3_i;
assign out_17_4_r = temp_b5_17_4_r;
assign out_17_4_i = temp_b5_17_4_i;
assign out_17_5_r = temp_b5_17_5_r;
assign out_17_5_i = temp_b5_17_5_i;
assign out_17_6_r = temp_b5_17_6_r;
assign out_17_6_i = temp_b5_17_6_i;
assign out_17_7_r = temp_b5_17_7_r;
assign out_17_7_i = temp_b5_17_7_i;
assign out_17_8_r = temp_b5_17_8_r;
assign out_17_8_i = temp_b5_17_8_i;
assign out_17_9_r = temp_b5_17_9_r;
assign out_17_9_i = temp_b5_17_9_i;
assign out_17_10_r = temp_b5_17_10_r;
assign out_17_10_i = temp_b5_17_10_i;
assign out_17_11_r = temp_b5_17_11_r;
assign out_17_11_i = temp_b5_17_11_i;
assign out_17_12_r = temp_b5_17_12_r;
assign out_17_12_i = temp_b5_17_12_i;
assign out_17_13_r = temp_b5_17_13_r;
assign out_17_13_i = temp_b5_17_13_i;
assign out_17_14_r = temp_b5_17_14_r;
assign out_17_14_i = temp_b5_17_14_i;
assign out_17_15_r = temp_b5_17_15_r;
assign out_17_15_i = temp_b5_17_15_i;
assign out_17_16_r = temp_b5_17_16_r;
assign out_17_16_i = temp_b5_17_16_i;
assign out_17_17_r = temp_b5_17_17_r;
assign out_17_17_i = temp_b5_17_17_i;
assign out_17_18_r = temp_b5_17_18_r;
assign out_17_18_i = temp_b5_17_18_i;
assign out_17_19_r = temp_b5_17_19_r;
assign out_17_19_i = temp_b5_17_19_i;
assign out_17_20_r = temp_b5_17_20_r;
assign out_17_20_i = temp_b5_17_20_i;
assign out_17_21_r = temp_b5_17_21_r;
assign out_17_21_i = temp_b5_17_21_i;
assign out_17_22_r = temp_b5_17_22_r;
assign out_17_22_i = temp_b5_17_22_i;
assign out_17_23_r = temp_b5_17_23_r;
assign out_17_23_i = temp_b5_17_23_i;
assign out_17_24_r = temp_b5_17_24_r;
assign out_17_24_i = temp_b5_17_24_i;
assign out_17_25_r = temp_b5_17_25_r;
assign out_17_25_i = temp_b5_17_25_i;
assign out_17_26_r = temp_b5_17_26_r;
assign out_17_26_i = temp_b5_17_26_i;
assign out_17_27_r = temp_b5_17_27_r;
assign out_17_27_i = temp_b5_17_27_i;
assign out_17_28_r = temp_b5_17_28_r;
assign out_17_28_i = temp_b5_17_28_i;
assign out_17_29_r = temp_b5_17_29_r;
assign out_17_29_i = temp_b5_17_29_i;
assign out_17_30_r = temp_b5_17_30_r;
assign out_17_30_i = temp_b5_17_30_i;
assign out_17_31_r = temp_b5_17_31_r;
assign out_17_31_i = temp_b5_17_31_i;
assign out_17_32_r = temp_b5_17_32_r;
assign out_17_32_i = temp_b5_17_32_i;
assign out_18_1_r = temp_b5_18_1_r;
assign out_18_1_i = temp_b5_18_1_i;
assign out_18_2_r = temp_b5_18_2_r;
assign out_18_2_i = temp_b5_18_2_i;
assign out_18_3_r = temp_b5_18_3_r;
assign out_18_3_i = temp_b5_18_3_i;
assign out_18_4_r = temp_b5_18_4_r;
assign out_18_4_i = temp_b5_18_4_i;
assign out_18_5_r = temp_b5_18_5_r;
assign out_18_5_i = temp_b5_18_5_i;
assign out_18_6_r = temp_b5_18_6_r;
assign out_18_6_i = temp_b5_18_6_i;
assign out_18_7_r = temp_b5_18_7_r;
assign out_18_7_i = temp_b5_18_7_i;
assign out_18_8_r = temp_b5_18_8_r;
assign out_18_8_i = temp_b5_18_8_i;
assign out_18_9_r = temp_b5_18_9_r;
assign out_18_9_i = temp_b5_18_9_i;
assign out_18_10_r = temp_b5_18_10_r;
assign out_18_10_i = temp_b5_18_10_i;
assign out_18_11_r = temp_b5_18_11_r;
assign out_18_11_i = temp_b5_18_11_i;
assign out_18_12_r = temp_b5_18_12_r;
assign out_18_12_i = temp_b5_18_12_i;
assign out_18_13_r = temp_b5_18_13_r;
assign out_18_13_i = temp_b5_18_13_i;
assign out_18_14_r = temp_b5_18_14_r;
assign out_18_14_i = temp_b5_18_14_i;
assign out_18_15_r = temp_b5_18_15_r;
assign out_18_15_i = temp_b5_18_15_i;
assign out_18_16_r = temp_b5_18_16_r;
assign out_18_16_i = temp_b5_18_16_i;
assign out_18_17_r = temp_b5_18_17_r;
assign out_18_17_i = temp_b5_18_17_i;
assign out_18_18_r = temp_b5_18_18_r;
assign out_18_18_i = temp_b5_18_18_i;
assign out_18_19_r = temp_b5_18_19_r;
assign out_18_19_i = temp_b5_18_19_i;
assign out_18_20_r = temp_b5_18_20_r;
assign out_18_20_i = temp_b5_18_20_i;
assign out_18_21_r = temp_b5_18_21_r;
assign out_18_21_i = temp_b5_18_21_i;
assign out_18_22_r = temp_b5_18_22_r;
assign out_18_22_i = temp_b5_18_22_i;
assign out_18_23_r = temp_b5_18_23_r;
assign out_18_23_i = temp_b5_18_23_i;
assign out_18_24_r = temp_b5_18_24_r;
assign out_18_24_i = temp_b5_18_24_i;
assign out_18_25_r = temp_b5_18_25_r;
assign out_18_25_i = temp_b5_18_25_i;
assign out_18_26_r = temp_b5_18_26_r;
assign out_18_26_i = temp_b5_18_26_i;
assign out_18_27_r = temp_b5_18_27_r;
assign out_18_27_i = temp_b5_18_27_i;
assign out_18_28_r = temp_b5_18_28_r;
assign out_18_28_i = temp_b5_18_28_i;
assign out_18_29_r = temp_b5_18_29_r;
assign out_18_29_i = temp_b5_18_29_i;
assign out_18_30_r = temp_b5_18_30_r;
assign out_18_30_i = temp_b5_18_30_i;
assign out_18_31_r = temp_b5_18_31_r;
assign out_18_31_i = temp_b5_18_31_i;
assign out_18_32_r = temp_b5_18_32_r;
assign out_18_32_i = temp_b5_18_32_i;
assign out_19_1_r = temp_b5_19_1_r;
assign out_19_1_i = temp_b5_19_1_i;
assign out_19_2_r = temp_b5_19_2_r;
assign out_19_2_i = temp_b5_19_2_i;
assign out_19_3_r = temp_b5_19_3_r;
assign out_19_3_i = temp_b5_19_3_i;
assign out_19_4_r = temp_b5_19_4_r;
assign out_19_4_i = temp_b5_19_4_i;
assign out_19_5_r = temp_b5_19_5_r;
assign out_19_5_i = temp_b5_19_5_i;
assign out_19_6_r = temp_b5_19_6_r;
assign out_19_6_i = temp_b5_19_6_i;
assign out_19_7_r = temp_b5_19_7_r;
assign out_19_7_i = temp_b5_19_7_i;
assign out_19_8_r = temp_b5_19_8_r;
assign out_19_8_i = temp_b5_19_8_i;
assign out_19_9_r = temp_b5_19_9_r;
assign out_19_9_i = temp_b5_19_9_i;
assign out_19_10_r = temp_b5_19_10_r;
assign out_19_10_i = temp_b5_19_10_i;
assign out_19_11_r = temp_b5_19_11_r;
assign out_19_11_i = temp_b5_19_11_i;
assign out_19_12_r = temp_b5_19_12_r;
assign out_19_12_i = temp_b5_19_12_i;
assign out_19_13_r = temp_b5_19_13_r;
assign out_19_13_i = temp_b5_19_13_i;
assign out_19_14_r = temp_b5_19_14_r;
assign out_19_14_i = temp_b5_19_14_i;
assign out_19_15_r = temp_b5_19_15_r;
assign out_19_15_i = temp_b5_19_15_i;
assign out_19_16_r = temp_b5_19_16_r;
assign out_19_16_i = temp_b5_19_16_i;
assign out_19_17_r = temp_b5_19_17_r;
assign out_19_17_i = temp_b5_19_17_i;
assign out_19_18_r = temp_b5_19_18_r;
assign out_19_18_i = temp_b5_19_18_i;
assign out_19_19_r = temp_b5_19_19_r;
assign out_19_19_i = temp_b5_19_19_i;
assign out_19_20_r = temp_b5_19_20_r;
assign out_19_20_i = temp_b5_19_20_i;
assign out_19_21_r = temp_b5_19_21_r;
assign out_19_21_i = temp_b5_19_21_i;
assign out_19_22_r = temp_b5_19_22_r;
assign out_19_22_i = temp_b5_19_22_i;
assign out_19_23_r = temp_b5_19_23_r;
assign out_19_23_i = temp_b5_19_23_i;
assign out_19_24_r = temp_b5_19_24_r;
assign out_19_24_i = temp_b5_19_24_i;
assign out_19_25_r = temp_b5_19_25_r;
assign out_19_25_i = temp_b5_19_25_i;
assign out_19_26_r = temp_b5_19_26_r;
assign out_19_26_i = temp_b5_19_26_i;
assign out_19_27_r = temp_b5_19_27_r;
assign out_19_27_i = temp_b5_19_27_i;
assign out_19_28_r = temp_b5_19_28_r;
assign out_19_28_i = temp_b5_19_28_i;
assign out_19_29_r = temp_b5_19_29_r;
assign out_19_29_i = temp_b5_19_29_i;
assign out_19_30_r = temp_b5_19_30_r;
assign out_19_30_i = temp_b5_19_30_i;
assign out_19_31_r = temp_b5_19_31_r;
assign out_19_31_i = temp_b5_19_31_i;
assign out_19_32_r = temp_b5_19_32_r;
assign out_19_32_i = temp_b5_19_32_i;
assign out_20_1_r = temp_b5_20_1_r;
assign out_20_1_i = temp_b5_20_1_i;
assign out_20_2_r = temp_b5_20_2_r;
assign out_20_2_i = temp_b5_20_2_i;
assign out_20_3_r = temp_b5_20_3_r;
assign out_20_3_i = temp_b5_20_3_i;
assign out_20_4_r = temp_b5_20_4_r;
assign out_20_4_i = temp_b5_20_4_i;
assign out_20_5_r = temp_b5_20_5_r;
assign out_20_5_i = temp_b5_20_5_i;
assign out_20_6_r = temp_b5_20_6_r;
assign out_20_6_i = temp_b5_20_6_i;
assign out_20_7_r = temp_b5_20_7_r;
assign out_20_7_i = temp_b5_20_7_i;
assign out_20_8_r = temp_b5_20_8_r;
assign out_20_8_i = temp_b5_20_8_i;
assign out_20_9_r = temp_b5_20_9_r;
assign out_20_9_i = temp_b5_20_9_i;
assign out_20_10_r = temp_b5_20_10_r;
assign out_20_10_i = temp_b5_20_10_i;
assign out_20_11_r = temp_b5_20_11_r;
assign out_20_11_i = temp_b5_20_11_i;
assign out_20_12_r = temp_b5_20_12_r;
assign out_20_12_i = temp_b5_20_12_i;
assign out_20_13_r = temp_b5_20_13_r;
assign out_20_13_i = temp_b5_20_13_i;
assign out_20_14_r = temp_b5_20_14_r;
assign out_20_14_i = temp_b5_20_14_i;
assign out_20_15_r = temp_b5_20_15_r;
assign out_20_15_i = temp_b5_20_15_i;
assign out_20_16_r = temp_b5_20_16_r;
assign out_20_16_i = temp_b5_20_16_i;
assign out_20_17_r = temp_b5_20_17_r;
assign out_20_17_i = temp_b5_20_17_i;
assign out_20_18_r = temp_b5_20_18_r;
assign out_20_18_i = temp_b5_20_18_i;
assign out_20_19_r = temp_b5_20_19_r;
assign out_20_19_i = temp_b5_20_19_i;
assign out_20_20_r = temp_b5_20_20_r;
assign out_20_20_i = temp_b5_20_20_i;
assign out_20_21_r = temp_b5_20_21_r;
assign out_20_21_i = temp_b5_20_21_i;
assign out_20_22_r = temp_b5_20_22_r;
assign out_20_22_i = temp_b5_20_22_i;
assign out_20_23_r = temp_b5_20_23_r;
assign out_20_23_i = temp_b5_20_23_i;
assign out_20_24_r = temp_b5_20_24_r;
assign out_20_24_i = temp_b5_20_24_i;
assign out_20_25_r = temp_b5_20_25_r;
assign out_20_25_i = temp_b5_20_25_i;
assign out_20_26_r = temp_b5_20_26_r;
assign out_20_26_i = temp_b5_20_26_i;
assign out_20_27_r = temp_b5_20_27_r;
assign out_20_27_i = temp_b5_20_27_i;
assign out_20_28_r = temp_b5_20_28_r;
assign out_20_28_i = temp_b5_20_28_i;
assign out_20_29_r = temp_b5_20_29_r;
assign out_20_29_i = temp_b5_20_29_i;
assign out_20_30_r = temp_b5_20_30_r;
assign out_20_30_i = temp_b5_20_30_i;
assign out_20_31_r = temp_b5_20_31_r;
assign out_20_31_i = temp_b5_20_31_i;
assign out_20_32_r = temp_b5_20_32_r;
assign out_20_32_i = temp_b5_20_32_i;
assign out_21_1_r = temp_b5_21_1_r;
assign out_21_1_i = temp_b5_21_1_i;
assign out_21_2_r = temp_b5_21_2_r;
assign out_21_2_i = temp_b5_21_2_i;
assign out_21_3_r = temp_b5_21_3_r;
assign out_21_3_i = temp_b5_21_3_i;
assign out_21_4_r = temp_b5_21_4_r;
assign out_21_4_i = temp_b5_21_4_i;
assign out_21_5_r = temp_b5_21_5_r;
assign out_21_5_i = temp_b5_21_5_i;
assign out_21_6_r = temp_b5_21_6_r;
assign out_21_6_i = temp_b5_21_6_i;
assign out_21_7_r = temp_b5_21_7_r;
assign out_21_7_i = temp_b5_21_7_i;
assign out_21_8_r = temp_b5_21_8_r;
assign out_21_8_i = temp_b5_21_8_i;
assign out_21_9_r = temp_b5_21_9_r;
assign out_21_9_i = temp_b5_21_9_i;
assign out_21_10_r = temp_b5_21_10_r;
assign out_21_10_i = temp_b5_21_10_i;
assign out_21_11_r = temp_b5_21_11_r;
assign out_21_11_i = temp_b5_21_11_i;
assign out_21_12_r = temp_b5_21_12_r;
assign out_21_12_i = temp_b5_21_12_i;
assign out_21_13_r = temp_b5_21_13_r;
assign out_21_13_i = temp_b5_21_13_i;
assign out_21_14_r = temp_b5_21_14_r;
assign out_21_14_i = temp_b5_21_14_i;
assign out_21_15_r = temp_b5_21_15_r;
assign out_21_15_i = temp_b5_21_15_i;
assign out_21_16_r = temp_b5_21_16_r;
assign out_21_16_i = temp_b5_21_16_i;
assign out_21_17_r = temp_b5_21_17_r;
assign out_21_17_i = temp_b5_21_17_i;
assign out_21_18_r = temp_b5_21_18_r;
assign out_21_18_i = temp_b5_21_18_i;
assign out_21_19_r = temp_b5_21_19_r;
assign out_21_19_i = temp_b5_21_19_i;
assign out_21_20_r = temp_b5_21_20_r;
assign out_21_20_i = temp_b5_21_20_i;
assign out_21_21_r = temp_b5_21_21_r;
assign out_21_21_i = temp_b5_21_21_i;
assign out_21_22_r = temp_b5_21_22_r;
assign out_21_22_i = temp_b5_21_22_i;
assign out_21_23_r = temp_b5_21_23_r;
assign out_21_23_i = temp_b5_21_23_i;
assign out_21_24_r = temp_b5_21_24_r;
assign out_21_24_i = temp_b5_21_24_i;
assign out_21_25_r = temp_b5_21_25_r;
assign out_21_25_i = temp_b5_21_25_i;
assign out_21_26_r = temp_b5_21_26_r;
assign out_21_26_i = temp_b5_21_26_i;
assign out_21_27_r = temp_b5_21_27_r;
assign out_21_27_i = temp_b5_21_27_i;
assign out_21_28_r = temp_b5_21_28_r;
assign out_21_28_i = temp_b5_21_28_i;
assign out_21_29_r = temp_b5_21_29_r;
assign out_21_29_i = temp_b5_21_29_i;
assign out_21_30_r = temp_b5_21_30_r;
assign out_21_30_i = temp_b5_21_30_i;
assign out_21_31_r = temp_b5_21_31_r;
assign out_21_31_i = temp_b5_21_31_i;
assign out_21_32_r = temp_b5_21_32_r;
assign out_21_32_i = temp_b5_21_32_i;
assign out_22_1_r = temp_b5_22_1_r;
assign out_22_1_i = temp_b5_22_1_i;
assign out_22_2_r = temp_b5_22_2_r;
assign out_22_2_i = temp_b5_22_2_i;
assign out_22_3_r = temp_b5_22_3_r;
assign out_22_3_i = temp_b5_22_3_i;
assign out_22_4_r = temp_b5_22_4_r;
assign out_22_4_i = temp_b5_22_4_i;
assign out_22_5_r = temp_b5_22_5_r;
assign out_22_5_i = temp_b5_22_5_i;
assign out_22_6_r = temp_b5_22_6_r;
assign out_22_6_i = temp_b5_22_6_i;
assign out_22_7_r = temp_b5_22_7_r;
assign out_22_7_i = temp_b5_22_7_i;
assign out_22_8_r = temp_b5_22_8_r;
assign out_22_8_i = temp_b5_22_8_i;
assign out_22_9_r = temp_b5_22_9_r;
assign out_22_9_i = temp_b5_22_9_i;
assign out_22_10_r = temp_b5_22_10_r;
assign out_22_10_i = temp_b5_22_10_i;
assign out_22_11_r = temp_b5_22_11_r;
assign out_22_11_i = temp_b5_22_11_i;
assign out_22_12_r = temp_b5_22_12_r;
assign out_22_12_i = temp_b5_22_12_i;
assign out_22_13_r = temp_b5_22_13_r;
assign out_22_13_i = temp_b5_22_13_i;
assign out_22_14_r = temp_b5_22_14_r;
assign out_22_14_i = temp_b5_22_14_i;
assign out_22_15_r = temp_b5_22_15_r;
assign out_22_15_i = temp_b5_22_15_i;
assign out_22_16_r = temp_b5_22_16_r;
assign out_22_16_i = temp_b5_22_16_i;
assign out_22_17_r = temp_b5_22_17_r;
assign out_22_17_i = temp_b5_22_17_i;
assign out_22_18_r = temp_b5_22_18_r;
assign out_22_18_i = temp_b5_22_18_i;
assign out_22_19_r = temp_b5_22_19_r;
assign out_22_19_i = temp_b5_22_19_i;
assign out_22_20_r = temp_b5_22_20_r;
assign out_22_20_i = temp_b5_22_20_i;
assign out_22_21_r = temp_b5_22_21_r;
assign out_22_21_i = temp_b5_22_21_i;
assign out_22_22_r = temp_b5_22_22_r;
assign out_22_22_i = temp_b5_22_22_i;
assign out_22_23_r = temp_b5_22_23_r;
assign out_22_23_i = temp_b5_22_23_i;
assign out_22_24_r = temp_b5_22_24_r;
assign out_22_24_i = temp_b5_22_24_i;
assign out_22_25_r = temp_b5_22_25_r;
assign out_22_25_i = temp_b5_22_25_i;
assign out_22_26_r = temp_b5_22_26_r;
assign out_22_26_i = temp_b5_22_26_i;
assign out_22_27_r = temp_b5_22_27_r;
assign out_22_27_i = temp_b5_22_27_i;
assign out_22_28_r = temp_b5_22_28_r;
assign out_22_28_i = temp_b5_22_28_i;
assign out_22_29_r = temp_b5_22_29_r;
assign out_22_29_i = temp_b5_22_29_i;
assign out_22_30_r = temp_b5_22_30_r;
assign out_22_30_i = temp_b5_22_30_i;
assign out_22_31_r = temp_b5_22_31_r;
assign out_22_31_i = temp_b5_22_31_i;
assign out_22_32_r = temp_b5_22_32_r;
assign out_22_32_i = temp_b5_22_32_i;
assign out_23_1_r = temp_b5_23_1_r;
assign out_23_1_i = temp_b5_23_1_i;
assign out_23_2_r = temp_b5_23_2_r;
assign out_23_2_i = temp_b5_23_2_i;
assign out_23_3_r = temp_b5_23_3_r;
assign out_23_3_i = temp_b5_23_3_i;
assign out_23_4_r = temp_b5_23_4_r;
assign out_23_4_i = temp_b5_23_4_i;
assign out_23_5_r = temp_b5_23_5_r;
assign out_23_5_i = temp_b5_23_5_i;
assign out_23_6_r = temp_b5_23_6_r;
assign out_23_6_i = temp_b5_23_6_i;
assign out_23_7_r = temp_b5_23_7_r;
assign out_23_7_i = temp_b5_23_7_i;
assign out_23_8_r = temp_b5_23_8_r;
assign out_23_8_i = temp_b5_23_8_i;
assign out_23_9_r = temp_b5_23_9_r;
assign out_23_9_i = temp_b5_23_9_i;
assign out_23_10_r = temp_b5_23_10_r;
assign out_23_10_i = temp_b5_23_10_i;
assign out_23_11_r = temp_b5_23_11_r;
assign out_23_11_i = temp_b5_23_11_i;
assign out_23_12_r = temp_b5_23_12_r;
assign out_23_12_i = temp_b5_23_12_i;
assign out_23_13_r = temp_b5_23_13_r;
assign out_23_13_i = temp_b5_23_13_i;
assign out_23_14_r = temp_b5_23_14_r;
assign out_23_14_i = temp_b5_23_14_i;
assign out_23_15_r = temp_b5_23_15_r;
assign out_23_15_i = temp_b5_23_15_i;
assign out_23_16_r = temp_b5_23_16_r;
assign out_23_16_i = temp_b5_23_16_i;
assign out_23_17_r = temp_b5_23_17_r;
assign out_23_17_i = temp_b5_23_17_i;
assign out_23_18_r = temp_b5_23_18_r;
assign out_23_18_i = temp_b5_23_18_i;
assign out_23_19_r = temp_b5_23_19_r;
assign out_23_19_i = temp_b5_23_19_i;
assign out_23_20_r = temp_b5_23_20_r;
assign out_23_20_i = temp_b5_23_20_i;
assign out_23_21_r = temp_b5_23_21_r;
assign out_23_21_i = temp_b5_23_21_i;
assign out_23_22_r = temp_b5_23_22_r;
assign out_23_22_i = temp_b5_23_22_i;
assign out_23_23_r = temp_b5_23_23_r;
assign out_23_23_i = temp_b5_23_23_i;
assign out_23_24_r = temp_b5_23_24_r;
assign out_23_24_i = temp_b5_23_24_i;
assign out_23_25_r = temp_b5_23_25_r;
assign out_23_25_i = temp_b5_23_25_i;
assign out_23_26_r = temp_b5_23_26_r;
assign out_23_26_i = temp_b5_23_26_i;
assign out_23_27_r = temp_b5_23_27_r;
assign out_23_27_i = temp_b5_23_27_i;
assign out_23_28_r = temp_b5_23_28_r;
assign out_23_28_i = temp_b5_23_28_i;
assign out_23_29_r = temp_b5_23_29_r;
assign out_23_29_i = temp_b5_23_29_i;
assign out_23_30_r = temp_b5_23_30_r;
assign out_23_30_i = temp_b5_23_30_i;
assign out_23_31_r = temp_b5_23_31_r;
assign out_23_31_i = temp_b5_23_31_i;
assign out_23_32_r = temp_b5_23_32_r;
assign out_23_32_i = temp_b5_23_32_i;
assign out_24_1_r = temp_b5_24_1_r;
assign out_24_1_i = temp_b5_24_1_i;
assign out_24_2_r = temp_b5_24_2_r;
assign out_24_2_i = temp_b5_24_2_i;
assign out_24_3_r = temp_b5_24_3_r;
assign out_24_3_i = temp_b5_24_3_i;
assign out_24_4_r = temp_b5_24_4_r;
assign out_24_4_i = temp_b5_24_4_i;
assign out_24_5_r = temp_b5_24_5_r;
assign out_24_5_i = temp_b5_24_5_i;
assign out_24_6_r = temp_b5_24_6_r;
assign out_24_6_i = temp_b5_24_6_i;
assign out_24_7_r = temp_b5_24_7_r;
assign out_24_7_i = temp_b5_24_7_i;
assign out_24_8_r = temp_b5_24_8_r;
assign out_24_8_i = temp_b5_24_8_i;
assign out_24_9_r = temp_b5_24_9_r;
assign out_24_9_i = temp_b5_24_9_i;
assign out_24_10_r = temp_b5_24_10_r;
assign out_24_10_i = temp_b5_24_10_i;
assign out_24_11_r = temp_b5_24_11_r;
assign out_24_11_i = temp_b5_24_11_i;
assign out_24_12_r = temp_b5_24_12_r;
assign out_24_12_i = temp_b5_24_12_i;
assign out_24_13_r = temp_b5_24_13_r;
assign out_24_13_i = temp_b5_24_13_i;
assign out_24_14_r = temp_b5_24_14_r;
assign out_24_14_i = temp_b5_24_14_i;
assign out_24_15_r = temp_b5_24_15_r;
assign out_24_15_i = temp_b5_24_15_i;
assign out_24_16_r = temp_b5_24_16_r;
assign out_24_16_i = temp_b5_24_16_i;
assign out_24_17_r = temp_b5_24_17_r;
assign out_24_17_i = temp_b5_24_17_i;
assign out_24_18_r = temp_b5_24_18_r;
assign out_24_18_i = temp_b5_24_18_i;
assign out_24_19_r = temp_b5_24_19_r;
assign out_24_19_i = temp_b5_24_19_i;
assign out_24_20_r = temp_b5_24_20_r;
assign out_24_20_i = temp_b5_24_20_i;
assign out_24_21_r = temp_b5_24_21_r;
assign out_24_21_i = temp_b5_24_21_i;
assign out_24_22_r = temp_b5_24_22_r;
assign out_24_22_i = temp_b5_24_22_i;
assign out_24_23_r = temp_b5_24_23_r;
assign out_24_23_i = temp_b5_24_23_i;
assign out_24_24_r = temp_b5_24_24_r;
assign out_24_24_i = temp_b5_24_24_i;
assign out_24_25_r = temp_b5_24_25_r;
assign out_24_25_i = temp_b5_24_25_i;
assign out_24_26_r = temp_b5_24_26_r;
assign out_24_26_i = temp_b5_24_26_i;
assign out_24_27_r = temp_b5_24_27_r;
assign out_24_27_i = temp_b5_24_27_i;
assign out_24_28_r = temp_b5_24_28_r;
assign out_24_28_i = temp_b5_24_28_i;
assign out_24_29_r = temp_b5_24_29_r;
assign out_24_29_i = temp_b5_24_29_i;
assign out_24_30_r = temp_b5_24_30_r;
assign out_24_30_i = temp_b5_24_30_i;
assign out_24_31_r = temp_b5_24_31_r;
assign out_24_31_i = temp_b5_24_31_i;
assign out_24_32_r = temp_b5_24_32_r;
assign out_24_32_i = temp_b5_24_32_i;
assign out_25_1_r = temp_b5_25_1_r;
assign out_25_1_i = temp_b5_25_1_i;
assign out_25_2_r = temp_b5_25_2_r;
assign out_25_2_i = temp_b5_25_2_i;
assign out_25_3_r = temp_b5_25_3_r;
assign out_25_3_i = temp_b5_25_3_i;
assign out_25_4_r = temp_b5_25_4_r;
assign out_25_4_i = temp_b5_25_4_i;
assign out_25_5_r = temp_b5_25_5_r;
assign out_25_5_i = temp_b5_25_5_i;
assign out_25_6_r = temp_b5_25_6_r;
assign out_25_6_i = temp_b5_25_6_i;
assign out_25_7_r = temp_b5_25_7_r;
assign out_25_7_i = temp_b5_25_7_i;
assign out_25_8_r = temp_b5_25_8_r;
assign out_25_8_i = temp_b5_25_8_i;
assign out_25_9_r = temp_b5_25_9_r;
assign out_25_9_i = temp_b5_25_9_i;
assign out_25_10_r = temp_b5_25_10_r;
assign out_25_10_i = temp_b5_25_10_i;
assign out_25_11_r = temp_b5_25_11_r;
assign out_25_11_i = temp_b5_25_11_i;
assign out_25_12_r = temp_b5_25_12_r;
assign out_25_12_i = temp_b5_25_12_i;
assign out_25_13_r = temp_b5_25_13_r;
assign out_25_13_i = temp_b5_25_13_i;
assign out_25_14_r = temp_b5_25_14_r;
assign out_25_14_i = temp_b5_25_14_i;
assign out_25_15_r = temp_b5_25_15_r;
assign out_25_15_i = temp_b5_25_15_i;
assign out_25_16_r = temp_b5_25_16_r;
assign out_25_16_i = temp_b5_25_16_i;
assign out_25_17_r = temp_b5_25_17_r;
assign out_25_17_i = temp_b5_25_17_i;
assign out_25_18_r = temp_b5_25_18_r;
assign out_25_18_i = temp_b5_25_18_i;
assign out_25_19_r = temp_b5_25_19_r;
assign out_25_19_i = temp_b5_25_19_i;
assign out_25_20_r = temp_b5_25_20_r;
assign out_25_20_i = temp_b5_25_20_i;
assign out_25_21_r = temp_b5_25_21_r;
assign out_25_21_i = temp_b5_25_21_i;
assign out_25_22_r = temp_b5_25_22_r;
assign out_25_22_i = temp_b5_25_22_i;
assign out_25_23_r = temp_b5_25_23_r;
assign out_25_23_i = temp_b5_25_23_i;
assign out_25_24_r = temp_b5_25_24_r;
assign out_25_24_i = temp_b5_25_24_i;
assign out_25_25_r = temp_b5_25_25_r;
assign out_25_25_i = temp_b5_25_25_i;
assign out_25_26_r = temp_b5_25_26_r;
assign out_25_26_i = temp_b5_25_26_i;
assign out_25_27_r = temp_b5_25_27_r;
assign out_25_27_i = temp_b5_25_27_i;
assign out_25_28_r = temp_b5_25_28_r;
assign out_25_28_i = temp_b5_25_28_i;
assign out_25_29_r = temp_b5_25_29_r;
assign out_25_29_i = temp_b5_25_29_i;
assign out_25_30_r = temp_b5_25_30_r;
assign out_25_30_i = temp_b5_25_30_i;
assign out_25_31_r = temp_b5_25_31_r;
assign out_25_31_i = temp_b5_25_31_i;
assign out_25_32_r = temp_b5_25_32_r;
assign out_25_32_i = temp_b5_25_32_i;
assign out_26_1_r = temp_b5_26_1_r;
assign out_26_1_i = temp_b5_26_1_i;
assign out_26_2_r = temp_b5_26_2_r;
assign out_26_2_i = temp_b5_26_2_i;
assign out_26_3_r = temp_b5_26_3_r;
assign out_26_3_i = temp_b5_26_3_i;
assign out_26_4_r = temp_b5_26_4_r;
assign out_26_4_i = temp_b5_26_4_i;
assign out_26_5_r = temp_b5_26_5_r;
assign out_26_5_i = temp_b5_26_5_i;
assign out_26_6_r = temp_b5_26_6_r;
assign out_26_6_i = temp_b5_26_6_i;
assign out_26_7_r = temp_b5_26_7_r;
assign out_26_7_i = temp_b5_26_7_i;
assign out_26_8_r = temp_b5_26_8_r;
assign out_26_8_i = temp_b5_26_8_i;
assign out_26_9_r = temp_b5_26_9_r;
assign out_26_9_i = temp_b5_26_9_i;
assign out_26_10_r = temp_b5_26_10_r;
assign out_26_10_i = temp_b5_26_10_i;
assign out_26_11_r = temp_b5_26_11_r;
assign out_26_11_i = temp_b5_26_11_i;
assign out_26_12_r = temp_b5_26_12_r;
assign out_26_12_i = temp_b5_26_12_i;
assign out_26_13_r = temp_b5_26_13_r;
assign out_26_13_i = temp_b5_26_13_i;
assign out_26_14_r = temp_b5_26_14_r;
assign out_26_14_i = temp_b5_26_14_i;
assign out_26_15_r = temp_b5_26_15_r;
assign out_26_15_i = temp_b5_26_15_i;
assign out_26_16_r = temp_b5_26_16_r;
assign out_26_16_i = temp_b5_26_16_i;
assign out_26_17_r = temp_b5_26_17_r;
assign out_26_17_i = temp_b5_26_17_i;
assign out_26_18_r = temp_b5_26_18_r;
assign out_26_18_i = temp_b5_26_18_i;
assign out_26_19_r = temp_b5_26_19_r;
assign out_26_19_i = temp_b5_26_19_i;
assign out_26_20_r = temp_b5_26_20_r;
assign out_26_20_i = temp_b5_26_20_i;
assign out_26_21_r = temp_b5_26_21_r;
assign out_26_21_i = temp_b5_26_21_i;
assign out_26_22_r = temp_b5_26_22_r;
assign out_26_22_i = temp_b5_26_22_i;
assign out_26_23_r = temp_b5_26_23_r;
assign out_26_23_i = temp_b5_26_23_i;
assign out_26_24_r = temp_b5_26_24_r;
assign out_26_24_i = temp_b5_26_24_i;
assign out_26_25_r = temp_b5_26_25_r;
assign out_26_25_i = temp_b5_26_25_i;
assign out_26_26_r = temp_b5_26_26_r;
assign out_26_26_i = temp_b5_26_26_i;
assign out_26_27_r = temp_b5_26_27_r;
assign out_26_27_i = temp_b5_26_27_i;
assign out_26_28_r = temp_b5_26_28_r;
assign out_26_28_i = temp_b5_26_28_i;
assign out_26_29_r = temp_b5_26_29_r;
assign out_26_29_i = temp_b5_26_29_i;
assign out_26_30_r = temp_b5_26_30_r;
assign out_26_30_i = temp_b5_26_30_i;
assign out_26_31_r = temp_b5_26_31_r;
assign out_26_31_i = temp_b5_26_31_i;
assign out_26_32_r = temp_b5_26_32_r;
assign out_26_32_i = temp_b5_26_32_i;
assign out_27_1_r = temp_b5_27_1_r;
assign out_27_1_i = temp_b5_27_1_i;
assign out_27_2_r = temp_b5_27_2_r;
assign out_27_2_i = temp_b5_27_2_i;
assign out_27_3_r = temp_b5_27_3_r;
assign out_27_3_i = temp_b5_27_3_i;
assign out_27_4_r = temp_b5_27_4_r;
assign out_27_4_i = temp_b5_27_4_i;
assign out_27_5_r = temp_b5_27_5_r;
assign out_27_5_i = temp_b5_27_5_i;
assign out_27_6_r = temp_b5_27_6_r;
assign out_27_6_i = temp_b5_27_6_i;
assign out_27_7_r = temp_b5_27_7_r;
assign out_27_7_i = temp_b5_27_7_i;
assign out_27_8_r = temp_b5_27_8_r;
assign out_27_8_i = temp_b5_27_8_i;
assign out_27_9_r = temp_b5_27_9_r;
assign out_27_9_i = temp_b5_27_9_i;
assign out_27_10_r = temp_b5_27_10_r;
assign out_27_10_i = temp_b5_27_10_i;
assign out_27_11_r = temp_b5_27_11_r;
assign out_27_11_i = temp_b5_27_11_i;
assign out_27_12_r = temp_b5_27_12_r;
assign out_27_12_i = temp_b5_27_12_i;
assign out_27_13_r = temp_b5_27_13_r;
assign out_27_13_i = temp_b5_27_13_i;
assign out_27_14_r = temp_b5_27_14_r;
assign out_27_14_i = temp_b5_27_14_i;
assign out_27_15_r = temp_b5_27_15_r;
assign out_27_15_i = temp_b5_27_15_i;
assign out_27_16_r = temp_b5_27_16_r;
assign out_27_16_i = temp_b5_27_16_i;
assign out_27_17_r = temp_b5_27_17_r;
assign out_27_17_i = temp_b5_27_17_i;
assign out_27_18_r = temp_b5_27_18_r;
assign out_27_18_i = temp_b5_27_18_i;
assign out_27_19_r = temp_b5_27_19_r;
assign out_27_19_i = temp_b5_27_19_i;
assign out_27_20_r = temp_b5_27_20_r;
assign out_27_20_i = temp_b5_27_20_i;
assign out_27_21_r = temp_b5_27_21_r;
assign out_27_21_i = temp_b5_27_21_i;
assign out_27_22_r = temp_b5_27_22_r;
assign out_27_22_i = temp_b5_27_22_i;
assign out_27_23_r = temp_b5_27_23_r;
assign out_27_23_i = temp_b5_27_23_i;
assign out_27_24_r = temp_b5_27_24_r;
assign out_27_24_i = temp_b5_27_24_i;
assign out_27_25_r = temp_b5_27_25_r;
assign out_27_25_i = temp_b5_27_25_i;
assign out_27_26_r = temp_b5_27_26_r;
assign out_27_26_i = temp_b5_27_26_i;
assign out_27_27_r = temp_b5_27_27_r;
assign out_27_27_i = temp_b5_27_27_i;
assign out_27_28_r = temp_b5_27_28_r;
assign out_27_28_i = temp_b5_27_28_i;
assign out_27_29_r = temp_b5_27_29_r;
assign out_27_29_i = temp_b5_27_29_i;
assign out_27_30_r = temp_b5_27_30_r;
assign out_27_30_i = temp_b5_27_30_i;
assign out_27_31_r = temp_b5_27_31_r;
assign out_27_31_i = temp_b5_27_31_i;
assign out_27_32_r = temp_b5_27_32_r;
assign out_27_32_i = temp_b5_27_32_i;
assign out_28_1_r = temp_b5_28_1_r;
assign out_28_1_i = temp_b5_28_1_i;
assign out_28_2_r = temp_b5_28_2_r;
assign out_28_2_i = temp_b5_28_2_i;
assign out_28_3_r = temp_b5_28_3_r;
assign out_28_3_i = temp_b5_28_3_i;
assign out_28_4_r = temp_b5_28_4_r;
assign out_28_4_i = temp_b5_28_4_i;
assign out_28_5_r = temp_b5_28_5_r;
assign out_28_5_i = temp_b5_28_5_i;
assign out_28_6_r = temp_b5_28_6_r;
assign out_28_6_i = temp_b5_28_6_i;
assign out_28_7_r = temp_b5_28_7_r;
assign out_28_7_i = temp_b5_28_7_i;
assign out_28_8_r = temp_b5_28_8_r;
assign out_28_8_i = temp_b5_28_8_i;
assign out_28_9_r = temp_b5_28_9_r;
assign out_28_9_i = temp_b5_28_9_i;
assign out_28_10_r = temp_b5_28_10_r;
assign out_28_10_i = temp_b5_28_10_i;
assign out_28_11_r = temp_b5_28_11_r;
assign out_28_11_i = temp_b5_28_11_i;
assign out_28_12_r = temp_b5_28_12_r;
assign out_28_12_i = temp_b5_28_12_i;
assign out_28_13_r = temp_b5_28_13_r;
assign out_28_13_i = temp_b5_28_13_i;
assign out_28_14_r = temp_b5_28_14_r;
assign out_28_14_i = temp_b5_28_14_i;
assign out_28_15_r = temp_b5_28_15_r;
assign out_28_15_i = temp_b5_28_15_i;
assign out_28_16_r = temp_b5_28_16_r;
assign out_28_16_i = temp_b5_28_16_i;
assign out_28_17_r = temp_b5_28_17_r;
assign out_28_17_i = temp_b5_28_17_i;
assign out_28_18_r = temp_b5_28_18_r;
assign out_28_18_i = temp_b5_28_18_i;
assign out_28_19_r = temp_b5_28_19_r;
assign out_28_19_i = temp_b5_28_19_i;
assign out_28_20_r = temp_b5_28_20_r;
assign out_28_20_i = temp_b5_28_20_i;
assign out_28_21_r = temp_b5_28_21_r;
assign out_28_21_i = temp_b5_28_21_i;
assign out_28_22_r = temp_b5_28_22_r;
assign out_28_22_i = temp_b5_28_22_i;
assign out_28_23_r = temp_b5_28_23_r;
assign out_28_23_i = temp_b5_28_23_i;
assign out_28_24_r = temp_b5_28_24_r;
assign out_28_24_i = temp_b5_28_24_i;
assign out_28_25_r = temp_b5_28_25_r;
assign out_28_25_i = temp_b5_28_25_i;
assign out_28_26_r = temp_b5_28_26_r;
assign out_28_26_i = temp_b5_28_26_i;
assign out_28_27_r = temp_b5_28_27_r;
assign out_28_27_i = temp_b5_28_27_i;
assign out_28_28_r = temp_b5_28_28_r;
assign out_28_28_i = temp_b5_28_28_i;
assign out_28_29_r = temp_b5_28_29_r;
assign out_28_29_i = temp_b5_28_29_i;
assign out_28_30_r = temp_b5_28_30_r;
assign out_28_30_i = temp_b5_28_30_i;
assign out_28_31_r = temp_b5_28_31_r;
assign out_28_31_i = temp_b5_28_31_i;
assign out_28_32_r = temp_b5_28_32_r;
assign out_28_32_i = temp_b5_28_32_i;
assign out_29_1_r = temp_b5_29_1_r;
assign out_29_1_i = temp_b5_29_1_i;
assign out_29_2_r = temp_b5_29_2_r;
assign out_29_2_i = temp_b5_29_2_i;
assign out_29_3_r = temp_b5_29_3_r;
assign out_29_3_i = temp_b5_29_3_i;
assign out_29_4_r = temp_b5_29_4_r;
assign out_29_4_i = temp_b5_29_4_i;
assign out_29_5_r = temp_b5_29_5_r;
assign out_29_5_i = temp_b5_29_5_i;
assign out_29_6_r = temp_b5_29_6_r;
assign out_29_6_i = temp_b5_29_6_i;
assign out_29_7_r = temp_b5_29_7_r;
assign out_29_7_i = temp_b5_29_7_i;
assign out_29_8_r = temp_b5_29_8_r;
assign out_29_8_i = temp_b5_29_8_i;
assign out_29_9_r = temp_b5_29_9_r;
assign out_29_9_i = temp_b5_29_9_i;
assign out_29_10_r = temp_b5_29_10_r;
assign out_29_10_i = temp_b5_29_10_i;
assign out_29_11_r = temp_b5_29_11_r;
assign out_29_11_i = temp_b5_29_11_i;
assign out_29_12_r = temp_b5_29_12_r;
assign out_29_12_i = temp_b5_29_12_i;
assign out_29_13_r = temp_b5_29_13_r;
assign out_29_13_i = temp_b5_29_13_i;
assign out_29_14_r = temp_b5_29_14_r;
assign out_29_14_i = temp_b5_29_14_i;
assign out_29_15_r = temp_b5_29_15_r;
assign out_29_15_i = temp_b5_29_15_i;
assign out_29_16_r = temp_b5_29_16_r;
assign out_29_16_i = temp_b5_29_16_i;
assign out_29_17_r = temp_b5_29_17_r;
assign out_29_17_i = temp_b5_29_17_i;
assign out_29_18_r = temp_b5_29_18_r;
assign out_29_18_i = temp_b5_29_18_i;
assign out_29_19_r = temp_b5_29_19_r;
assign out_29_19_i = temp_b5_29_19_i;
assign out_29_20_r = temp_b5_29_20_r;
assign out_29_20_i = temp_b5_29_20_i;
assign out_29_21_r = temp_b5_29_21_r;
assign out_29_21_i = temp_b5_29_21_i;
assign out_29_22_r = temp_b5_29_22_r;
assign out_29_22_i = temp_b5_29_22_i;
assign out_29_23_r = temp_b5_29_23_r;
assign out_29_23_i = temp_b5_29_23_i;
assign out_29_24_r = temp_b5_29_24_r;
assign out_29_24_i = temp_b5_29_24_i;
assign out_29_25_r = temp_b5_29_25_r;
assign out_29_25_i = temp_b5_29_25_i;
assign out_29_26_r = temp_b5_29_26_r;
assign out_29_26_i = temp_b5_29_26_i;
assign out_29_27_r = temp_b5_29_27_r;
assign out_29_27_i = temp_b5_29_27_i;
assign out_29_28_r = temp_b5_29_28_r;
assign out_29_28_i = temp_b5_29_28_i;
assign out_29_29_r = temp_b5_29_29_r;
assign out_29_29_i = temp_b5_29_29_i;
assign out_29_30_r = temp_b5_29_30_r;
assign out_29_30_i = temp_b5_29_30_i;
assign out_29_31_r = temp_b5_29_31_r;
assign out_29_31_i = temp_b5_29_31_i;
assign out_29_32_r = temp_b5_29_32_r;
assign out_29_32_i = temp_b5_29_32_i;
assign out_30_1_r = temp_b5_30_1_r;
assign out_30_1_i = temp_b5_30_1_i;
assign out_30_2_r = temp_b5_30_2_r;
assign out_30_2_i = temp_b5_30_2_i;
assign out_30_3_r = temp_b5_30_3_r;
assign out_30_3_i = temp_b5_30_3_i;
assign out_30_4_r = temp_b5_30_4_r;
assign out_30_4_i = temp_b5_30_4_i;
assign out_30_5_r = temp_b5_30_5_r;
assign out_30_5_i = temp_b5_30_5_i;
assign out_30_6_r = temp_b5_30_6_r;
assign out_30_6_i = temp_b5_30_6_i;
assign out_30_7_r = temp_b5_30_7_r;
assign out_30_7_i = temp_b5_30_7_i;
assign out_30_8_r = temp_b5_30_8_r;
assign out_30_8_i = temp_b5_30_8_i;
assign out_30_9_r = temp_b5_30_9_r;
assign out_30_9_i = temp_b5_30_9_i;
assign out_30_10_r = temp_b5_30_10_r;
assign out_30_10_i = temp_b5_30_10_i;
assign out_30_11_r = temp_b5_30_11_r;
assign out_30_11_i = temp_b5_30_11_i;
assign out_30_12_r = temp_b5_30_12_r;
assign out_30_12_i = temp_b5_30_12_i;
assign out_30_13_r = temp_b5_30_13_r;
assign out_30_13_i = temp_b5_30_13_i;
assign out_30_14_r = temp_b5_30_14_r;
assign out_30_14_i = temp_b5_30_14_i;
assign out_30_15_r = temp_b5_30_15_r;
assign out_30_15_i = temp_b5_30_15_i;
assign out_30_16_r = temp_b5_30_16_r;
assign out_30_16_i = temp_b5_30_16_i;
assign out_30_17_r = temp_b5_30_17_r;
assign out_30_17_i = temp_b5_30_17_i;
assign out_30_18_r = temp_b5_30_18_r;
assign out_30_18_i = temp_b5_30_18_i;
assign out_30_19_r = temp_b5_30_19_r;
assign out_30_19_i = temp_b5_30_19_i;
assign out_30_20_r = temp_b5_30_20_r;
assign out_30_20_i = temp_b5_30_20_i;
assign out_30_21_r = temp_b5_30_21_r;
assign out_30_21_i = temp_b5_30_21_i;
assign out_30_22_r = temp_b5_30_22_r;
assign out_30_22_i = temp_b5_30_22_i;
assign out_30_23_r = temp_b5_30_23_r;
assign out_30_23_i = temp_b5_30_23_i;
assign out_30_24_r = temp_b5_30_24_r;
assign out_30_24_i = temp_b5_30_24_i;
assign out_30_25_r = temp_b5_30_25_r;
assign out_30_25_i = temp_b5_30_25_i;
assign out_30_26_r = temp_b5_30_26_r;
assign out_30_26_i = temp_b5_30_26_i;
assign out_30_27_r = temp_b5_30_27_r;
assign out_30_27_i = temp_b5_30_27_i;
assign out_30_28_r = temp_b5_30_28_r;
assign out_30_28_i = temp_b5_30_28_i;
assign out_30_29_r = temp_b5_30_29_r;
assign out_30_29_i = temp_b5_30_29_i;
assign out_30_30_r = temp_b5_30_30_r;
assign out_30_30_i = temp_b5_30_30_i;
assign out_30_31_r = temp_b5_30_31_r;
assign out_30_31_i = temp_b5_30_31_i;
assign out_30_32_r = temp_b5_30_32_r;
assign out_30_32_i = temp_b5_30_32_i;
assign out_31_1_r = temp_b5_31_1_r;
assign out_31_1_i = temp_b5_31_1_i;
assign out_31_2_r = temp_b5_31_2_r;
assign out_31_2_i = temp_b5_31_2_i;
assign out_31_3_r = temp_b5_31_3_r;
assign out_31_3_i = temp_b5_31_3_i;
assign out_31_4_r = temp_b5_31_4_r;
assign out_31_4_i = temp_b5_31_4_i;
assign out_31_5_r = temp_b5_31_5_r;
assign out_31_5_i = temp_b5_31_5_i;
assign out_31_6_r = temp_b5_31_6_r;
assign out_31_6_i = temp_b5_31_6_i;
assign out_31_7_r = temp_b5_31_7_r;
assign out_31_7_i = temp_b5_31_7_i;
assign out_31_8_r = temp_b5_31_8_r;
assign out_31_8_i = temp_b5_31_8_i;
assign out_31_9_r = temp_b5_31_9_r;
assign out_31_9_i = temp_b5_31_9_i;
assign out_31_10_r = temp_b5_31_10_r;
assign out_31_10_i = temp_b5_31_10_i;
assign out_31_11_r = temp_b5_31_11_r;
assign out_31_11_i = temp_b5_31_11_i;
assign out_31_12_r = temp_b5_31_12_r;
assign out_31_12_i = temp_b5_31_12_i;
assign out_31_13_r = temp_b5_31_13_r;
assign out_31_13_i = temp_b5_31_13_i;
assign out_31_14_r = temp_b5_31_14_r;
assign out_31_14_i = temp_b5_31_14_i;
assign out_31_15_r = temp_b5_31_15_r;
assign out_31_15_i = temp_b5_31_15_i;
assign out_31_16_r = temp_b5_31_16_r;
assign out_31_16_i = temp_b5_31_16_i;
assign out_31_17_r = temp_b5_31_17_r;
assign out_31_17_i = temp_b5_31_17_i;
assign out_31_18_r = temp_b5_31_18_r;
assign out_31_18_i = temp_b5_31_18_i;
assign out_31_19_r = temp_b5_31_19_r;
assign out_31_19_i = temp_b5_31_19_i;
assign out_31_20_r = temp_b5_31_20_r;
assign out_31_20_i = temp_b5_31_20_i;
assign out_31_21_r = temp_b5_31_21_r;
assign out_31_21_i = temp_b5_31_21_i;
assign out_31_22_r = temp_b5_31_22_r;
assign out_31_22_i = temp_b5_31_22_i;
assign out_31_23_r = temp_b5_31_23_r;
assign out_31_23_i = temp_b5_31_23_i;
assign out_31_24_r = temp_b5_31_24_r;
assign out_31_24_i = temp_b5_31_24_i;
assign out_31_25_r = temp_b5_31_25_r;
assign out_31_25_i = temp_b5_31_25_i;
assign out_31_26_r = temp_b5_31_26_r;
assign out_31_26_i = temp_b5_31_26_i;
assign out_31_27_r = temp_b5_31_27_r;
assign out_31_27_i = temp_b5_31_27_i;
assign out_31_28_r = temp_b5_31_28_r;
assign out_31_28_i = temp_b5_31_28_i;
assign out_31_29_r = temp_b5_31_29_r;
assign out_31_29_i = temp_b5_31_29_i;
assign out_31_30_r = temp_b5_31_30_r;
assign out_31_30_i = temp_b5_31_30_i;
assign out_31_31_r = temp_b5_31_31_r;
assign out_31_31_i = temp_b5_31_31_i;
assign out_31_32_r = temp_b5_31_32_r;
assign out_31_32_i = temp_b5_31_32_i;
assign out_32_1_r = temp_b5_32_1_r;
assign out_32_1_i = temp_b5_32_1_i;
assign out_32_2_r = temp_b5_32_2_r;
assign out_32_2_i = temp_b5_32_2_i;
assign out_32_3_r = temp_b5_32_3_r;
assign out_32_3_i = temp_b5_32_3_i;
assign out_32_4_r = temp_b5_32_4_r;
assign out_32_4_i = temp_b5_32_4_i;
assign out_32_5_r = temp_b5_32_5_r;
assign out_32_5_i = temp_b5_32_5_i;
assign out_32_6_r = temp_b5_32_6_r;
assign out_32_6_i = temp_b5_32_6_i;
assign out_32_7_r = temp_b5_32_7_r;
assign out_32_7_i = temp_b5_32_7_i;
assign out_32_8_r = temp_b5_32_8_r;
assign out_32_8_i = temp_b5_32_8_i;
assign out_32_9_r = temp_b5_32_9_r;
assign out_32_9_i = temp_b5_32_9_i;
assign out_32_10_r = temp_b5_32_10_r;
assign out_32_10_i = temp_b5_32_10_i;
assign out_32_11_r = temp_b5_32_11_r;
assign out_32_11_i = temp_b5_32_11_i;
assign out_32_12_r = temp_b5_32_12_r;
assign out_32_12_i = temp_b5_32_12_i;
assign out_32_13_r = temp_b5_32_13_r;
assign out_32_13_i = temp_b5_32_13_i;
assign out_32_14_r = temp_b5_32_14_r;
assign out_32_14_i = temp_b5_32_14_i;
assign out_32_15_r = temp_b5_32_15_r;
assign out_32_15_i = temp_b5_32_15_i;
assign out_32_16_r = temp_b5_32_16_r;
assign out_32_16_i = temp_b5_32_16_i;
assign out_32_17_r = temp_b5_32_17_r;
assign out_32_17_i = temp_b5_32_17_i;
assign out_32_18_r = temp_b5_32_18_r;
assign out_32_18_i = temp_b5_32_18_i;
assign out_32_19_r = temp_b5_32_19_r;
assign out_32_19_i = temp_b5_32_19_i;
assign out_32_20_r = temp_b5_32_20_r;
assign out_32_20_i = temp_b5_32_20_i;
assign out_32_21_r = temp_b5_32_21_r;
assign out_32_21_i = temp_b5_32_21_i;
assign out_32_22_r = temp_b5_32_22_r;
assign out_32_22_i = temp_b5_32_22_i;
assign out_32_23_r = temp_b5_32_23_r;
assign out_32_23_i = temp_b5_32_23_i;
assign out_32_24_r = temp_b5_32_24_r;
assign out_32_24_i = temp_b5_32_24_i;
assign out_32_25_r = temp_b5_32_25_r;
assign out_32_25_i = temp_b5_32_25_i;
assign out_32_26_r = temp_b5_32_26_r;
assign out_32_26_i = temp_b5_32_26_i;
assign out_32_27_r = temp_b5_32_27_r;
assign out_32_27_i = temp_b5_32_27_i;
assign out_32_28_r = temp_b5_32_28_r;
assign out_32_28_i = temp_b5_32_28_i;
assign out_32_29_r = temp_b5_32_29_r;
assign out_32_29_i = temp_b5_32_29_i;
assign out_32_30_r = temp_b5_32_30_r;
assign out_32_30_i = temp_b5_32_30_i;
assign out_32_31_r = temp_b5_32_31_r;
assign out_32_31_i = temp_b5_32_31_i;
assign out_32_32_r = temp_b5_32_32_r;
assign out_32_32_i = temp_b5_32_32_i;

assign out_r = out_1_1_r;
assign out_i = out_1_1_i;



endmodule
