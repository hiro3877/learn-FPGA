`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/08/25 18:20:35
// Design Name: 
// Module Name: top_sim
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module top_sim();

reg		clk;

reg signed [`InBus]		in_1_1_r;
reg signed [`InBus]		in_1_1_i;
reg signed [`InBus]		in_1_2_r;
reg signed [`InBus]		in_1_2_i;
reg signed [`InBus]		in_1_3_r;
reg signed [`InBus]		in_1_3_i;
reg signed [`InBus]		in_1_4_r;
reg signed [`InBus]		in_1_4_i;
reg signed [`InBus]		in_1_5_r;
reg signed [`InBus]		in_1_5_i;
reg signed [`InBus]		in_1_6_r;
reg signed [`InBus]		in_1_6_i;
reg signed [`InBus]		in_1_7_r;
reg signed [`InBus]		in_1_7_i;
reg signed [`InBus]		in_1_8_r;
reg signed [`InBus]		in_1_8_i;
reg signed [`InBus]		in_1_9_r;
reg signed [`InBus]		in_1_9_i;
reg signed [`InBus]		in_1_10_r;
reg signed [`InBus]		in_1_10_i;
reg signed [`InBus]		in_1_11_r;
reg signed [`InBus]		in_1_11_i;
reg signed [`InBus]		in_1_12_r;
reg signed [`InBus]		in_1_12_i;
reg signed [`InBus]		in_1_13_r;
reg signed [`InBus]		in_1_13_i;
reg signed [`InBus]		in_1_14_r;
reg signed [`InBus]		in_1_14_i;
reg signed [`InBus]		in_1_15_r;
reg signed [`InBus]		in_1_15_i;
reg signed [`InBus]		in_1_16_r;
reg signed [`InBus]		in_1_16_i;
reg signed [`InBus]		in_1_17_r;
reg signed [`InBus]		in_1_17_i;
reg signed [`InBus]		in_1_18_r;
reg signed [`InBus]		in_1_18_i;
reg signed [`InBus]		in_1_19_r;
reg signed [`InBus]		in_1_19_i;
reg signed [`InBus]		in_1_20_r;
reg signed [`InBus]		in_1_20_i;
reg signed [`InBus]		in_1_21_r;
reg signed [`InBus]		in_1_21_i;
reg signed [`InBus]		in_1_22_r;
reg signed [`InBus]		in_1_22_i;
reg signed [`InBus]		in_1_23_r;
reg signed [`InBus]		in_1_23_i;
reg signed [`InBus]		in_1_24_r;
reg signed [`InBus]		in_1_24_i;
reg signed [`InBus]		in_1_25_r;
reg signed [`InBus]		in_1_25_i;
reg signed [`InBus]		in_1_26_r;
reg signed [`InBus]		in_1_26_i;
reg signed [`InBus]		in_1_27_r;
reg signed [`InBus]		in_1_27_i;
reg signed [`InBus]		in_1_28_r;
reg signed [`InBus]		in_1_28_i;
reg signed [`InBus]		in_1_29_r;
reg signed [`InBus]		in_1_29_i;
reg signed [`InBus]		in_1_30_r;
reg signed [`InBus]		in_1_30_i;
reg signed [`InBus]		in_1_31_r;
reg signed [`InBus]		in_1_31_i;
reg signed [`InBus]		in_1_32_r;
reg signed [`InBus]		in_1_32_i;
reg signed [`InBus]		in_2_1_r;
reg signed [`InBus]		in_2_1_i;
reg signed [`InBus]		in_2_2_r;
reg signed [`InBus]		in_2_2_i;
reg signed [`InBus]		in_2_3_r;
reg signed [`InBus]		in_2_3_i;
reg signed [`InBus]		in_2_4_r;
reg signed [`InBus]		in_2_4_i;
reg signed [`InBus]		in_2_5_r;
reg signed [`InBus]		in_2_5_i;
reg signed [`InBus]		in_2_6_r;
reg signed [`InBus]		in_2_6_i;
reg signed [`InBus]		in_2_7_r;
reg signed [`InBus]		in_2_7_i;
reg signed [`InBus]		in_2_8_r;
reg signed [`InBus]		in_2_8_i;
reg signed [`InBus]		in_2_9_r;
reg signed [`InBus]		in_2_9_i;
reg signed [`InBus]		in_2_10_r;
reg signed [`InBus]		in_2_10_i;
reg signed [`InBus]		in_2_11_r;
reg signed [`InBus]		in_2_11_i;
reg signed [`InBus]		in_2_12_r;
reg signed [`InBus]		in_2_12_i;
reg signed [`InBus]		in_2_13_r;
reg signed [`InBus]		in_2_13_i;
reg signed [`InBus]		in_2_14_r;
reg signed [`InBus]		in_2_14_i;
reg signed [`InBus]		in_2_15_r;
reg signed [`InBus]		in_2_15_i;
reg signed [`InBus]		in_2_16_r;
reg signed [`InBus]		in_2_16_i;
reg signed [`InBus]		in_2_17_r;
reg signed [`InBus]		in_2_17_i;
reg signed [`InBus]		in_2_18_r;
reg signed [`InBus]		in_2_18_i;
reg signed [`InBus]		in_2_19_r;
reg signed [`InBus]		in_2_19_i;
reg signed [`InBus]		in_2_20_r;
reg signed [`InBus]		in_2_20_i;
reg signed [`InBus]		in_2_21_r;
reg signed [`InBus]		in_2_21_i;
reg signed [`InBus]		in_2_22_r;
reg signed [`InBus]		in_2_22_i;
reg signed [`InBus]		in_2_23_r;
reg signed [`InBus]		in_2_23_i;
reg signed [`InBus]		in_2_24_r;
reg signed [`InBus]		in_2_24_i;
reg signed [`InBus]		in_2_25_r;
reg signed [`InBus]		in_2_25_i;
reg signed [`InBus]		in_2_26_r;
reg signed [`InBus]		in_2_26_i;
reg signed [`InBus]		in_2_27_r;
reg signed [`InBus]		in_2_27_i;
reg signed [`InBus]		in_2_28_r;
reg signed [`InBus]		in_2_28_i;
reg signed [`InBus]		in_2_29_r;
reg signed [`InBus]		in_2_29_i;
reg signed [`InBus]		in_2_30_r;
reg signed [`InBus]		in_2_30_i;
reg signed [`InBus]		in_2_31_r;
reg signed [`InBus]		in_2_31_i;
reg signed [`InBus]		in_2_32_r;
reg signed [`InBus]		in_2_32_i;
reg signed [`InBus]		in_3_1_r;
reg signed [`InBus]		in_3_1_i;
reg signed [`InBus]		in_3_2_r;
reg signed [`InBus]		in_3_2_i;
reg signed [`InBus]		in_3_3_r;
reg signed [`InBus]		in_3_3_i;
reg signed [`InBus]		in_3_4_r;
reg signed [`InBus]		in_3_4_i;
reg signed [`InBus]		in_3_5_r;
reg signed [`InBus]		in_3_5_i;
reg signed [`InBus]		in_3_6_r;
reg signed [`InBus]		in_3_6_i;
reg signed [`InBus]		in_3_7_r;
reg signed [`InBus]		in_3_7_i;
reg signed [`InBus]		in_3_8_r;
reg signed [`InBus]		in_3_8_i;
reg signed [`InBus]		in_3_9_r;
reg signed [`InBus]		in_3_9_i;
reg signed [`InBus]		in_3_10_r;
reg signed [`InBus]		in_3_10_i;
reg signed [`InBus]		in_3_11_r;
reg signed [`InBus]		in_3_11_i;
reg signed [`InBus]		in_3_12_r;
reg signed [`InBus]		in_3_12_i;
reg signed [`InBus]		in_3_13_r;
reg signed [`InBus]		in_3_13_i;
reg signed [`InBus]		in_3_14_r;
reg signed [`InBus]		in_3_14_i;
reg signed [`InBus]		in_3_15_r;
reg signed [`InBus]		in_3_15_i;
reg signed [`InBus]		in_3_16_r;
reg signed [`InBus]		in_3_16_i;
reg signed [`InBus]		in_3_17_r;
reg signed [`InBus]		in_3_17_i;
reg signed [`InBus]		in_3_18_r;
reg signed [`InBus]		in_3_18_i;
reg signed [`InBus]		in_3_19_r;
reg signed [`InBus]		in_3_19_i;
reg signed [`InBus]		in_3_20_r;
reg signed [`InBus]		in_3_20_i;
reg signed [`InBus]		in_3_21_r;
reg signed [`InBus]		in_3_21_i;
reg signed [`InBus]		in_3_22_r;
reg signed [`InBus]		in_3_22_i;
reg signed [`InBus]		in_3_23_r;
reg signed [`InBus]		in_3_23_i;
reg signed [`InBus]		in_3_24_r;
reg signed [`InBus]		in_3_24_i;
reg signed [`InBus]		in_3_25_r;
reg signed [`InBus]		in_3_25_i;
reg signed [`InBus]		in_3_26_r;
reg signed [`InBus]		in_3_26_i;
reg signed [`InBus]		in_3_27_r;
reg signed [`InBus]		in_3_27_i;
reg signed [`InBus]		in_3_28_r;
reg signed [`InBus]		in_3_28_i;
reg signed [`InBus]		in_3_29_r;
reg signed [`InBus]		in_3_29_i;
reg signed [`InBus]		in_3_30_r;
reg signed [`InBus]		in_3_30_i;
reg signed [`InBus]		in_3_31_r;
reg signed [`InBus]		in_3_31_i;
reg signed [`InBus]		in_3_32_r;
reg signed [`InBus]		in_3_32_i;
reg signed [`InBus]		in_4_1_r;
reg signed [`InBus]		in_4_1_i;
reg signed [`InBus]		in_4_2_r;
reg signed [`InBus]		in_4_2_i;
reg signed [`InBus]		in_4_3_r;
reg signed [`InBus]		in_4_3_i;
reg signed [`InBus]		in_4_4_r;
reg signed [`InBus]		in_4_4_i;
reg signed [`InBus]		in_4_5_r;
reg signed [`InBus]		in_4_5_i;
reg signed [`InBus]		in_4_6_r;
reg signed [`InBus]		in_4_6_i;
reg signed [`InBus]		in_4_7_r;
reg signed [`InBus]		in_4_7_i;
reg signed [`InBus]		in_4_8_r;
reg signed [`InBus]		in_4_8_i;
reg signed [`InBus]		in_4_9_r;
reg signed [`InBus]		in_4_9_i;
reg signed [`InBus]		in_4_10_r;
reg signed [`InBus]		in_4_10_i;
reg signed [`InBus]		in_4_11_r;
reg signed [`InBus]		in_4_11_i;
reg signed [`InBus]		in_4_12_r;
reg signed [`InBus]		in_4_12_i;
reg signed [`InBus]		in_4_13_r;
reg signed [`InBus]		in_4_13_i;
reg signed [`InBus]		in_4_14_r;
reg signed [`InBus]		in_4_14_i;
reg signed [`InBus]		in_4_15_r;
reg signed [`InBus]		in_4_15_i;
reg signed [`InBus]		in_4_16_r;
reg signed [`InBus]		in_4_16_i;
reg signed [`InBus]		in_4_17_r;
reg signed [`InBus]		in_4_17_i;
reg signed [`InBus]		in_4_18_r;
reg signed [`InBus]		in_4_18_i;
reg signed [`InBus]		in_4_19_r;
reg signed [`InBus]		in_4_19_i;
reg signed [`InBus]		in_4_20_r;
reg signed [`InBus]		in_4_20_i;
reg signed [`InBus]		in_4_21_r;
reg signed [`InBus]		in_4_21_i;
reg signed [`InBus]		in_4_22_r;
reg signed [`InBus]		in_4_22_i;
reg signed [`InBus]		in_4_23_r;
reg signed [`InBus]		in_4_23_i;
reg signed [`InBus]		in_4_24_r;
reg signed [`InBus]		in_4_24_i;
reg signed [`InBus]		in_4_25_r;
reg signed [`InBus]		in_4_25_i;
reg signed [`InBus]		in_4_26_r;
reg signed [`InBus]		in_4_26_i;
reg signed [`InBus]		in_4_27_r;
reg signed [`InBus]		in_4_27_i;
reg signed [`InBus]		in_4_28_r;
reg signed [`InBus]		in_4_28_i;
reg signed [`InBus]		in_4_29_r;
reg signed [`InBus]		in_4_29_i;
reg signed [`InBus]		in_4_30_r;
reg signed [`InBus]		in_4_30_i;
reg signed [`InBus]		in_4_31_r;
reg signed [`InBus]		in_4_31_i;
reg signed [`InBus]		in_4_32_r;
reg signed [`InBus]		in_4_32_i;
reg signed [`InBus]		in_5_1_r;
reg signed [`InBus]		in_5_1_i;
reg signed [`InBus]		in_5_2_r;
reg signed [`InBus]		in_5_2_i;
reg signed [`InBus]		in_5_3_r;
reg signed [`InBus]		in_5_3_i;
reg signed [`InBus]		in_5_4_r;
reg signed [`InBus]		in_5_4_i;
reg signed [`InBus]		in_5_5_r;
reg signed [`InBus]		in_5_5_i;
reg signed [`InBus]		in_5_6_r;
reg signed [`InBus]		in_5_6_i;
reg signed [`InBus]		in_5_7_r;
reg signed [`InBus]		in_5_7_i;
reg signed [`InBus]		in_5_8_r;
reg signed [`InBus]		in_5_8_i;
reg signed [`InBus]		in_5_9_r;
reg signed [`InBus]		in_5_9_i;
reg signed [`InBus]		in_5_10_r;
reg signed [`InBus]		in_5_10_i;
reg signed [`InBus]		in_5_11_r;
reg signed [`InBus]		in_5_11_i;
reg signed [`InBus]		in_5_12_r;
reg signed [`InBus]		in_5_12_i;
reg signed [`InBus]		in_5_13_r;
reg signed [`InBus]		in_5_13_i;
reg signed [`InBus]		in_5_14_r;
reg signed [`InBus]		in_5_14_i;
reg signed [`InBus]		in_5_15_r;
reg signed [`InBus]		in_5_15_i;
reg signed [`InBus]		in_5_16_r;
reg signed [`InBus]		in_5_16_i;
reg signed [`InBus]		in_5_17_r;
reg signed [`InBus]		in_5_17_i;
reg signed [`InBus]		in_5_18_r;
reg signed [`InBus]		in_5_18_i;
reg signed [`InBus]		in_5_19_r;
reg signed [`InBus]		in_5_19_i;
reg signed [`InBus]		in_5_20_r;
reg signed [`InBus]		in_5_20_i;
reg signed [`InBus]		in_5_21_r;
reg signed [`InBus]		in_5_21_i;
reg signed [`InBus]		in_5_22_r;
reg signed [`InBus]		in_5_22_i;
reg signed [`InBus]		in_5_23_r;
reg signed [`InBus]		in_5_23_i;
reg signed [`InBus]		in_5_24_r;
reg signed [`InBus]		in_5_24_i;
reg signed [`InBus]		in_5_25_r;
reg signed [`InBus]		in_5_25_i;
reg signed [`InBus]		in_5_26_r;
reg signed [`InBus]		in_5_26_i;
reg signed [`InBus]		in_5_27_r;
reg signed [`InBus]		in_5_27_i;
reg signed [`InBus]		in_5_28_r;
reg signed [`InBus]		in_5_28_i;
reg signed [`InBus]		in_5_29_r;
reg signed [`InBus]		in_5_29_i;
reg signed [`InBus]		in_5_30_r;
reg signed [`InBus]		in_5_30_i;
reg signed [`InBus]		in_5_31_r;
reg signed [`InBus]		in_5_31_i;
reg signed [`InBus]		in_5_32_r;
reg signed [`InBus]		in_5_32_i;
reg signed [`InBus]		in_6_1_r;
reg signed [`InBus]		in_6_1_i;
reg signed [`InBus]		in_6_2_r;
reg signed [`InBus]		in_6_2_i;
reg signed [`InBus]		in_6_3_r;
reg signed [`InBus]		in_6_3_i;
reg signed [`InBus]		in_6_4_r;
reg signed [`InBus]		in_6_4_i;
reg signed [`InBus]		in_6_5_r;
reg signed [`InBus]		in_6_5_i;
reg signed [`InBus]		in_6_6_r;
reg signed [`InBus]		in_6_6_i;
reg signed [`InBus]		in_6_7_r;
reg signed [`InBus]		in_6_7_i;
reg signed [`InBus]		in_6_8_r;
reg signed [`InBus]		in_6_8_i;
reg signed [`InBus]		in_6_9_r;
reg signed [`InBus]		in_6_9_i;
reg signed [`InBus]		in_6_10_r;
reg signed [`InBus]		in_6_10_i;
reg signed [`InBus]		in_6_11_r;
reg signed [`InBus]		in_6_11_i;
reg signed [`InBus]		in_6_12_r;
reg signed [`InBus]		in_6_12_i;
reg signed [`InBus]		in_6_13_r;
reg signed [`InBus]		in_6_13_i;
reg signed [`InBus]		in_6_14_r;
reg signed [`InBus]		in_6_14_i;
reg signed [`InBus]		in_6_15_r;
reg signed [`InBus]		in_6_15_i;
reg signed [`InBus]		in_6_16_r;
reg signed [`InBus]		in_6_16_i;
reg signed [`InBus]		in_6_17_r;
reg signed [`InBus]		in_6_17_i;
reg signed [`InBus]		in_6_18_r;
reg signed [`InBus]		in_6_18_i;
reg signed [`InBus]		in_6_19_r;
reg signed [`InBus]		in_6_19_i;
reg signed [`InBus]		in_6_20_r;
reg signed [`InBus]		in_6_20_i;
reg signed [`InBus]		in_6_21_r;
reg signed [`InBus]		in_6_21_i;
reg signed [`InBus]		in_6_22_r;
reg signed [`InBus]		in_6_22_i;
reg signed [`InBus]		in_6_23_r;
reg signed [`InBus]		in_6_23_i;
reg signed [`InBus]		in_6_24_r;
reg signed [`InBus]		in_6_24_i;
reg signed [`InBus]		in_6_25_r;
reg signed [`InBus]		in_6_25_i;
reg signed [`InBus]		in_6_26_r;
reg signed [`InBus]		in_6_26_i;
reg signed [`InBus]		in_6_27_r;
reg signed [`InBus]		in_6_27_i;
reg signed [`InBus]		in_6_28_r;
reg signed [`InBus]		in_6_28_i;
reg signed [`InBus]		in_6_29_r;
reg signed [`InBus]		in_6_29_i;
reg signed [`InBus]		in_6_30_r;
reg signed [`InBus]		in_6_30_i;
reg signed [`InBus]		in_6_31_r;
reg signed [`InBus]		in_6_31_i;
reg signed [`InBus]		in_6_32_r;
reg signed [`InBus]		in_6_32_i;
reg signed [`InBus]		in_7_1_r;
reg signed [`InBus]		in_7_1_i;
reg signed [`InBus]		in_7_2_r;
reg signed [`InBus]		in_7_2_i;
reg signed [`InBus]		in_7_3_r;
reg signed [`InBus]		in_7_3_i;
reg signed [`InBus]		in_7_4_r;
reg signed [`InBus]		in_7_4_i;
reg signed [`InBus]		in_7_5_r;
reg signed [`InBus]		in_7_5_i;
reg signed [`InBus]		in_7_6_r;
reg signed [`InBus]		in_7_6_i;
reg signed [`InBus]		in_7_7_r;
reg signed [`InBus]		in_7_7_i;
reg signed [`InBus]		in_7_8_r;
reg signed [`InBus]		in_7_8_i;
reg signed [`InBus]		in_7_9_r;
reg signed [`InBus]		in_7_9_i;
reg signed [`InBus]		in_7_10_r;
reg signed [`InBus]		in_7_10_i;
reg signed [`InBus]		in_7_11_r;
reg signed [`InBus]		in_7_11_i;
reg signed [`InBus]		in_7_12_r;
reg signed [`InBus]		in_7_12_i;
reg signed [`InBus]		in_7_13_r;
reg signed [`InBus]		in_7_13_i;
reg signed [`InBus]		in_7_14_r;
reg signed [`InBus]		in_7_14_i;
reg signed [`InBus]		in_7_15_r;
reg signed [`InBus]		in_7_15_i;
reg signed [`InBus]		in_7_16_r;
reg signed [`InBus]		in_7_16_i;
reg signed [`InBus]		in_7_17_r;
reg signed [`InBus]		in_7_17_i;
reg signed [`InBus]		in_7_18_r;
reg signed [`InBus]		in_7_18_i;
reg signed [`InBus]		in_7_19_r;
reg signed [`InBus]		in_7_19_i;
reg signed [`InBus]		in_7_20_r;
reg signed [`InBus]		in_7_20_i;
reg signed [`InBus]		in_7_21_r;
reg signed [`InBus]		in_7_21_i;
reg signed [`InBus]		in_7_22_r;
reg signed [`InBus]		in_7_22_i;
reg signed [`InBus]		in_7_23_r;
reg signed [`InBus]		in_7_23_i;
reg signed [`InBus]		in_7_24_r;
reg signed [`InBus]		in_7_24_i;
reg signed [`InBus]		in_7_25_r;
reg signed [`InBus]		in_7_25_i;
reg signed [`InBus]		in_7_26_r;
reg signed [`InBus]		in_7_26_i;
reg signed [`InBus]		in_7_27_r;
reg signed [`InBus]		in_7_27_i;
reg signed [`InBus]		in_7_28_r;
reg signed [`InBus]		in_7_28_i;
reg signed [`InBus]		in_7_29_r;
reg signed [`InBus]		in_7_29_i;
reg signed [`InBus]		in_7_30_r;
reg signed [`InBus]		in_7_30_i;
reg signed [`InBus]		in_7_31_r;
reg signed [`InBus]		in_7_31_i;
reg signed [`InBus]		in_7_32_r;
reg signed [`InBus]		in_7_32_i;
reg signed [`InBus]		in_8_1_r;
reg signed [`InBus]		in_8_1_i;
reg signed [`InBus]		in_8_2_r;
reg signed [`InBus]		in_8_2_i;
reg signed [`InBus]		in_8_3_r;
reg signed [`InBus]		in_8_3_i;
reg signed [`InBus]		in_8_4_r;
reg signed [`InBus]		in_8_4_i;
reg signed [`InBus]		in_8_5_r;
reg signed [`InBus]		in_8_5_i;
reg signed [`InBus]		in_8_6_r;
reg signed [`InBus]		in_8_6_i;
reg signed [`InBus]		in_8_7_r;
reg signed [`InBus]		in_8_7_i;
reg signed [`InBus]		in_8_8_r;
reg signed [`InBus]		in_8_8_i;
reg signed [`InBus]		in_8_9_r;
reg signed [`InBus]		in_8_9_i;
reg signed [`InBus]		in_8_10_r;
reg signed [`InBus]		in_8_10_i;
reg signed [`InBus]		in_8_11_r;
reg signed [`InBus]		in_8_11_i;
reg signed [`InBus]		in_8_12_r;
reg signed [`InBus]		in_8_12_i;
reg signed [`InBus]		in_8_13_r;
reg signed [`InBus]		in_8_13_i;
reg signed [`InBus]		in_8_14_r;
reg signed [`InBus]		in_8_14_i;
reg signed [`InBus]		in_8_15_r;
reg signed [`InBus]		in_8_15_i;
reg signed [`InBus]		in_8_16_r;
reg signed [`InBus]		in_8_16_i;
reg signed [`InBus]		in_8_17_r;
reg signed [`InBus]		in_8_17_i;
reg signed [`InBus]		in_8_18_r;
reg signed [`InBus]		in_8_18_i;
reg signed [`InBus]		in_8_19_r;
reg signed [`InBus]		in_8_19_i;
reg signed [`InBus]		in_8_20_r;
reg signed [`InBus]		in_8_20_i;
reg signed [`InBus]		in_8_21_r;
reg signed [`InBus]		in_8_21_i;
reg signed [`InBus]		in_8_22_r;
reg signed [`InBus]		in_8_22_i;
reg signed [`InBus]		in_8_23_r;
reg signed [`InBus]		in_8_23_i;
reg signed [`InBus]		in_8_24_r;
reg signed [`InBus]		in_8_24_i;
reg signed [`InBus]		in_8_25_r;
reg signed [`InBus]		in_8_25_i;
reg signed [`InBus]		in_8_26_r;
reg signed [`InBus]		in_8_26_i;
reg signed [`InBus]		in_8_27_r;
reg signed [`InBus]		in_8_27_i;
reg signed [`InBus]		in_8_28_r;
reg signed [`InBus]		in_8_28_i;
reg signed [`InBus]		in_8_29_r;
reg signed [`InBus]		in_8_29_i;
reg signed [`InBus]		in_8_30_r;
reg signed [`InBus]		in_8_30_i;
reg signed [`InBus]		in_8_31_r;
reg signed [`InBus]		in_8_31_i;
reg signed [`InBus]		in_8_32_r;
reg signed [`InBus]		in_8_32_i;
reg signed [`InBus]		in_9_1_r;
reg signed [`InBus]		in_9_1_i;
reg signed [`InBus]		in_9_2_r;
reg signed [`InBus]		in_9_2_i;
reg signed [`InBus]		in_9_3_r;
reg signed [`InBus]		in_9_3_i;
reg signed [`InBus]		in_9_4_r;
reg signed [`InBus]		in_9_4_i;
reg signed [`InBus]		in_9_5_r;
reg signed [`InBus]		in_9_5_i;
reg signed [`InBus]		in_9_6_r;
reg signed [`InBus]		in_9_6_i;
reg signed [`InBus]		in_9_7_r;
reg signed [`InBus]		in_9_7_i;
reg signed [`InBus]		in_9_8_r;
reg signed [`InBus]		in_9_8_i;
reg signed [`InBus]		in_9_9_r;
reg signed [`InBus]		in_9_9_i;
reg signed [`InBus]		in_9_10_r;
reg signed [`InBus]		in_9_10_i;
reg signed [`InBus]		in_9_11_r;
reg signed [`InBus]		in_9_11_i;
reg signed [`InBus]		in_9_12_r;
reg signed [`InBus]		in_9_12_i;
reg signed [`InBus]		in_9_13_r;
reg signed [`InBus]		in_9_13_i;
reg signed [`InBus]		in_9_14_r;
reg signed [`InBus]		in_9_14_i;
reg signed [`InBus]		in_9_15_r;
reg signed [`InBus]		in_9_15_i;
reg signed [`InBus]		in_9_16_r;
reg signed [`InBus]		in_9_16_i;
reg signed [`InBus]		in_9_17_r;
reg signed [`InBus]		in_9_17_i;
reg signed [`InBus]		in_9_18_r;
reg signed [`InBus]		in_9_18_i;
reg signed [`InBus]		in_9_19_r;
reg signed [`InBus]		in_9_19_i;
reg signed [`InBus]		in_9_20_r;
reg signed [`InBus]		in_9_20_i;
reg signed [`InBus]		in_9_21_r;
reg signed [`InBus]		in_9_21_i;
reg signed [`InBus]		in_9_22_r;
reg signed [`InBus]		in_9_22_i;
reg signed [`InBus]		in_9_23_r;
reg signed [`InBus]		in_9_23_i;
reg signed [`InBus]		in_9_24_r;
reg signed [`InBus]		in_9_24_i;
reg signed [`InBus]		in_9_25_r;
reg signed [`InBus]		in_9_25_i;
reg signed [`InBus]		in_9_26_r;
reg signed [`InBus]		in_9_26_i;
reg signed [`InBus]		in_9_27_r;
reg signed [`InBus]		in_9_27_i;
reg signed [`InBus]		in_9_28_r;
reg signed [`InBus]		in_9_28_i;
reg signed [`InBus]		in_9_29_r;
reg signed [`InBus]		in_9_29_i;
reg signed [`InBus]		in_9_30_r;
reg signed [`InBus]		in_9_30_i;
reg signed [`InBus]		in_9_31_r;
reg signed [`InBus]		in_9_31_i;
reg signed [`InBus]		in_9_32_r;
reg signed [`InBus]		in_9_32_i;
reg signed [`InBus]		in_10_1_r;
reg signed [`InBus]		in_10_1_i;
reg signed [`InBus]		in_10_2_r;
reg signed [`InBus]		in_10_2_i;
reg signed [`InBus]		in_10_3_r;
reg signed [`InBus]		in_10_3_i;
reg signed [`InBus]		in_10_4_r;
reg signed [`InBus]		in_10_4_i;
reg signed [`InBus]		in_10_5_r;
reg signed [`InBus]		in_10_5_i;
reg signed [`InBus]		in_10_6_r;
reg signed [`InBus]		in_10_6_i;
reg signed [`InBus]		in_10_7_r;
reg signed [`InBus]		in_10_7_i;
reg signed [`InBus]		in_10_8_r;
reg signed [`InBus]		in_10_8_i;
reg signed [`InBus]		in_10_9_r;
reg signed [`InBus]		in_10_9_i;
reg signed [`InBus]		in_10_10_r;
reg signed [`InBus]		in_10_10_i;
reg signed [`InBus]		in_10_11_r;
reg signed [`InBus]		in_10_11_i;
reg signed [`InBus]		in_10_12_r;
reg signed [`InBus]		in_10_12_i;
reg signed [`InBus]		in_10_13_r;
reg signed [`InBus]		in_10_13_i;
reg signed [`InBus]		in_10_14_r;
reg signed [`InBus]		in_10_14_i;
reg signed [`InBus]		in_10_15_r;
reg signed [`InBus]		in_10_15_i;
reg signed [`InBus]		in_10_16_r;
reg signed [`InBus]		in_10_16_i;
reg signed [`InBus]		in_10_17_r;
reg signed [`InBus]		in_10_17_i;
reg signed [`InBus]		in_10_18_r;
reg signed [`InBus]		in_10_18_i;
reg signed [`InBus]		in_10_19_r;
reg signed [`InBus]		in_10_19_i;
reg signed [`InBus]		in_10_20_r;
reg signed [`InBus]		in_10_20_i;
reg signed [`InBus]		in_10_21_r;
reg signed [`InBus]		in_10_21_i;
reg signed [`InBus]		in_10_22_r;
reg signed [`InBus]		in_10_22_i;
reg signed [`InBus]		in_10_23_r;
reg signed [`InBus]		in_10_23_i;
reg signed [`InBus]		in_10_24_r;
reg signed [`InBus]		in_10_24_i;
reg signed [`InBus]		in_10_25_r;
reg signed [`InBus]		in_10_25_i;
reg signed [`InBus]		in_10_26_r;
reg signed [`InBus]		in_10_26_i;
reg signed [`InBus]		in_10_27_r;
reg signed [`InBus]		in_10_27_i;
reg signed [`InBus]		in_10_28_r;
reg signed [`InBus]		in_10_28_i;
reg signed [`InBus]		in_10_29_r;
reg signed [`InBus]		in_10_29_i;
reg signed [`InBus]		in_10_30_r;
reg signed [`InBus]		in_10_30_i;
reg signed [`InBus]		in_10_31_r;
reg signed [`InBus]		in_10_31_i;
reg signed [`InBus]		in_10_32_r;
reg signed [`InBus]		in_10_32_i;
reg signed [`InBus]		in_11_1_r;
reg signed [`InBus]		in_11_1_i;
reg signed [`InBus]		in_11_2_r;
reg signed [`InBus]		in_11_2_i;
reg signed [`InBus]		in_11_3_r;
reg signed [`InBus]		in_11_3_i;
reg signed [`InBus]		in_11_4_r;
reg signed [`InBus]		in_11_4_i;
reg signed [`InBus]		in_11_5_r;
reg signed [`InBus]		in_11_5_i;
reg signed [`InBus]		in_11_6_r;
reg signed [`InBus]		in_11_6_i;
reg signed [`InBus]		in_11_7_r;
reg signed [`InBus]		in_11_7_i;
reg signed [`InBus]		in_11_8_r;
reg signed [`InBus]		in_11_8_i;
reg signed [`InBus]		in_11_9_r;
reg signed [`InBus]		in_11_9_i;
reg signed [`InBus]		in_11_10_r;
reg signed [`InBus]		in_11_10_i;
reg signed [`InBus]		in_11_11_r;
reg signed [`InBus]		in_11_11_i;
reg signed [`InBus]		in_11_12_r;
reg signed [`InBus]		in_11_12_i;
reg signed [`InBus]		in_11_13_r;
reg signed [`InBus]		in_11_13_i;
reg signed [`InBus]		in_11_14_r;
reg signed [`InBus]		in_11_14_i;
reg signed [`InBus]		in_11_15_r;
reg signed [`InBus]		in_11_15_i;
reg signed [`InBus]		in_11_16_r;
reg signed [`InBus]		in_11_16_i;
reg signed [`InBus]		in_11_17_r;
reg signed [`InBus]		in_11_17_i;
reg signed [`InBus]		in_11_18_r;
reg signed [`InBus]		in_11_18_i;
reg signed [`InBus]		in_11_19_r;
reg signed [`InBus]		in_11_19_i;
reg signed [`InBus]		in_11_20_r;
reg signed [`InBus]		in_11_20_i;
reg signed [`InBus]		in_11_21_r;
reg signed [`InBus]		in_11_21_i;
reg signed [`InBus]		in_11_22_r;
reg signed [`InBus]		in_11_22_i;
reg signed [`InBus]		in_11_23_r;
reg signed [`InBus]		in_11_23_i;
reg signed [`InBus]		in_11_24_r;
reg signed [`InBus]		in_11_24_i;
reg signed [`InBus]		in_11_25_r;
reg signed [`InBus]		in_11_25_i;
reg signed [`InBus]		in_11_26_r;
reg signed [`InBus]		in_11_26_i;
reg signed [`InBus]		in_11_27_r;
reg signed [`InBus]		in_11_27_i;
reg signed [`InBus]		in_11_28_r;
reg signed [`InBus]		in_11_28_i;
reg signed [`InBus]		in_11_29_r;
reg signed [`InBus]		in_11_29_i;
reg signed [`InBus]		in_11_30_r;
reg signed [`InBus]		in_11_30_i;
reg signed [`InBus]		in_11_31_r;
reg signed [`InBus]		in_11_31_i;
reg signed [`InBus]		in_11_32_r;
reg signed [`InBus]		in_11_32_i;
reg signed [`InBus]		in_12_1_r;
reg signed [`InBus]		in_12_1_i;
reg signed [`InBus]		in_12_2_r;
reg signed [`InBus]		in_12_2_i;
reg signed [`InBus]		in_12_3_r;
reg signed [`InBus]		in_12_3_i;
reg signed [`InBus]		in_12_4_r;
reg signed [`InBus]		in_12_4_i;
reg signed [`InBus]		in_12_5_r;
reg signed [`InBus]		in_12_5_i;
reg signed [`InBus]		in_12_6_r;
reg signed [`InBus]		in_12_6_i;
reg signed [`InBus]		in_12_7_r;
reg signed [`InBus]		in_12_7_i;
reg signed [`InBus]		in_12_8_r;
reg signed [`InBus]		in_12_8_i;
reg signed [`InBus]		in_12_9_r;
reg signed [`InBus]		in_12_9_i;
reg signed [`InBus]		in_12_10_r;
reg signed [`InBus]		in_12_10_i;
reg signed [`InBus]		in_12_11_r;
reg signed [`InBus]		in_12_11_i;
reg signed [`InBus]		in_12_12_r;
reg signed [`InBus]		in_12_12_i;
reg signed [`InBus]		in_12_13_r;
reg signed [`InBus]		in_12_13_i;
reg signed [`InBus]		in_12_14_r;
reg signed [`InBus]		in_12_14_i;
reg signed [`InBus]		in_12_15_r;
reg signed [`InBus]		in_12_15_i;
reg signed [`InBus]		in_12_16_r;
reg signed [`InBus]		in_12_16_i;
reg signed [`InBus]		in_12_17_r;
reg signed [`InBus]		in_12_17_i;
reg signed [`InBus]		in_12_18_r;
reg signed [`InBus]		in_12_18_i;
reg signed [`InBus]		in_12_19_r;
reg signed [`InBus]		in_12_19_i;
reg signed [`InBus]		in_12_20_r;
reg signed [`InBus]		in_12_20_i;
reg signed [`InBus]		in_12_21_r;
reg signed [`InBus]		in_12_21_i;
reg signed [`InBus]		in_12_22_r;
reg signed [`InBus]		in_12_22_i;
reg signed [`InBus]		in_12_23_r;
reg signed [`InBus]		in_12_23_i;
reg signed [`InBus]		in_12_24_r;
reg signed [`InBus]		in_12_24_i;
reg signed [`InBus]		in_12_25_r;
reg signed [`InBus]		in_12_25_i;
reg signed [`InBus]		in_12_26_r;
reg signed [`InBus]		in_12_26_i;
reg signed [`InBus]		in_12_27_r;
reg signed [`InBus]		in_12_27_i;
reg signed [`InBus]		in_12_28_r;
reg signed [`InBus]		in_12_28_i;
reg signed [`InBus]		in_12_29_r;
reg signed [`InBus]		in_12_29_i;
reg signed [`InBus]		in_12_30_r;
reg signed [`InBus]		in_12_30_i;
reg signed [`InBus]		in_12_31_r;
reg signed [`InBus]		in_12_31_i;
reg signed [`InBus]		in_12_32_r;
reg signed [`InBus]		in_12_32_i;
reg signed [`InBus]		in_13_1_r;
reg signed [`InBus]		in_13_1_i;
reg signed [`InBus]		in_13_2_r;
reg signed [`InBus]		in_13_2_i;
reg signed [`InBus]		in_13_3_r;
reg signed [`InBus]		in_13_3_i;
reg signed [`InBus]		in_13_4_r;
reg signed [`InBus]		in_13_4_i;
reg signed [`InBus]		in_13_5_r;
reg signed [`InBus]		in_13_5_i;
reg signed [`InBus]		in_13_6_r;
reg signed [`InBus]		in_13_6_i;
reg signed [`InBus]		in_13_7_r;
reg signed [`InBus]		in_13_7_i;
reg signed [`InBus]		in_13_8_r;
reg signed [`InBus]		in_13_8_i;
reg signed [`InBus]		in_13_9_r;
reg signed [`InBus]		in_13_9_i;
reg signed [`InBus]		in_13_10_r;
reg signed [`InBus]		in_13_10_i;
reg signed [`InBus]		in_13_11_r;
reg signed [`InBus]		in_13_11_i;
reg signed [`InBus]		in_13_12_r;
reg signed [`InBus]		in_13_12_i;
reg signed [`InBus]		in_13_13_r;
reg signed [`InBus]		in_13_13_i;
reg signed [`InBus]		in_13_14_r;
reg signed [`InBus]		in_13_14_i;
reg signed [`InBus]		in_13_15_r;
reg signed [`InBus]		in_13_15_i;
reg signed [`InBus]		in_13_16_r;
reg signed [`InBus]		in_13_16_i;
reg signed [`InBus]		in_13_17_r;
reg signed [`InBus]		in_13_17_i;
reg signed [`InBus]		in_13_18_r;
reg signed [`InBus]		in_13_18_i;
reg signed [`InBus]		in_13_19_r;
reg signed [`InBus]		in_13_19_i;
reg signed [`InBus]		in_13_20_r;
reg signed [`InBus]		in_13_20_i;
reg signed [`InBus]		in_13_21_r;
reg signed [`InBus]		in_13_21_i;
reg signed [`InBus]		in_13_22_r;
reg signed [`InBus]		in_13_22_i;
reg signed [`InBus]		in_13_23_r;
reg signed [`InBus]		in_13_23_i;
reg signed [`InBus]		in_13_24_r;
reg signed [`InBus]		in_13_24_i;
reg signed [`InBus]		in_13_25_r;
reg signed [`InBus]		in_13_25_i;
reg signed [`InBus]		in_13_26_r;
reg signed [`InBus]		in_13_26_i;
reg signed [`InBus]		in_13_27_r;
reg signed [`InBus]		in_13_27_i;
reg signed [`InBus]		in_13_28_r;
reg signed [`InBus]		in_13_28_i;
reg signed [`InBus]		in_13_29_r;
reg signed [`InBus]		in_13_29_i;
reg signed [`InBus]		in_13_30_r;
reg signed [`InBus]		in_13_30_i;
reg signed [`InBus]		in_13_31_r;
reg signed [`InBus]		in_13_31_i;
reg signed [`InBus]		in_13_32_r;
reg signed [`InBus]		in_13_32_i;
reg signed [`InBus]		in_14_1_r;
reg signed [`InBus]		in_14_1_i;
reg signed [`InBus]		in_14_2_r;
reg signed [`InBus]		in_14_2_i;
reg signed [`InBus]		in_14_3_r;
reg signed [`InBus]		in_14_3_i;
reg signed [`InBus]		in_14_4_r;
reg signed [`InBus]		in_14_4_i;
reg signed [`InBus]		in_14_5_r;
reg signed [`InBus]		in_14_5_i;
reg signed [`InBus]		in_14_6_r;
reg signed [`InBus]		in_14_6_i;
reg signed [`InBus]		in_14_7_r;
reg signed [`InBus]		in_14_7_i;
reg signed [`InBus]		in_14_8_r;
reg signed [`InBus]		in_14_8_i;
reg signed [`InBus]		in_14_9_r;
reg signed [`InBus]		in_14_9_i;
reg signed [`InBus]		in_14_10_r;
reg signed [`InBus]		in_14_10_i;
reg signed [`InBus]		in_14_11_r;
reg signed [`InBus]		in_14_11_i;
reg signed [`InBus]		in_14_12_r;
reg signed [`InBus]		in_14_12_i;
reg signed [`InBus]		in_14_13_r;
reg signed [`InBus]		in_14_13_i;
reg signed [`InBus]		in_14_14_r;
reg signed [`InBus]		in_14_14_i;
reg signed [`InBus]		in_14_15_r;
reg signed [`InBus]		in_14_15_i;
reg signed [`InBus]		in_14_16_r;
reg signed [`InBus]		in_14_16_i;
reg signed [`InBus]		in_14_17_r;
reg signed [`InBus]		in_14_17_i;
reg signed [`InBus]		in_14_18_r;
reg signed [`InBus]		in_14_18_i;
reg signed [`InBus]		in_14_19_r;
reg signed [`InBus]		in_14_19_i;
reg signed [`InBus]		in_14_20_r;
reg signed [`InBus]		in_14_20_i;
reg signed [`InBus]		in_14_21_r;
reg signed [`InBus]		in_14_21_i;
reg signed [`InBus]		in_14_22_r;
reg signed [`InBus]		in_14_22_i;
reg signed [`InBus]		in_14_23_r;
reg signed [`InBus]		in_14_23_i;
reg signed [`InBus]		in_14_24_r;
reg signed [`InBus]		in_14_24_i;
reg signed [`InBus]		in_14_25_r;
reg signed [`InBus]		in_14_25_i;
reg signed [`InBus]		in_14_26_r;
reg signed [`InBus]		in_14_26_i;
reg signed [`InBus]		in_14_27_r;
reg signed [`InBus]		in_14_27_i;
reg signed [`InBus]		in_14_28_r;
reg signed [`InBus]		in_14_28_i;
reg signed [`InBus]		in_14_29_r;
reg signed [`InBus]		in_14_29_i;
reg signed [`InBus]		in_14_30_r;
reg signed [`InBus]		in_14_30_i;
reg signed [`InBus]		in_14_31_r;
reg signed [`InBus]		in_14_31_i;
reg signed [`InBus]		in_14_32_r;
reg signed [`InBus]		in_14_32_i;
reg signed [`InBus]		in_15_1_r;
reg signed [`InBus]		in_15_1_i;
reg signed [`InBus]		in_15_2_r;
reg signed [`InBus]		in_15_2_i;
reg signed [`InBus]		in_15_3_r;
reg signed [`InBus]		in_15_3_i;
reg signed [`InBus]		in_15_4_r;
reg signed [`InBus]		in_15_4_i;
reg signed [`InBus]		in_15_5_r;
reg signed [`InBus]		in_15_5_i;
reg signed [`InBus]		in_15_6_r;
reg signed [`InBus]		in_15_6_i;
reg signed [`InBus]		in_15_7_r;
reg signed [`InBus]		in_15_7_i;
reg signed [`InBus]		in_15_8_r;
reg signed [`InBus]		in_15_8_i;
reg signed [`InBus]		in_15_9_r;
reg signed [`InBus]		in_15_9_i;
reg signed [`InBus]		in_15_10_r;
reg signed [`InBus]		in_15_10_i;
reg signed [`InBus]		in_15_11_r;
reg signed [`InBus]		in_15_11_i;
reg signed [`InBus]		in_15_12_r;
reg signed [`InBus]		in_15_12_i;
reg signed [`InBus]		in_15_13_r;
reg signed [`InBus]		in_15_13_i;
reg signed [`InBus]		in_15_14_r;
reg signed [`InBus]		in_15_14_i;
reg signed [`InBus]		in_15_15_r;
reg signed [`InBus]		in_15_15_i;
reg signed [`InBus]		in_15_16_r;
reg signed [`InBus]		in_15_16_i;
reg signed [`InBus]		in_15_17_r;
reg signed [`InBus]		in_15_17_i;
reg signed [`InBus]		in_15_18_r;
reg signed [`InBus]		in_15_18_i;
reg signed [`InBus]		in_15_19_r;
reg signed [`InBus]		in_15_19_i;
reg signed [`InBus]		in_15_20_r;
reg signed [`InBus]		in_15_20_i;
reg signed [`InBus]		in_15_21_r;
reg signed [`InBus]		in_15_21_i;
reg signed [`InBus]		in_15_22_r;
reg signed [`InBus]		in_15_22_i;
reg signed [`InBus]		in_15_23_r;
reg signed [`InBus]		in_15_23_i;
reg signed [`InBus]		in_15_24_r;
reg signed [`InBus]		in_15_24_i;
reg signed [`InBus]		in_15_25_r;
reg signed [`InBus]		in_15_25_i;
reg signed [`InBus]		in_15_26_r;
reg signed [`InBus]		in_15_26_i;
reg signed [`InBus]		in_15_27_r;
reg signed [`InBus]		in_15_27_i;
reg signed [`InBus]		in_15_28_r;
reg signed [`InBus]		in_15_28_i;
reg signed [`InBus]		in_15_29_r;
reg signed [`InBus]		in_15_29_i;
reg signed [`InBus]		in_15_30_r;
reg signed [`InBus]		in_15_30_i;
reg signed [`InBus]		in_15_31_r;
reg signed [`InBus]		in_15_31_i;
reg signed [`InBus]		in_15_32_r;
reg signed [`InBus]		in_15_32_i;
reg signed [`InBus]		in_16_1_r;
reg signed [`InBus]		in_16_1_i;
reg signed [`InBus]		in_16_2_r;
reg signed [`InBus]		in_16_2_i;
reg signed [`InBus]		in_16_3_r;
reg signed [`InBus]		in_16_3_i;
reg signed [`InBus]		in_16_4_r;
reg signed [`InBus]		in_16_4_i;
reg signed [`InBus]		in_16_5_r;
reg signed [`InBus]		in_16_5_i;
reg signed [`InBus]		in_16_6_r;
reg signed [`InBus]		in_16_6_i;
reg signed [`InBus]		in_16_7_r;
reg signed [`InBus]		in_16_7_i;
reg signed [`InBus]		in_16_8_r;
reg signed [`InBus]		in_16_8_i;
reg signed [`InBus]		in_16_9_r;
reg signed [`InBus]		in_16_9_i;
reg signed [`InBus]		in_16_10_r;
reg signed [`InBus]		in_16_10_i;
reg signed [`InBus]		in_16_11_r;
reg signed [`InBus]		in_16_11_i;
reg signed [`InBus]		in_16_12_r;
reg signed [`InBus]		in_16_12_i;
reg signed [`InBus]		in_16_13_r;
reg signed [`InBus]		in_16_13_i;
reg signed [`InBus]		in_16_14_r;
reg signed [`InBus]		in_16_14_i;
reg signed [`InBus]		in_16_15_r;
reg signed [`InBus]		in_16_15_i;
reg signed [`InBus]		in_16_16_r;
reg signed [`InBus]		in_16_16_i;
reg signed [`InBus]		in_16_17_r;
reg signed [`InBus]		in_16_17_i;
reg signed [`InBus]		in_16_18_r;
reg signed [`InBus]		in_16_18_i;
reg signed [`InBus]		in_16_19_r;
reg signed [`InBus]		in_16_19_i;
reg signed [`InBus]		in_16_20_r;
reg signed [`InBus]		in_16_20_i;
reg signed [`InBus]		in_16_21_r;
reg signed [`InBus]		in_16_21_i;
reg signed [`InBus]		in_16_22_r;
reg signed [`InBus]		in_16_22_i;
reg signed [`InBus]		in_16_23_r;
reg signed [`InBus]		in_16_23_i;
reg signed [`InBus]		in_16_24_r;
reg signed [`InBus]		in_16_24_i;
reg signed [`InBus]		in_16_25_r;
reg signed [`InBus]		in_16_25_i;
reg signed [`InBus]		in_16_26_r;
reg signed [`InBus]		in_16_26_i;
reg signed [`InBus]		in_16_27_r;
reg signed [`InBus]		in_16_27_i;
reg signed [`InBus]		in_16_28_r;
reg signed [`InBus]		in_16_28_i;
reg signed [`InBus]		in_16_29_r;
reg signed [`InBus]		in_16_29_i;
reg signed [`InBus]		in_16_30_r;
reg signed [`InBus]		in_16_30_i;
reg signed [`InBus]		in_16_31_r;
reg signed [`InBus]		in_16_31_i;
reg signed [`InBus]		in_16_32_r;
reg signed [`InBus]		in_16_32_i;
reg signed [`InBus]		in_17_1_r;
reg signed [`InBus]		in_17_1_i;
reg signed [`InBus]		in_17_2_r;
reg signed [`InBus]		in_17_2_i;
reg signed [`InBus]		in_17_3_r;
reg signed [`InBus]		in_17_3_i;
reg signed [`InBus]		in_17_4_r;
reg signed [`InBus]		in_17_4_i;
reg signed [`InBus]		in_17_5_r;
reg signed [`InBus]		in_17_5_i;
reg signed [`InBus]		in_17_6_r;
reg signed [`InBus]		in_17_6_i;
reg signed [`InBus]		in_17_7_r;
reg signed [`InBus]		in_17_7_i;
reg signed [`InBus]		in_17_8_r;
reg signed [`InBus]		in_17_8_i;
reg signed [`InBus]		in_17_9_r;
reg signed [`InBus]		in_17_9_i;
reg signed [`InBus]		in_17_10_r;
reg signed [`InBus]		in_17_10_i;
reg signed [`InBus]		in_17_11_r;
reg signed [`InBus]		in_17_11_i;
reg signed [`InBus]		in_17_12_r;
reg signed [`InBus]		in_17_12_i;
reg signed [`InBus]		in_17_13_r;
reg signed [`InBus]		in_17_13_i;
reg signed [`InBus]		in_17_14_r;
reg signed [`InBus]		in_17_14_i;
reg signed [`InBus]		in_17_15_r;
reg signed [`InBus]		in_17_15_i;
reg signed [`InBus]		in_17_16_r;
reg signed [`InBus]		in_17_16_i;
reg signed [`InBus]		in_17_17_r;
reg signed [`InBus]		in_17_17_i;
reg signed [`InBus]		in_17_18_r;
reg signed [`InBus]		in_17_18_i;
reg signed [`InBus]		in_17_19_r;
reg signed [`InBus]		in_17_19_i;
reg signed [`InBus]		in_17_20_r;
reg signed [`InBus]		in_17_20_i;
reg signed [`InBus]		in_17_21_r;
reg signed [`InBus]		in_17_21_i;
reg signed [`InBus]		in_17_22_r;
reg signed [`InBus]		in_17_22_i;
reg signed [`InBus]		in_17_23_r;
reg signed [`InBus]		in_17_23_i;
reg signed [`InBus]		in_17_24_r;
reg signed [`InBus]		in_17_24_i;
reg signed [`InBus]		in_17_25_r;
reg signed [`InBus]		in_17_25_i;
reg signed [`InBus]		in_17_26_r;
reg signed [`InBus]		in_17_26_i;
reg signed [`InBus]		in_17_27_r;
reg signed [`InBus]		in_17_27_i;
reg signed [`InBus]		in_17_28_r;
reg signed [`InBus]		in_17_28_i;
reg signed [`InBus]		in_17_29_r;
reg signed [`InBus]		in_17_29_i;
reg signed [`InBus]		in_17_30_r;
reg signed [`InBus]		in_17_30_i;
reg signed [`InBus]		in_17_31_r;
reg signed [`InBus]		in_17_31_i;
reg signed [`InBus]		in_17_32_r;
reg signed [`InBus]		in_17_32_i;
reg signed [`InBus]		in_18_1_r;
reg signed [`InBus]		in_18_1_i;
reg signed [`InBus]		in_18_2_r;
reg signed [`InBus]		in_18_2_i;
reg signed [`InBus]		in_18_3_r;
reg signed [`InBus]		in_18_3_i;
reg signed [`InBus]		in_18_4_r;
reg signed [`InBus]		in_18_4_i;
reg signed [`InBus]		in_18_5_r;
reg signed [`InBus]		in_18_5_i;
reg signed [`InBus]		in_18_6_r;
reg signed [`InBus]		in_18_6_i;
reg signed [`InBus]		in_18_7_r;
reg signed [`InBus]		in_18_7_i;
reg signed [`InBus]		in_18_8_r;
reg signed [`InBus]		in_18_8_i;
reg signed [`InBus]		in_18_9_r;
reg signed [`InBus]		in_18_9_i;
reg signed [`InBus]		in_18_10_r;
reg signed [`InBus]		in_18_10_i;
reg signed [`InBus]		in_18_11_r;
reg signed [`InBus]		in_18_11_i;
reg signed [`InBus]		in_18_12_r;
reg signed [`InBus]		in_18_12_i;
reg signed [`InBus]		in_18_13_r;
reg signed [`InBus]		in_18_13_i;
reg signed [`InBus]		in_18_14_r;
reg signed [`InBus]		in_18_14_i;
reg signed [`InBus]		in_18_15_r;
reg signed [`InBus]		in_18_15_i;
reg signed [`InBus]		in_18_16_r;
reg signed [`InBus]		in_18_16_i;
reg signed [`InBus]		in_18_17_r;
reg signed [`InBus]		in_18_17_i;
reg signed [`InBus]		in_18_18_r;
reg signed [`InBus]		in_18_18_i;
reg signed [`InBus]		in_18_19_r;
reg signed [`InBus]		in_18_19_i;
reg signed [`InBus]		in_18_20_r;
reg signed [`InBus]		in_18_20_i;
reg signed [`InBus]		in_18_21_r;
reg signed [`InBus]		in_18_21_i;
reg signed [`InBus]		in_18_22_r;
reg signed [`InBus]		in_18_22_i;
reg signed [`InBus]		in_18_23_r;
reg signed [`InBus]		in_18_23_i;
reg signed [`InBus]		in_18_24_r;
reg signed [`InBus]		in_18_24_i;
reg signed [`InBus]		in_18_25_r;
reg signed [`InBus]		in_18_25_i;
reg signed [`InBus]		in_18_26_r;
reg signed [`InBus]		in_18_26_i;
reg signed [`InBus]		in_18_27_r;
reg signed [`InBus]		in_18_27_i;
reg signed [`InBus]		in_18_28_r;
reg signed [`InBus]		in_18_28_i;
reg signed [`InBus]		in_18_29_r;
reg signed [`InBus]		in_18_29_i;
reg signed [`InBus]		in_18_30_r;
reg signed [`InBus]		in_18_30_i;
reg signed [`InBus]		in_18_31_r;
reg signed [`InBus]		in_18_31_i;
reg signed [`InBus]		in_18_32_r;
reg signed [`InBus]		in_18_32_i;
reg signed [`InBus]		in_19_1_r;
reg signed [`InBus]		in_19_1_i;
reg signed [`InBus]		in_19_2_r;
reg signed [`InBus]		in_19_2_i;
reg signed [`InBus]		in_19_3_r;
reg signed [`InBus]		in_19_3_i;
reg signed [`InBus]		in_19_4_r;
reg signed [`InBus]		in_19_4_i;
reg signed [`InBus]		in_19_5_r;
reg signed [`InBus]		in_19_5_i;
reg signed [`InBus]		in_19_6_r;
reg signed [`InBus]		in_19_6_i;
reg signed [`InBus]		in_19_7_r;
reg signed [`InBus]		in_19_7_i;
reg signed [`InBus]		in_19_8_r;
reg signed [`InBus]		in_19_8_i;
reg signed [`InBus]		in_19_9_r;
reg signed [`InBus]		in_19_9_i;
reg signed [`InBus]		in_19_10_r;
reg signed [`InBus]		in_19_10_i;
reg signed [`InBus]		in_19_11_r;
reg signed [`InBus]		in_19_11_i;
reg signed [`InBus]		in_19_12_r;
reg signed [`InBus]		in_19_12_i;
reg signed [`InBus]		in_19_13_r;
reg signed [`InBus]		in_19_13_i;
reg signed [`InBus]		in_19_14_r;
reg signed [`InBus]		in_19_14_i;
reg signed [`InBus]		in_19_15_r;
reg signed [`InBus]		in_19_15_i;
reg signed [`InBus]		in_19_16_r;
reg signed [`InBus]		in_19_16_i;
reg signed [`InBus]		in_19_17_r;
reg signed [`InBus]		in_19_17_i;
reg signed [`InBus]		in_19_18_r;
reg signed [`InBus]		in_19_18_i;
reg signed [`InBus]		in_19_19_r;
reg signed [`InBus]		in_19_19_i;
reg signed [`InBus]		in_19_20_r;
reg signed [`InBus]		in_19_20_i;
reg signed [`InBus]		in_19_21_r;
reg signed [`InBus]		in_19_21_i;
reg signed [`InBus]		in_19_22_r;
reg signed [`InBus]		in_19_22_i;
reg signed [`InBus]		in_19_23_r;
reg signed [`InBus]		in_19_23_i;
reg signed [`InBus]		in_19_24_r;
reg signed [`InBus]		in_19_24_i;
reg signed [`InBus]		in_19_25_r;
reg signed [`InBus]		in_19_25_i;
reg signed [`InBus]		in_19_26_r;
reg signed [`InBus]		in_19_26_i;
reg signed [`InBus]		in_19_27_r;
reg signed [`InBus]		in_19_27_i;
reg signed [`InBus]		in_19_28_r;
reg signed [`InBus]		in_19_28_i;
reg signed [`InBus]		in_19_29_r;
reg signed [`InBus]		in_19_29_i;
reg signed [`InBus]		in_19_30_r;
reg signed [`InBus]		in_19_30_i;
reg signed [`InBus]		in_19_31_r;
reg signed [`InBus]		in_19_31_i;
reg signed [`InBus]		in_19_32_r;
reg signed [`InBus]		in_19_32_i;
reg signed [`InBus]		in_20_1_r;
reg signed [`InBus]		in_20_1_i;
reg signed [`InBus]		in_20_2_r;
reg signed [`InBus]		in_20_2_i;
reg signed [`InBus]		in_20_3_r;
reg signed [`InBus]		in_20_3_i;
reg signed [`InBus]		in_20_4_r;
reg signed [`InBus]		in_20_4_i;
reg signed [`InBus]		in_20_5_r;
reg signed [`InBus]		in_20_5_i;
reg signed [`InBus]		in_20_6_r;
reg signed [`InBus]		in_20_6_i;
reg signed [`InBus]		in_20_7_r;
reg signed [`InBus]		in_20_7_i;
reg signed [`InBus]		in_20_8_r;
reg signed [`InBus]		in_20_8_i;
reg signed [`InBus]		in_20_9_r;
reg signed [`InBus]		in_20_9_i;
reg signed [`InBus]		in_20_10_r;
reg signed [`InBus]		in_20_10_i;
reg signed [`InBus]		in_20_11_r;
reg signed [`InBus]		in_20_11_i;
reg signed [`InBus]		in_20_12_r;
reg signed [`InBus]		in_20_12_i;
reg signed [`InBus]		in_20_13_r;
reg signed [`InBus]		in_20_13_i;
reg signed [`InBus]		in_20_14_r;
reg signed [`InBus]		in_20_14_i;
reg signed [`InBus]		in_20_15_r;
reg signed [`InBus]		in_20_15_i;
reg signed [`InBus]		in_20_16_r;
reg signed [`InBus]		in_20_16_i;
reg signed [`InBus]		in_20_17_r;
reg signed [`InBus]		in_20_17_i;
reg signed [`InBus]		in_20_18_r;
reg signed [`InBus]		in_20_18_i;
reg signed [`InBus]		in_20_19_r;
reg signed [`InBus]		in_20_19_i;
reg signed [`InBus]		in_20_20_r;
reg signed [`InBus]		in_20_20_i;
reg signed [`InBus]		in_20_21_r;
reg signed [`InBus]		in_20_21_i;
reg signed [`InBus]		in_20_22_r;
reg signed [`InBus]		in_20_22_i;
reg signed [`InBus]		in_20_23_r;
reg signed [`InBus]		in_20_23_i;
reg signed [`InBus]		in_20_24_r;
reg signed [`InBus]		in_20_24_i;
reg signed [`InBus]		in_20_25_r;
reg signed [`InBus]		in_20_25_i;
reg signed [`InBus]		in_20_26_r;
reg signed [`InBus]		in_20_26_i;
reg signed [`InBus]		in_20_27_r;
reg signed [`InBus]		in_20_27_i;
reg signed [`InBus]		in_20_28_r;
reg signed [`InBus]		in_20_28_i;
reg signed [`InBus]		in_20_29_r;
reg signed [`InBus]		in_20_29_i;
reg signed [`InBus]		in_20_30_r;
reg signed [`InBus]		in_20_30_i;
reg signed [`InBus]		in_20_31_r;
reg signed [`InBus]		in_20_31_i;
reg signed [`InBus]		in_20_32_r;
reg signed [`InBus]		in_20_32_i;
reg signed [`InBus]		in_21_1_r;
reg signed [`InBus]		in_21_1_i;
reg signed [`InBus]		in_21_2_r;
reg signed [`InBus]		in_21_2_i;
reg signed [`InBus]		in_21_3_r;
reg signed [`InBus]		in_21_3_i;
reg signed [`InBus]		in_21_4_r;
reg signed [`InBus]		in_21_4_i;
reg signed [`InBus]		in_21_5_r;
reg signed [`InBus]		in_21_5_i;
reg signed [`InBus]		in_21_6_r;
reg signed [`InBus]		in_21_6_i;
reg signed [`InBus]		in_21_7_r;
reg signed [`InBus]		in_21_7_i;
reg signed [`InBus]		in_21_8_r;
reg signed [`InBus]		in_21_8_i;
reg signed [`InBus]		in_21_9_r;
reg signed [`InBus]		in_21_9_i;
reg signed [`InBus]		in_21_10_r;
reg signed [`InBus]		in_21_10_i;
reg signed [`InBus]		in_21_11_r;
reg signed [`InBus]		in_21_11_i;
reg signed [`InBus]		in_21_12_r;
reg signed [`InBus]		in_21_12_i;
reg signed [`InBus]		in_21_13_r;
reg signed [`InBus]		in_21_13_i;
reg signed [`InBus]		in_21_14_r;
reg signed [`InBus]		in_21_14_i;
reg signed [`InBus]		in_21_15_r;
reg signed [`InBus]		in_21_15_i;
reg signed [`InBus]		in_21_16_r;
reg signed [`InBus]		in_21_16_i;
reg signed [`InBus]		in_21_17_r;
reg signed [`InBus]		in_21_17_i;
reg signed [`InBus]		in_21_18_r;
reg signed [`InBus]		in_21_18_i;
reg signed [`InBus]		in_21_19_r;
reg signed [`InBus]		in_21_19_i;
reg signed [`InBus]		in_21_20_r;
reg signed [`InBus]		in_21_20_i;
reg signed [`InBus]		in_21_21_r;
reg signed [`InBus]		in_21_21_i;
reg signed [`InBus]		in_21_22_r;
reg signed [`InBus]		in_21_22_i;
reg signed [`InBus]		in_21_23_r;
reg signed [`InBus]		in_21_23_i;
reg signed [`InBus]		in_21_24_r;
reg signed [`InBus]		in_21_24_i;
reg signed [`InBus]		in_21_25_r;
reg signed [`InBus]		in_21_25_i;
reg signed [`InBus]		in_21_26_r;
reg signed [`InBus]		in_21_26_i;
reg signed [`InBus]		in_21_27_r;
reg signed [`InBus]		in_21_27_i;
reg signed [`InBus]		in_21_28_r;
reg signed [`InBus]		in_21_28_i;
reg signed [`InBus]		in_21_29_r;
reg signed [`InBus]		in_21_29_i;
reg signed [`InBus]		in_21_30_r;
reg signed [`InBus]		in_21_30_i;
reg signed [`InBus]		in_21_31_r;
reg signed [`InBus]		in_21_31_i;
reg signed [`InBus]		in_21_32_r;
reg signed [`InBus]		in_21_32_i;
reg signed [`InBus]		in_22_1_r;
reg signed [`InBus]		in_22_1_i;
reg signed [`InBus]		in_22_2_r;
reg signed [`InBus]		in_22_2_i;
reg signed [`InBus]		in_22_3_r;
reg signed [`InBus]		in_22_3_i;
reg signed [`InBus]		in_22_4_r;
reg signed [`InBus]		in_22_4_i;
reg signed [`InBus]		in_22_5_r;
reg signed [`InBus]		in_22_5_i;
reg signed [`InBus]		in_22_6_r;
reg signed [`InBus]		in_22_6_i;
reg signed [`InBus]		in_22_7_r;
reg signed [`InBus]		in_22_7_i;
reg signed [`InBus]		in_22_8_r;
reg signed [`InBus]		in_22_8_i;
reg signed [`InBus]		in_22_9_r;
reg signed [`InBus]		in_22_9_i;
reg signed [`InBus]		in_22_10_r;
reg signed [`InBus]		in_22_10_i;
reg signed [`InBus]		in_22_11_r;
reg signed [`InBus]		in_22_11_i;
reg signed [`InBus]		in_22_12_r;
reg signed [`InBus]		in_22_12_i;
reg signed [`InBus]		in_22_13_r;
reg signed [`InBus]		in_22_13_i;
reg signed [`InBus]		in_22_14_r;
reg signed [`InBus]		in_22_14_i;
reg signed [`InBus]		in_22_15_r;
reg signed [`InBus]		in_22_15_i;
reg signed [`InBus]		in_22_16_r;
reg signed [`InBus]		in_22_16_i;
reg signed [`InBus]		in_22_17_r;
reg signed [`InBus]		in_22_17_i;
reg signed [`InBus]		in_22_18_r;
reg signed [`InBus]		in_22_18_i;
reg signed [`InBus]		in_22_19_r;
reg signed [`InBus]		in_22_19_i;
reg signed [`InBus]		in_22_20_r;
reg signed [`InBus]		in_22_20_i;
reg signed [`InBus]		in_22_21_r;
reg signed [`InBus]		in_22_21_i;
reg signed [`InBus]		in_22_22_r;
reg signed [`InBus]		in_22_22_i;
reg signed [`InBus]		in_22_23_r;
reg signed [`InBus]		in_22_23_i;
reg signed [`InBus]		in_22_24_r;
reg signed [`InBus]		in_22_24_i;
reg signed [`InBus]		in_22_25_r;
reg signed [`InBus]		in_22_25_i;
reg signed [`InBus]		in_22_26_r;
reg signed [`InBus]		in_22_26_i;
reg signed [`InBus]		in_22_27_r;
reg signed [`InBus]		in_22_27_i;
reg signed [`InBus]		in_22_28_r;
reg signed [`InBus]		in_22_28_i;
reg signed [`InBus]		in_22_29_r;
reg signed [`InBus]		in_22_29_i;
reg signed [`InBus]		in_22_30_r;
reg signed [`InBus]		in_22_30_i;
reg signed [`InBus]		in_22_31_r;
reg signed [`InBus]		in_22_31_i;
reg signed [`InBus]		in_22_32_r;
reg signed [`InBus]		in_22_32_i;
reg signed [`InBus]		in_23_1_r;
reg signed [`InBus]		in_23_1_i;
reg signed [`InBus]		in_23_2_r;
reg signed [`InBus]		in_23_2_i;
reg signed [`InBus]		in_23_3_r;
reg signed [`InBus]		in_23_3_i;
reg signed [`InBus]		in_23_4_r;
reg signed [`InBus]		in_23_4_i;
reg signed [`InBus]		in_23_5_r;
reg signed [`InBus]		in_23_5_i;
reg signed [`InBus]		in_23_6_r;
reg signed [`InBus]		in_23_6_i;
reg signed [`InBus]		in_23_7_r;
reg signed [`InBus]		in_23_7_i;
reg signed [`InBus]		in_23_8_r;
reg signed [`InBus]		in_23_8_i;
reg signed [`InBus]		in_23_9_r;
reg signed [`InBus]		in_23_9_i;
reg signed [`InBus]		in_23_10_r;
reg signed [`InBus]		in_23_10_i;
reg signed [`InBus]		in_23_11_r;
reg signed [`InBus]		in_23_11_i;
reg signed [`InBus]		in_23_12_r;
reg signed [`InBus]		in_23_12_i;
reg signed [`InBus]		in_23_13_r;
reg signed [`InBus]		in_23_13_i;
reg signed [`InBus]		in_23_14_r;
reg signed [`InBus]		in_23_14_i;
reg signed [`InBus]		in_23_15_r;
reg signed [`InBus]		in_23_15_i;
reg signed [`InBus]		in_23_16_r;
reg signed [`InBus]		in_23_16_i;
reg signed [`InBus]		in_23_17_r;
reg signed [`InBus]		in_23_17_i;
reg signed [`InBus]		in_23_18_r;
reg signed [`InBus]		in_23_18_i;
reg signed [`InBus]		in_23_19_r;
reg signed [`InBus]		in_23_19_i;
reg signed [`InBus]		in_23_20_r;
reg signed [`InBus]		in_23_20_i;
reg signed [`InBus]		in_23_21_r;
reg signed [`InBus]		in_23_21_i;
reg signed [`InBus]		in_23_22_r;
reg signed [`InBus]		in_23_22_i;
reg signed [`InBus]		in_23_23_r;
reg signed [`InBus]		in_23_23_i;
reg signed [`InBus]		in_23_24_r;
reg signed [`InBus]		in_23_24_i;
reg signed [`InBus]		in_23_25_r;
reg signed [`InBus]		in_23_25_i;
reg signed [`InBus]		in_23_26_r;
reg signed [`InBus]		in_23_26_i;
reg signed [`InBus]		in_23_27_r;
reg signed [`InBus]		in_23_27_i;
reg signed [`InBus]		in_23_28_r;
reg signed [`InBus]		in_23_28_i;
reg signed [`InBus]		in_23_29_r;
reg signed [`InBus]		in_23_29_i;
reg signed [`InBus]		in_23_30_r;
reg signed [`InBus]		in_23_30_i;
reg signed [`InBus]		in_23_31_r;
reg signed [`InBus]		in_23_31_i;
reg signed [`InBus]		in_23_32_r;
reg signed [`InBus]		in_23_32_i;
reg signed [`InBus]		in_24_1_r;
reg signed [`InBus]		in_24_1_i;
reg signed [`InBus]		in_24_2_r;
reg signed [`InBus]		in_24_2_i;
reg signed [`InBus]		in_24_3_r;
reg signed [`InBus]		in_24_3_i;
reg signed [`InBus]		in_24_4_r;
reg signed [`InBus]		in_24_4_i;
reg signed [`InBus]		in_24_5_r;
reg signed [`InBus]		in_24_5_i;
reg signed [`InBus]		in_24_6_r;
reg signed [`InBus]		in_24_6_i;
reg signed [`InBus]		in_24_7_r;
reg signed [`InBus]		in_24_7_i;
reg signed [`InBus]		in_24_8_r;
reg signed [`InBus]		in_24_8_i;
reg signed [`InBus]		in_24_9_r;
reg signed [`InBus]		in_24_9_i;
reg signed [`InBus]		in_24_10_r;
reg signed [`InBus]		in_24_10_i;
reg signed [`InBus]		in_24_11_r;
reg signed [`InBus]		in_24_11_i;
reg signed [`InBus]		in_24_12_r;
reg signed [`InBus]		in_24_12_i;
reg signed [`InBus]		in_24_13_r;
reg signed [`InBus]		in_24_13_i;
reg signed [`InBus]		in_24_14_r;
reg signed [`InBus]		in_24_14_i;
reg signed [`InBus]		in_24_15_r;
reg signed [`InBus]		in_24_15_i;
reg signed [`InBus]		in_24_16_r;
reg signed [`InBus]		in_24_16_i;
reg signed [`InBus]		in_24_17_r;
reg signed [`InBus]		in_24_17_i;
reg signed [`InBus]		in_24_18_r;
reg signed [`InBus]		in_24_18_i;
reg signed [`InBus]		in_24_19_r;
reg signed [`InBus]		in_24_19_i;
reg signed [`InBus]		in_24_20_r;
reg signed [`InBus]		in_24_20_i;
reg signed [`InBus]		in_24_21_r;
reg signed [`InBus]		in_24_21_i;
reg signed [`InBus]		in_24_22_r;
reg signed [`InBus]		in_24_22_i;
reg signed [`InBus]		in_24_23_r;
reg signed [`InBus]		in_24_23_i;
reg signed [`InBus]		in_24_24_r;
reg signed [`InBus]		in_24_24_i;
reg signed [`InBus]		in_24_25_r;
reg signed [`InBus]		in_24_25_i;
reg signed [`InBus]		in_24_26_r;
reg signed [`InBus]		in_24_26_i;
reg signed [`InBus]		in_24_27_r;
reg signed [`InBus]		in_24_27_i;
reg signed [`InBus]		in_24_28_r;
reg signed [`InBus]		in_24_28_i;
reg signed [`InBus]		in_24_29_r;
reg signed [`InBus]		in_24_29_i;
reg signed [`InBus]		in_24_30_r;
reg signed [`InBus]		in_24_30_i;
reg signed [`InBus]		in_24_31_r;
reg signed [`InBus]		in_24_31_i;
reg signed [`InBus]		in_24_32_r;
reg signed [`InBus]		in_24_32_i;
reg signed [`InBus]		in_25_1_r;
reg signed [`InBus]		in_25_1_i;
reg signed [`InBus]		in_25_2_r;
reg signed [`InBus]		in_25_2_i;
reg signed [`InBus]		in_25_3_r;
reg signed [`InBus]		in_25_3_i;
reg signed [`InBus]		in_25_4_r;
reg signed [`InBus]		in_25_4_i;
reg signed [`InBus]		in_25_5_r;
reg signed [`InBus]		in_25_5_i;
reg signed [`InBus]		in_25_6_r;
reg signed [`InBus]		in_25_6_i;
reg signed [`InBus]		in_25_7_r;
reg signed [`InBus]		in_25_7_i;
reg signed [`InBus]		in_25_8_r;
reg signed [`InBus]		in_25_8_i;
reg signed [`InBus]		in_25_9_r;
reg signed [`InBus]		in_25_9_i;
reg signed [`InBus]		in_25_10_r;
reg signed [`InBus]		in_25_10_i;
reg signed [`InBus]		in_25_11_r;
reg signed [`InBus]		in_25_11_i;
reg signed [`InBus]		in_25_12_r;
reg signed [`InBus]		in_25_12_i;
reg signed [`InBus]		in_25_13_r;
reg signed [`InBus]		in_25_13_i;
reg signed [`InBus]		in_25_14_r;
reg signed [`InBus]		in_25_14_i;
reg signed [`InBus]		in_25_15_r;
reg signed [`InBus]		in_25_15_i;
reg signed [`InBus]		in_25_16_r;
reg signed [`InBus]		in_25_16_i;
reg signed [`InBus]		in_25_17_r;
reg signed [`InBus]		in_25_17_i;
reg signed [`InBus]		in_25_18_r;
reg signed [`InBus]		in_25_18_i;
reg signed [`InBus]		in_25_19_r;
reg signed [`InBus]		in_25_19_i;
reg signed [`InBus]		in_25_20_r;
reg signed [`InBus]		in_25_20_i;
reg signed [`InBus]		in_25_21_r;
reg signed [`InBus]		in_25_21_i;
reg signed [`InBus]		in_25_22_r;
reg signed [`InBus]		in_25_22_i;
reg signed [`InBus]		in_25_23_r;
reg signed [`InBus]		in_25_23_i;
reg signed [`InBus]		in_25_24_r;
reg signed [`InBus]		in_25_24_i;
reg signed [`InBus]		in_25_25_r;
reg signed [`InBus]		in_25_25_i;
reg signed [`InBus]		in_25_26_r;
reg signed [`InBus]		in_25_26_i;
reg signed [`InBus]		in_25_27_r;
reg signed [`InBus]		in_25_27_i;
reg signed [`InBus]		in_25_28_r;
reg signed [`InBus]		in_25_28_i;
reg signed [`InBus]		in_25_29_r;
reg signed [`InBus]		in_25_29_i;
reg signed [`InBus]		in_25_30_r;
reg signed [`InBus]		in_25_30_i;
reg signed [`InBus]		in_25_31_r;
reg signed [`InBus]		in_25_31_i;
reg signed [`InBus]		in_25_32_r;
reg signed [`InBus]		in_25_32_i;
reg signed [`InBus]		in_26_1_r;
reg signed [`InBus]		in_26_1_i;
reg signed [`InBus]		in_26_2_r;
reg signed [`InBus]		in_26_2_i;
reg signed [`InBus]		in_26_3_r;
reg signed [`InBus]		in_26_3_i;
reg signed [`InBus]		in_26_4_r;
reg signed [`InBus]		in_26_4_i;
reg signed [`InBus]		in_26_5_r;
reg signed [`InBus]		in_26_5_i;
reg signed [`InBus]		in_26_6_r;
reg signed [`InBus]		in_26_6_i;
reg signed [`InBus]		in_26_7_r;
reg signed [`InBus]		in_26_7_i;
reg signed [`InBus]		in_26_8_r;
reg signed [`InBus]		in_26_8_i;
reg signed [`InBus]		in_26_9_r;
reg signed [`InBus]		in_26_9_i;
reg signed [`InBus]		in_26_10_r;
reg signed [`InBus]		in_26_10_i;
reg signed [`InBus]		in_26_11_r;
reg signed [`InBus]		in_26_11_i;
reg signed [`InBus]		in_26_12_r;
reg signed [`InBus]		in_26_12_i;
reg signed [`InBus]		in_26_13_r;
reg signed [`InBus]		in_26_13_i;
reg signed [`InBus]		in_26_14_r;
reg signed [`InBus]		in_26_14_i;
reg signed [`InBus]		in_26_15_r;
reg signed [`InBus]		in_26_15_i;
reg signed [`InBus]		in_26_16_r;
reg signed [`InBus]		in_26_16_i;
reg signed [`InBus]		in_26_17_r;
reg signed [`InBus]		in_26_17_i;
reg signed [`InBus]		in_26_18_r;
reg signed [`InBus]		in_26_18_i;
reg signed [`InBus]		in_26_19_r;
reg signed [`InBus]		in_26_19_i;
reg signed [`InBus]		in_26_20_r;
reg signed [`InBus]		in_26_20_i;
reg signed [`InBus]		in_26_21_r;
reg signed [`InBus]		in_26_21_i;
reg signed [`InBus]		in_26_22_r;
reg signed [`InBus]		in_26_22_i;
reg signed [`InBus]		in_26_23_r;
reg signed [`InBus]		in_26_23_i;
reg signed [`InBus]		in_26_24_r;
reg signed [`InBus]		in_26_24_i;
reg signed [`InBus]		in_26_25_r;
reg signed [`InBus]		in_26_25_i;
reg signed [`InBus]		in_26_26_r;
reg signed [`InBus]		in_26_26_i;
reg signed [`InBus]		in_26_27_r;
reg signed [`InBus]		in_26_27_i;
reg signed [`InBus]		in_26_28_r;
reg signed [`InBus]		in_26_28_i;
reg signed [`InBus]		in_26_29_r;
reg signed [`InBus]		in_26_29_i;
reg signed [`InBus]		in_26_30_r;
reg signed [`InBus]		in_26_30_i;
reg signed [`InBus]		in_26_31_r;
reg signed [`InBus]		in_26_31_i;
reg signed [`InBus]		in_26_32_r;
reg signed [`InBus]		in_26_32_i;
reg signed [`InBus]		in_27_1_r;
reg signed [`InBus]		in_27_1_i;
reg signed [`InBus]		in_27_2_r;
reg signed [`InBus]		in_27_2_i;
reg signed [`InBus]		in_27_3_r;
reg signed [`InBus]		in_27_3_i;
reg signed [`InBus]		in_27_4_r;
reg signed [`InBus]		in_27_4_i;
reg signed [`InBus]		in_27_5_r;
reg signed [`InBus]		in_27_5_i;
reg signed [`InBus]		in_27_6_r;
reg signed [`InBus]		in_27_6_i;
reg signed [`InBus]		in_27_7_r;
reg signed [`InBus]		in_27_7_i;
reg signed [`InBus]		in_27_8_r;
reg signed [`InBus]		in_27_8_i;
reg signed [`InBus]		in_27_9_r;
reg signed [`InBus]		in_27_9_i;
reg signed [`InBus]		in_27_10_r;
reg signed [`InBus]		in_27_10_i;
reg signed [`InBus]		in_27_11_r;
reg signed [`InBus]		in_27_11_i;
reg signed [`InBus]		in_27_12_r;
reg signed [`InBus]		in_27_12_i;
reg signed [`InBus]		in_27_13_r;
reg signed [`InBus]		in_27_13_i;
reg signed [`InBus]		in_27_14_r;
reg signed [`InBus]		in_27_14_i;
reg signed [`InBus]		in_27_15_r;
reg signed [`InBus]		in_27_15_i;
reg signed [`InBus]		in_27_16_r;
reg signed [`InBus]		in_27_16_i;
reg signed [`InBus]		in_27_17_r;
reg signed [`InBus]		in_27_17_i;
reg signed [`InBus]		in_27_18_r;
reg signed [`InBus]		in_27_18_i;
reg signed [`InBus]		in_27_19_r;
reg signed [`InBus]		in_27_19_i;
reg signed [`InBus]		in_27_20_r;
reg signed [`InBus]		in_27_20_i;
reg signed [`InBus]		in_27_21_r;
reg signed [`InBus]		in_27_21_i;
reg signed [`InBus]		in_27_22_r;
reg signed [`InBus]		in_27_22_i;
reg signed [`InBus]		in_27_23_r;
reg signed [`InBus]		in_27_23_i;
reg signed [`InBus]		in_27_24_r;
reg signed [`InBus]		in_27_24_i;
reg signed [`InBus]		in_27_25_r;
reg signed [`InBus]		in_27_25_i;
reg signed [`InBus]		in_27_26_r;
reg signed [`InBus]		in_27_26_i;
reg signed [`InBus]		in_27_27_r;
reg signed [`InBus]		in_27_27_i;
reg signed [`InBus]		in_27_28_r;
reg signed [`InBus]		in_27_28_i;
reg signed [`InBus]		in_27_29_r;
reg signed [`InBus]		in_27_29_i;
reg signed [`InBus]		in_27_30_r;
reg signed [`InBus]		in_27_30_i;
reg signed [`InBus]		in_27_31_r;
reg signed [`InBus]		in_27_31_i;
reg signed [`InBus]		in_27_32_r;
reg signed [`InBus]		in_27_32_i;
reg signed [`InBus]		in_28_1_r;
reg signed [`InBus]		in_28_1_i;
reg signed [`InBus]		in_28_2_r;
reg signed [`InBus]		in_28_2_i;
reg signed [`InBus]		in_28_3_r;
reg signed [`InBus]		in_28_3_i;
reg signed [`InBus]		in_28_4_r;
reg signed [`InBus]		in_28_4_i;
reg signed [`InBus]		in_28_5_r;
reg signed [`InBus]		in_28_5_i;
reg signed [`InBus]		in_28_6_r;
reg signed [`InBus]		in_28_6_i;
reg signed [`InBus]		in_28_7_r;
reg signed [`InBus]		in_28_7_i;
reg signed [`InBus]		in_28_8_r;
reg signed [`InBus]		in_28_8_i;
reg signed [`InBus]		in_28_9_r;
reg signed [`InBus]		in_28_9_i;
reg signed [`InBus]		in_28_10_r;
reg signed [`InBus]		in_28_10_i;
reg signed [`InBus]		in_28_11_r;
reg signed [`InBus]		in_28_11_i;
reg signed [`InBus]		in_28_12_r;
reg signed [`InBus]		in_28_12_i;
reg signed [`InBus]		in_28_13_r;
reg signed [`InBus]		in_28_13_i;
reg signed [`InBus]		in_28_14_r;
reg signed [`InBus]		in_28_14_i;
reg signed [`InBus]		in_28_15_r;
reg signed [`InBus]		in_28_15_i;
reg signed [`InBus]		in_28_16_r;
reg signed [`InBus]		in_28_16_i;
reg signed [`InBus]		in_28_17_r;
reg signed [`InBus]		in_28_17_i;
reg signed [`InBus]		in_28_18_r;
reg signed [`InBus]		in_28_18_i;
reg signed [`InBus]		in_28_19_r;
reg signed [`InBus]		in_28_19_i;
reg signed [`InBus]		in_28_20_r;
reg signed [`InBus]		in_28_20_i;
reg signed [`InBus]		in_28_21_r;
reg signed [`InBus]		in_28_21_i;
reg signed [`InBus]		in_28_22_r;
reg signed [`InBus]		in_28_22_i;
reg signed [`InBus]		in_28_23_r;
reg signed [`InBus]		in_28_23_i;
reg signed [`InBus]		in_28_24_r;
reg signed [`InBus]		in_28_24_i;
reg signed [`InBus]		in_28_25_r;
reg signed [`InBus]		in_28_25_i;
reg signed [`InBus]		in_28_26_r;
reg signed [`InBus]		in_28_26_i;
reg signed [`InBus]		in_28_27_r;
reg signed [`InBus]		in_28_27_i;
reg signed [`InBus]		in_28_28_r;
reg signed [`InBus]		in_28_28_i;
reg signed [`InBus]		in_28_29_r;
reg signed [`InBus]		in_28_29_i;
reg signed [`InBus]		in_28_30_r;
reg signed [`InBus]		in_28_30_i;
reg signed [`InBus]		in_28_31_r;
reg signed [`InBus]		in_28_31_i;
reg signed [`InBus]		in_28_32_r;
reg signed [`InBus]		in_28_32_i;
reg signed [`InBus]		in_29_1_r;
reg signed [`InBus]		in_29_1_i;
reg signed [`InBus]		in_29_2_r;
reg signed [`InBus]		in_29_2_i;
reg signed [`InBus]		in_29_3_r;
reg signed [`InBus]		in_29_3_i;
reg signed [`InBus]		in_29_4_r;
reg signed [`InBus]		in_29_4_i;
reg signed [`InBus]		in_29_5_r;
reg signed [`InBus]		in_29_5_i;
reg signed [`InBus]		in_29_6_r;
reg signed [`InBus]		in_29_6_i;
reg signed [`InBus]		in_29_7_r;
reg signed [`InBus]		in_29_7_i;
reg signed [`InBus]		in_29_8_r;
reg signed [`InBus]		in_29_8_i;
reg signed [`InBus]		in_29_9_r;
reg signed [`InBus]		in_29_9_i;
reg signed [`InBus]		in_29_10_r;
reg signed [`InBus]		in_29_10_i;
reg signed [`InBus]		in_29_11_r;
reg signed [`InBus]		in_29_11_i;
reg signed [`InBus]		in_29_12_r;
reg signed [`InBus]		in_29_12_i;
reg signed [`InBus]		in_29_13_r;
reg signed [`InBus]		in_29_13_i;
reg signed [`InBus]		in_29_14_r;
reg signed [`InBus]		in_29_14_i;
reg signed [`InBus]		in_29_15_r;
reg signed [`InBus]		in_29_15_i;
reg signed [`InBus]		in_29_16_r;
reg signed [`InBus]		in_29_16_i;
reg signed [`InBus]		in_29_17_r;
reg signed [`InBus]		in_29_17_i;
reg signed [`InBus]		in_29_18_r;
reg signed [`InBus]		in_29_18_i;
reg signed [`InBus]		in_29_19_r;
reg signed [`InBus]		in_29_19_i;
reg signed [`InBus]		in_29_20_r;
reg signed [`InBus]		in_29_20_i;
reg signed [`InBus]		in_29_21_r;
reg signed [`InBus]		in_29_21_i;
reg signed [`InBus]		in_29_22_r;
reg signed [`InBus]		in_29_22_i;
reg signed [`InBus]		in_29_23_r;
reg signed [`InBus]		in_29_23_i;
reg signed [`InBus]		in_29_24_r;
reg signed [`InBus]		in_29_24_i;
reg signed [`InBus]		in_29_25_r;
reg signed [`InBus]		in_29_25_i;
reg signed [`InBus]		in_29_26_r;
reg signed [`InBus]		in_29_26_i;
reg signed [`InBus]		in_29_27_r;
reg signed [`InBus]		in_29_27_i;
reg signed [`InBus]		in_29_28_r;
reg signed [`InBus]		in_29_28_i;
reg signed [`InBus]		in_29_29_r;
reg signed [`InBus]		in_29_29_i;
reg signed [`InBus]		in_29_30_r;
reg signed [`InBus]		in_29_30_i;
reg signed [`InBus]		in_29_31_r;
reg signed [`InBus]		in_29_31_i;
reg signed [`InBus]		in_29_32_r;
reg signed [`InBus]		in_29_32_i;
reg signed [`InBus]		in_30_1_r;
reg signed [`InBus]		in_30_1_i;
reg signed [`InBus]		in_30_2_r;
reg signed [`InBus]		in_30_2_i;
reg signed [`InBus]		in_30_3_r;
reg signed [`InBus]		in_30_3_i;
reg signed [`InBus]		in_30_4_r;
reg signed [`InBus]		in_30_4_i;
reg signed [`InBus]		in_30_5_r;
reg signed [`InBus]		in_30_5_i;
reg signed [`InBus]		in_30_6_r;
reg signed [`InBus]		in_30_6_i;
reg signed [`InBus]		in_30_7_r;
reg signed [`InBus]		in_30_7_i;
reg signed [`InBus]		in_30_8_r;
reg signed [`InBus]		in_30_8_i;
reg signed [`InBus]		in_30_9_r;
reg signed [`InBus]		in_30_9_i;
reg signed [`InBus]		in_30_10_r;
reg signed [`InBus]		in_30_10_i;
reg signed [`InBus]		in_30_11_r;
reg signed [`InBus]		in_30_11_i;
reg signed [`InBus]		in_30_12_r;
reg signed [`InBus]		in_30_12_i;
reg signed [`InBus]		in_30_13_r;
reg signed [`InBus]		in_30_13_i;
reg signed [`InBus]		in_30_14_r;
reg signed [`InBus]		in_30_14_i;
reg signed [`InBus]		in_30_15_r;
reg signed [`InBus]		in_30_15_i;
reg signed [`InBus]		in_30_16_r;
reg signed [`InBus]		in_30_16_i;
reg signed [`InBus]		in_30_17_r;
reg signed [`InBus]		in_30_17_i;
reg signed [`InBus]		in_30_18_r;
reg signed [`InBus]		in_30_18_i;
reg signed [`InBus]		in_30_19_r;
reg signed [`InBus]		in_30_19_i;
reg signed [`InBus]		in_30_20_r;
reg signed [`InBus]		in_30_20_i;
reg signed [`InBus]		in_30_21_r;
reg signed [`InBus]		in_30_21_i;
reg signed [`InBus]		in_30_22_r;
reg signed [`InBus]		in_30_22_i;
reg signed [`InBus]		in_30_23_r;
reg signed [`InBus]		in_30_23_i;
reg signed [`InBus]		in_30_24_r;
reg signed [`InBus]		in_30_24_i;
reg signed [`InBus]		in_30_25_r;
reg signed [`InBus]		in_30_25_i;
reg signed [`InBus]		in_30_26_r;
reg signed [`InBus]		in_30_26_i;
reg signed [`InBus]		in_30_27_r;
reg signed [`InBus]		in_30_27_i;
reg signed [`InBus]		in_30_28_r;
reg signed [`InBus]		in_30_28_i;
reg signed [`InBus]		in_30_29_r;
reg signed [`InBus]		in_30_29_i;
reg signed [`InBus]		in_30_30_r;
reg signed [`InBus]		in_30_30_i;
reg signed [`InBus]		in_30_31_r;
reg signed [`InBus]		in_30_31_i;
reg signed [`InBus]		in_30_32_r;
reg signed [`InBus]		in_30_32_i;
reg signed [`InBus]		in_31_1_r;
reg signed [`InBus]		in_31_1_i;
reg signed [`InBus]		in_31_2_r;
reg signed [`InBus]		in_31_2_i;
reg signed [`InBus]		in_31_3_r;
reg signed [`InBus]		in_31_3_i;
reg signed [`InBus]		in_31_4_r;
reg signed [`InBus]		in_31_4_i;
reg signed [`InBus]		in_31_5_r;
reg signed [`InBus]		in_31_5_i;
reg signed [`InBus]		in_31_6_r;
reg signed [`InBus]		in_31_6_i;
reg signed [`InBus]		in_31_7_r;
reg signed [`InBus]		in_31_7_i;
reg signed [`InBus]		in_31_8_r;
reg signed [`InBus]		in_31_8_i;
reg signed [`InBus]		in_31_9_r;
reg signed [`InBus]		in_31_9_i;
reg signed [`InBus]		in_31_10_r;
reg signed [`InBus]		in_31_10_i;
reg signed [`InBus]		in_31_11_r;
reg signed [`InBus]		in_31_11_i;
reg signed [`InBus]		in_31_12_r;
reg signed [`InBus]		in_31_12_i;
reg signed [`InBus]		in_31_13_r;
reg signed [`InBus]		in_31_13_i;
reg signed [`InBus]		in_31_14_r;
reg signed [`InBus]		in_31_14_i;
reg signed [`InBus]		in_31_15_r;
reg signed [`InBus]		in_31_15_i;
reg signed [`InBus]		in_31_16_r;
reg signed [`InBus]		in_31_16_i;
reg signed [`InBus]		in_31_17_r;
reg signed [`InBus]		in_31_17_i;
reg signed [`InBus]		in_31_18_r;
reg signed [`InBus]		in_31_18_i;
reg signed [`InBus]		in_31_19_r;
reg signed [`InBus]		in_31_19_i;
reg signed [`InBus]		in_31_20_r;
reg signed [`InBus]		in_31_20_i;
reg signed [`InBus]		in_31_21_r;
reg signed [`InBus]		in_31_21_i;
reg signed [`InBus]		in_31_22_r;
reg signed [`InBus]		in_31_22_i;
reg signed [`InBus]		in_31_23_r;
reg signed [`InBus]		in_31_23_i;
reg signed [`InBus]		in_31_24_r;
reg signed [`InBus]		in_31_24_i;
reg signed [`InBus]		in_31_25_r;
reg signed [`InBus]		in_31_25_i;
reg signed [`InBus]		in_31_26_r;
reg signed [`InBus]		in_31_26_i;
reg signed [`InBus]		in_31_27_r;
reg signed [`InBus]		in_31_27_i;
reg signed [`InBus]		in_31_28_r;
reg signed [`InBus]		in_31_28_i;
reg signed [`InBus]		in_31_29_r;
reg signed [`InBus]		in_31_29_i;
reg signed [`InBus]		in_31_30_r;
reg signed [`InBus]		in_31_30_i;
reg signed [`InBus]		in_31_31_r;
reg signed [`InBus]		in_31_31_i;
reg signed [`InBus]		in_31_32_r;
reg signed [`InBus]		in_31_32_i;
reg signed [`InBus]		in_32_1_r;
reg signed [`InBus]		in_32_1_i;
reg signed [`InBus]		in_32_2_r;
reg signed [`InBus]		in_32_2_i;
reg signed [`InBus]		in_32_3_r;
reg signed [`InBus]		in_32_3_i;
reg signed [`InBus]		in_32_4_r;
reg signed [`InBus]		in_32_4_i;
reg signed [`InBus]		in_32_5_r;
reg signed [`InBus]		in_32_5_i;
reg signed [`InBus]		in_32_6_r;
reg signed [`InBus]		in_32_6_i;
reg signed [`InBus]		in_32_7_r;
reg signed [`InBus]		in_32_7_i;
reg signed [`InBus]		in_32_8_r;
reg signed [`InBus]		in_32_8_i;
reg signed [`InBus]		in_32_9_r;
reg signed [`InBus]		in_32_9_i;
reg signed [`InBus]		in_32_10_r;
reg signed [`InBus]		in_32_10_i;
reg signed [`InBus]		in_32_11_r;
reg signed [`InBus]		in_32_11_i;
reg signed [`InBus]		in_32_12_r;
reg signed [`InBus]		in_32_12_i;
reg signed [`InBus]		in_32_13_r;
reg signed [`InBus]		in_32_13_i;
reg signed [`InBus]		in_32_14_r;
reg signed [`InBus]		in_32_14_i;
reg signed [`InBus]		in_32_15_r;
reg signed [`InBus]		in_32_15_i;
reg signed [`InBus]		in_32_16_r;
reg signed [`InBus]		in_32_16_i;
reg signed [`InBus]		in_32_17_r;
reg signed [`InBus]		in_32_17_i;
reg signed [`InBus]		in_32_18_r;
reg signed [`InBus]		in_32_18_i;
reg signed [`InBus]		in_32_19_r;
reg signed [`InBus]		in_32_19_i;
reg signed [`InBus]		in_32_20_r;
reg signed [`InBus]		in_32_20_i;
reg signed [`InBus]		in_32_21_r;
reg signed [`InBus]		in_32_21_i;
reg signed [`InBus]		in_32_22_r;
reg signed [`InBus]		in_32_22_i;
reg signed [`InBus]		in_32_23_r;
reg signed [`InBus]		in_32_23_i;
reg signed [`InBus]		in_32_24_r;
reg signed [`InBus]		in_32_24_i;
reg signed [`InBus]		in_32_25_r;
reg signed [`InBus]		in_32_25_i;
reg signed [`InBus]		in_32_26_r;
reg signed [`InBus]		in_32_26_i;
reg signed [`InBus]		in_32_27_r;
reg signed [`InBus]		in_32_27_i;
reg signed [`InBus]		in_32_28_r;
reg signed [`InBus]		in_32_28_i;
reg signed [`InBus]		in_32_29_r;
reg signed [`InBus]		in_32_29_i;
reg signed [`InBus]		in_32_30_r;
reg signed [`InBus]		in_32_30_i;
reg signed [`InBus]		in_32_31_r;
reg signed [`InBus]		in_32_31_i;
reg signed [`InBus]		in_32_32_r;
reg signed [`InBus]		in_32_32_i;

wire signed [`OutBus]		out_1_1_r;
wire signed [`OutBus]		out_1_1_i;
wire signed [`OutBus]		out_1_2_r;
wire signed [`OutBus]		out_1_2_i;
wire signed [`OutBus]		out_1_3_r;
wire signed [`OutBus]		out_1_3_i;
wire signed [`OutBus]		out_1_4_r;
wire signed [`OutBus]		out_1_4_i;
wire signed [`OutBus]		out_1_5_r;
wire signed [`OutBus]		out_1_5_i;
wire signed [`OutBus]		out_1_6_r;
wire signed [`OutBus]		out_1_6_i;
wire signed [`OutBus]		out_1_7_r;
wire signed [`OutBus]		out_1_7_i;
wire signed [`OutBus]		out_1_8_r;
wire signed [`OutBus]		out_1_8_i;
wire signed [`OutBus]		out_1_9_r;
wire signed [`OutBus]		out_1_9_i;
wire signed [`OutBus]		out_1_10_r;
wire signed [`OutBus]		out_1_10_i;
wire signed [`OutBus]		out_1_11_r;
wire signed [`OutBus]		out_1_11_i;
wire signed [`OutBus]		out_1_12_r;
wire signed [`OutBus]		out_1_12_i;
wire signed [`OutBus]		out_1_13_r;
wire signed [`OutBus]		out_1_13_i;
wire signed [`OutBus]		out_1_14_r;
wire signed [`OutBus]		out_1_14_i;
wire signed [`OutBus]		out_1_15_r;
wire signed [`OutBus]		out_1_15_i;
wire signed [`OutBus]		out_1_16_r;
wire signed [`OutBus]		out_1_16_i;
wire signed [`OutBus]		out_1_17_r;
wire signed [`OutBus]		out_1_17_i;
wire signed [`OutBus]		out_1_18_r;
wire signed [`OutBus]		out_1_18_i;
wire signed [`OutBus]		out_1_19_r;
wire signed [`OutBus]		out_1_19_i;
wire signed [`OutBus]		out_1_20_r;
wire signed [`OutBus]		out_1_20_i;
wire signed [`OutBus]		out_1_21_r;
wire signed [`OutBus]		out_1_21_i;
wire signed [`OutBus]		out_1_22_r;
wire signed [`OutBus]		out_1_22_i;
wire signed [`OutBus]		out_1_23_r;
wire signed [`OutBus]		out_1_23_i;
wire signed [`OutBus]		out_1_24_r;
wire signed [`OutBus]		out_1_24_i;
wire signed [`OutBus]		out_1_25_r;
wire signed [`OutBus]		out_1_25_i;
wire signed [`OutBus]		out_1_26_r;
wire signed [`OutBus]		out_1_26_i;
wire signed [`OutBus]		out_1_27_r;
wire signed [`OutBus]		out_1_27_i;
wire signed [`OutBus]		out_1_28_r;
wire signed [`OutBus]		out_1_28_i;
wire signed [`OutBus]		out_1_29_r;
wire signed [`OutBus]		out_1_29_i;
wire signed [`OutBus]		out_1_30_r;
wire signed [`OutBus]		out_1_30_i;
wire signed [`OutBus]		out_1_31_r;
wire signed [`OutBus]		out_1_31_i;
wire signed [`OutBus]		out_1_32_r;
wire signed [`OutBus]		out_1_32_i;
wire signed [`OutBus]		out_2_1_r;
wire signed [`OutBus]		out_2_1_i;
wire signed [`OutBus]		out_2_2_r;
wire signed [`OutBus]		out_2_2_i;
wire signed [`OutBus]		out_2_3_r;
wire signed [`OutBus]		out_2_3_i;
wire signed [`OutBus]		out_2_4_r;
wire signed [`OutBus]		out_2_4_i;
wire signed [`OutBus]		out_2_5_r;
wire signed [`OutBus]		out_2_5_i;
wire signed [`OutBus]		out_2_6_r;
wire signed [`OutBus]		out_2_6_i;
wire signed [`OutBus]		out_2_7_r;
wire signed [`OutBus]		out_2_7_i;
wire signed [`OutBus]		out_2_8_r;
wire signed [`OutBus]		out_2_8_i;
wire signed [`OutBus]		out_2_9_r;
wire signed [`OutBus]		out_2_9_i;
wire signed [`OutBus]		out_2_10_r;
wire signed [`OutBus]		out_2_10_i;
wire signed [`OutBus]		out_2_11_r;
wire signed [`OutBus]		out_2_11_i;
wire signed [`OutBus]		out_2_12_r;
wire signed [`OutBus]		out_2_12_i;
wire signed [`OutBus]		out_2_13_r;
wire signed [`OutBus]		out_2_13_i;
wire signed [`OutBus]		out_2_14_r;
wire signed [`OutBus]		out_2_14_i;
wire signed [`OutBus]		out_2_15_r;
wire signed [`OutBus]		out_2_15_i;
wire signed [`OutBus]		out_2_16_r;
wire signed [`OutBus]		out_2_16_i;
wire signed [`OutBus]		out_2_17_r;
wire signed [`OutBus]		out_2_17_i;
wire signed [`OutBus]		out_2_18_r;
wire signed [`OutBus]		out_2_18_i;
wire signed [`OutBus]		out_2_19_r;
wire signed [`OutBus]		out_2_19_i;
wire signed [`OutBus]		out_2_20_r;
wire signed [`OutBus]		out_2_20_i;
wire signed [`OutBus]		out_2_21_r;
wire signed [`OutBus]		out_2_21_i;
wire signed [`OutBus]		out_2_22_r;
wire signed [`OutBus]		out_2_22_i;
wire signed [`OutBus]		out_2_23_r;
wire signed [`OutBus]		out_2_23_i;
wire signed [`OutBus]		out_2_24_r;
wire signed [`OutBus]		out_2_24_i;
wire signed [`OutBus]		out_2_25_r;
wire signed [`OutBus]		out_2_25_i;
wire signed [`OutBus]		out_2_26_r;
wire signed [`OutBus]		out_2_26_i;
wire signed [`OutBus]		out_2_27_r;
wire signed [`OutBus]		out_2_27_i;
wire signed [`OutBus]		out_2_28_r;
wire signed [`OutBus]		out_2_28_i;
wire signed [`OutBus]		out_2_29_r;
wire signed [`OutBus]		out_2_29_i;
wire signed [`OutBus]		out_2_30_r;
wire signed [`OutBus]		out_2_30_i;
wire signed [`OutBus]		out_2_31_r;
wire signed [`OutBus]		out_2_31_i;
wire signed [`OutBus]		out_2_32_r;
wire signed [`OutBus]		out_2_32_i;
wire signed [`OutBus]		out_3_1_r;
wire signed [`OutBus]		out_3_1_i;
wire signed [`OutBus]		out_3_2_r;
wire signed [`OutBus]		out_3_2_i;
wire signed [`OutBus]		out_3_3_r;
wire signed [`OutBus]		out_3_3_i;
wire signed [`OutBus]		out_3_4_r;
wire signed [`OutBus]		out_3_4_i;
wire signed [`OutBus]		out_3_5_r;
wire signed [`OutBus]		out_3_5_i;
wire signed [`OutBus]		out_3_6_r;
wire signed [`OutBus]		out_3_6_i;
wire signed [`OutBus]		out_3_7_r;
wire signed [`OutBus]		out_3_7_i;
wire signed [`OutBus]		out_3_8_r;
wire signed [`OutBus]		out_3_8_i;
wire signed [`OutBus]		out_3_9_r;
wire signed [`OutBus]		out_3_9_i;
wire signed [`OutBus]		out_3_10_r;
wire signed [`OutBus]		out_3_10_i;
wire signed [`OutBus]		out_3_11_r;
wire signed [`OutBus]		out_3_11_i;
wire signed [`OutBus]		out_3_12_r;
wire signed [`OutBus]		out_3_12_i;
wire signed [`OutBus]		out_3_13_r;
wire signed [`OutBus]		out_3_13_i;
wire signed [`OutBus]		out_3_14_r;
wire signed [`OutBus]		out_3_14_i;
wire signed [`OutBus]		out_3_15_r;
wire signed [`OutBus]		out_3_15_i;
wire signed [`OutBus]		out_3_16_r;
wire signed [`OutBus]		out_3_16_i;
wire signed [`OutBus]		out_3_17_r;
wire signed [`OutBus]		out_3_17_i;
wire signed [`OutBus]		out_3_18_r;
wire signed [`OutBus]		out_3_18_i;
wire signed [`OutBus]		out_3_19_r;
wire signed [`OutBus]		out_3_19_i;
wire signed [`OutBus]		out_3_20_r;
wire signed [`OutBus]		out_3_20_i;
wire signed [`OutBus]		out_3_21_r;
wire signed [`OutBus]		out_3_21_i;
wire signed [`OutBus]		out_3_22_r;
wire signed [`OutBus]		out_3_22_i;
wire signed [`OutBus]		out_3_23_r;
wire signed [`OutBus]		out_3_23_i;
wire signed [`OutBus]		out_3_24_r;
wire signed [`OutBus]		out_3_24_i;
wire signed [`OutBus]		out_3_25_r;
wire signed [`OutBus]		out_3_25_i;
wire signed [`OutBus]		out_3_26_r;
wire signed [`OutBus]		out_3_26_i;
wire signed [`OutBus]		out_3_27_r;
wire signed [`OutBus]		out_3_27_i;
wire signed [`OutBus]		out_3_28_r;
wire signed [`OutBus]		out_3_28_i;
wire signed [`OutBus]		out_3_29_r;
wire signed [`OutBus]		out_3_29_i;
wire signed [`OutBus]		out_3_30_r;
wire signed [`OutBus]		out_3_30_i;
wire signed [`OutBus]		out_3_31_r;
wire signed [`OutBus]		out_3_31_i;
wire signed [`OutBus]		out_3_32_r;
wire signed [`OutBus]		out_3_32_i;
wire signed [`OutBus]		out_4_1_r;
wire signed [`OutBus]		out_4_1_i;
wire signed [`OutBus]		out_4_2_r;
wire signed [`OutBus]		out_4_2_i;
wire signed [`OutBus]		out_4_3_r;
wire signed [`OutBus]		out_4_3_i;
wire signed [`OutBus]		out_4_4_r;
wire signed [`OutBus]		out_4_4_i;
wire signed [`OutBus]		out_4_5_r;
wire signed [`OutBus]		out_4_5_i;
wire signed [`OutBus]		out_4_6_r;
wire signed [`OutBus]		out_4_6_i;
wire signed [`OutBus]		out_4_7_r;
wire signed [`OutBus]		out_4_7_i;
wire signed [`OutBus]		out_4_8_r;
wire signed [`OutBus]		out_4_8_i;
wire signed [`OutBus]		out_4_9_r;
wire signed [`OutBus]		out_4_9_i;
wire signed [`OutBus]		out_4_10_r;
wire signed [`OutBus]		out_4_10_i;
wire signed [`OutBus]		out_4_11_r;
wire signed [`OutBus]		out_4_11_i;
wire signed [`OutBus]		out_4_12_r;
wire signed [`OutBus]		out_4_12_i;
wire signed [`OutBus]		out_4_13_r;
wire signed [`OutBus]		out_4_13_i;
wire signed [`OutBus]		out_4_14_r;
wire signed [`OutBus]		out_4_14_i;
wire signed [`OutBus]		out_4_15_r;
wire signed [`OutBus]		out_4_15_i;
wire signed [`OutBus]		out_4_16_r;
wire signed [`OutBus]		out_4_16_i;
wire signed [`OutBus]		out_4_17_r;
wire signed [`OutBus]		out_4_17_i;
wire signed [`OutBus]		out_4_18_r;
wire signed [`OutBus]		out_4_18_i;
wire signed [`OutBus]		out_4_19_r;
wire signed [`OutBus]		out_4_19_i;
wire signed [`OutBus]		out_4_20_r;
wire signed [`OutBus]		out_4_20_i;
wire signed [`OutBus]		out_4_21_r;
wire signed [`OutBus]		out_4_21_i;
wire signed [`OutBus]		out_4_22_r;
wire signed [`OutBus]		out_4_22_i;
wire signed [`OutBus]		out_4_23_r;
wire signed [`OutBus]		out_4_23_i;
wire signed [`OutBus]		out_4_24_r;
wire signed [`OutBus]		out_4_24_i;
wire signed [`OutBus]		out_4_25_r;
wire signed [`OutBus]		out_4_25_i;
wire signed [`OutBus]		out_4_26_r;
wire signed [`OutBus]		out_4_26_i;
wire signed [`OutBus]		out_4_27_r;
wire signed [`OutBus]		out_4_27_i;
wire signed [`OutBus]		out_4_28_r;
wire signed [`OutBus]		out_4_28_i;
wire signed [`OutBus]		out_4_29_r;
wire signed [`OutBus]		out_4_29_i;
wire signed [`OutBus]		out_4_30_r;
wire signed [`OutBus]		out_4_30_i;
wire signed [`OutBus]		out_4_31_r;
wire signed [`OutBus]		out_4_31_i;
wire signed [`OutBus]		out_4_32_r;
wire signed [`OutBus]		out_4_32_i;
wire signed [`OutBus]		out_5_1_r;
wire signed [`OutBus]		out_5_1_i;
wire signed [`OutBus]		out_5_2_r;
wire signed [`OutBus]		out_5_2_i;
wire signed [`OutBus]		out_5_3_r;
wire signed [`OutBus]		out_5_3_i;
wire signed [`OutBus]		out_5_4_r;
wire signed [`OutBus]		out_5_4_i;
wire signed [`OutBus]		out_5_5_r;
wire signed [`OutBus]		out_5_5_i;
wire signed [`OutBus]		out_5_6_r;
wire signed [`OutBus]		out_5_6_i;
wire signed [`OutBus]		out_5_7_r;
wire signed [`OutBus]		out_5_7_i;
wire signed [`OutBus]		out_5_8_r;
wire signed [`OutBus]		out_5_8_i;
wire signed [`OutBus]		out_5_9_r;
wire signed [`OutBus]		out_5_9_i;
wire signed [`OutBus]		out_5_10_r;
wire signed [`OutBus]		out_5_10_i;
wire signed [`OutBus]		out_5_11_r;
wire signed [`OutBus]		out_5_11_i;
wire signed [`OutBus]		out_5_12_r;
wire signed [`OutBus]		out_5_12_i;
wire signed [`OutBus]		out_5_13_r;
wire signed [`OutBus]		out_5_13_i;
wire signed [`OutBus]		out_5_14_r;
wire signed [`OutBus]		out_5_14_i;
wire signed [`OutBus]		out_5_15_r;
wire signed [`OutBus]		out_5_15_i;
wire signed [`OutBus]		out_5_16_r;
wire signed [`OutBus]		out_5_16_i;
wire signed [`OutBus]		out_5_17_r;
wire signed [`OutBus]		out_5_17_i;
wire signed [`OutBus]		out_5_18_r;
wire signed [`OutBus]		out_5_18_i;
wire signed [`OutBus]		out_5_19_r;
wire signed [`OutBus]		out_5_19_i;
wire signed [`OutBus]		out_5_20_r;
wire signed [`OutBus]		out_5_20_i;
wire signed [`OutBus]		out_5_21_r;
wire signed [`OutBus]		out_5_21_i;
wire signed [`OutBus]		out_5_22_r;
wire signed [`OutBus]		out_5_22_i;
wire signed [`OutBus]		out_5_23_r;
wire signed [`OutBus]		out_5_23_i;
wire signed [`OutBus]		out_5_24_r;
wire signed [`OutBus]		out_5_24_i;
wire signed [`OutBus]		out_5_25_r;
wire signed [`OutBus]		out_5_25_i;
wire signed [`OutBus]		out_5_26_r;
wire signed [`OutBus]		out_5_26_i;
wire signed [`OutBus]		out_5_27_r;
wire signed [`OutBus]		out_5_27_i;
wire signed [`OutBus]		out_5_28_r;
wire signed [`OutBus]		out_5_28_i;
wire signed [`OutBus]		out_5_29_r;
wire signed [`OutBus]		out_5_29_i;
wire signed [`OutBus]		out_5_30_r;
wire signed [`OutBus]		out_5_30_i;
wire signed [`OutBus]		out_5_31_r;
wire signed [`OutBus]		out_5_31_i;
wire signed [`OutBus]		out_5_32_r;
wire signed [`OutBus]		out_5_32_i;
wire signed [`OutBus]		out_6_1_r;
wire signed [`OutBus]		out_6_1_i;
wire signed [`OutBus]		out_6_2_r;
wire signed [`OutBus]		out_6_2_i;
wire signed [`OutBus]		out_6_3_r;
wire signed [`OutBus]		out_6_3_i;
wire signed [`OutBus]		out_6_4_r;
wire signed [`OutBus]		out_6_4_i;
wire signed [`OutBus]		out_6_5_r;
wire signed [`OutBus]		out_6_5_i;
wire signed [`OutBus]		out_6_6_r;
wire signed [`OutBus]		out_6_6_i;
wire signed [`OutBus]		out_6_7_r;
wire signed [`OutBus]		out_6_7_i;
wire signed [`OutBus]		out_6_8_r;
wire signed [`OutBus]		out_6_8_i;
wire signed [`OutBus]		out_6_9_r;
wire signed [`OutBus]		out_6_9_i;
wire signed [`OutBus]		out_6_10_r;
wire signed [`OutBus]		out_6_10_i;
wire signed [`OutBus]		out_6_11_r;
wire signed [`OutBus]		out_6_11_i;
wire signed [`OutBus]		out_6_12_r;
wire signed [`OutBus]		out_6_12_i;
wire signed [`OutBus]		out_6_13_r;
wire signed [`OutBus]		out_6_13_i;
wire signed [`OutBus]		out_6_14_r;
wire signed [`OutBus]		out_6_14_i;
wire signed [`OutBus]		out_6_15_r;
wire signed [`OutBus]		out_6_15_i;
wire signed [`OutBus]		out_6_16_r;
wire signed [`OutBus]		out_6_16_i;
wire signed [`OutBus]		out_6_17_r;
wire signed [`OutBus]		out_6_17_i;
wire signed [`OutBus]		out_6_18_r;
wire signed [`OutBus]		out_6_18_i;
wire signed [`OutBus]		out_6_19_r;
wire signed [`OutBus]		out_6_19_i;
wire signed [`OutBus]		out_6_20_r;
wire signed [`OutBus]		out_6_20_i;
wire signed [`OutBus]		out_6_21_r;
wire signed [`OutBus]		out_6_21_i;
wire signed [`OutBus]		out_6_22_r;
wire signed [`OutBus]		out_6_22_i;
wire signed [`OutBus]		out_6_23_r;
wire signed [`OutBus]		out_6_23_i;
wire signed [`OutBus]		out_6_24_r;
wire signed [`OutBus]		out_6_24_i;
wire signed [`OutBus]		out_6_25_r;
wire signed [`OutBus]		out_6_25_i;
wire signed [`OutBus]		out_6_26_r;
wire signed [`OutBus]		out_6_26_i;
wire signed [`OutBus]		out_6_27_r;
wire signed [`OutBus]		out_6_27_i;
wire signed [`OutBus]		out_6_28_r;
wire signed [`OutBus]		out_6_28_i;
wire signed [`OutBus]		out_6_29_r;
wire signed [`OutBus]		out_6_29_i;
wire signed [`OutBus]		out_6_30_r;
wire signed [`OutBus]		out_6_30_i;
wire signed [`OutBus]		out_6_31_r;
wire signed [`OutBus]		out_6_31_i;
wire signed [`OutBus]		out_6_32_r;
wire signed [`OutBus]		out_6_32_i;
wire signed [`OutBus]		out_7_1_r;
wire signed [`OutBus]		out_7_1_i;
wire signed [`OutBus]		out_7_2_r;
wire signed [`OutBus]		out_7_2_i;
wire signed [`OutBus]		out_7_3_r;
wire signed [`OutBus]		out_7_3_i;
wire signed [`OutBus]		out_7_4_r;
wire signed [`OutBus]		out_7_4_i;
wire signed [`OutBus]		out_7_5_r;
wire signed [`OutBus]		out_7_5_i;
wire signed [`OutBus]		out_7_6_r;
wire signed [`OutBus]		out_7_6_i;
wire signed [`OutBus]		out_7_7_r;
wire signed [`OutBus]		out_7_7_i;
wire signed [`OutBus]		out_7_8_r;
wire signed [`OutBus]		out_7_8_i;
wire signed [`OutBus]		out_7_9_r;
wire signed [`OutBus]		out_7_9_i;
wire signed [`OutBus]		out_7_10_r;
wire signed [`OutBus]		out_7_10_i;
wire signed [`OutBus]		out_7_11_r;
wire signed [`OutBus]		out_7_11_i;
wire signed [`OutBus]		out_7_12_r;
wire signed [`OutBus]		out_7_12_i;
wire signed [`OutBus]		out_7_13_r;
wire signed [`OutBus]		out_7_13_i;
wire signed [`OutBus]		out_7_14_r;
wire signed [`OutBus]		out_7_14_i;
wire signed [`OutBus]		out_7_15_r;
wire signed [`OutBus]		out_7_15_i;
wire signed [`OutBus]		out_7_16_r;
wire signed [`OutBus]		out_7_16_i;
wire signed [`OutBus]		out_7_17_r;
wire signed [`OutBus]		out_7_17_i;
wire signed [`OutBus]		out_7_18_r;
wire signed [`OutBus]		out_7_18_i;
wire signed [`OutBus]		out_7_19_r;
wire signed [`OutBus]		out_7_19_i;
wire signed [`OutBus]		out_7_20_r;
wire signed [`OutBus]		out_7_20_i;
wire signed [`OutBus]		out_7_21_r;
wire signed [`OutBus]		out_7_21_i;
wire signed [`OutBus]		out_7_22_r;
wire signed [`OutBus]		out_7_22_i;
wire signed [`OutBus]		out_7_23_r;
wire signed [`OutBus]		out_7_23_i;
wire signed [`OutBus]		out_7_24_r;
wire signed [`OutBus]		out_7_24_i;
wire signed [`OutBus]		out_7_25_r;
wire signed [`OutBus]		out_7_25_i;
wire signed [`OutBus]		out_7_26_r;
wire signed [`OutBus]		out_7_26_i;
wire signed [`OutBus]		out_7_27_r;
wire signed [`OutBus]		out_7_27_i;
wire signed [`OutBus]		out_7_28_r;
wire signed [`OutBus]		out_7_28_i;
wire signed [`OutBus]		out_7_29_r;
wire signed [`OutBus]		out_7_29_i;
wire signed [`OutBus]		out_7_30_r;
wire signed [`OutBus]		out_7_30_i;
wire signed [`OutBus]		out_7_31_r;
wire signed [`OutBus]		out_7_31_i;
wire signed [`OutBus]		out_7_32_r;
wire signed [`OutBus]		out_7_32_i;
wire signed [`OutBus]		out_8_1_r;
wire signed [`OutBus]		out_8_1_i;
wire signed [`OutBus]		out_8_2_r;
wire signed [`OutBus]		out_8_2_i;
wire signed [`OutBus]		out_8_3_r;
wire signed [`OutBus]		out_8_3_i;
wire signed [`OutBus]		out_8_4_r;
wire signed [`OutBus]		out_8_4_i;
wire signed [`OutBus]		out_8_5_r;
wire signed [`OutBus]		out_8_5_i;
wire signed [`OutBus]		out_8_6_r;
wire signed [`OutBus]		out_8_6_i;
wire signed [`OutBus]		out_8_7_r;
wire signed [`OutBus]		out_8_7_i;
wire signed [`OutBus]		out_8_8_r;
wire signed [`OutBus]		out_8_8_i;
wire signed [`OutBus]		out_8_9_r;
wire signed [`OutBus]		out_8_9_i;
wire signed [`OutBus]		out_8_10_r;
wire signed [`OutBus]		out_8_10_i;
wire signed [`OutBus]		out_8_11_r;
wire signed [`OutBus]		out_8_11_i;
wire signed [`OutBus]		out_8_12_r;
wire signed [`OutBus]		out_8_12_i;
wire signed [`OutBus]		out_8_13_r;
wire signed [`OutBus]		out_8_13_i;
wire signed [`OutBus]		out_8_14_r;
wire signed [`OutBus]		out_8_14_i;
wire signed [`OutBus]		out_8_15_r;
wire signed [`OutBus]		out_8_15_i;
wire signed [`OutBus]		out_8_16_r;
wire signed [`OutBus]		out_8_16_i;
wire signed [`OutBus]		out_8_17_r;
wire signed [`OutBus]		out_8_17_i;
wire signed [`OutBus]		out_8_18_r;
wire signed [`OutBus]		out_8_18_i;
wire signed [`OutBus]		out_8_19_r;
wire signed [`OutBus]		out_8_19_i;
wire signed [`OutBus]		out_8_20_r;
wire signed [`OutBus]		out_8_20_i;
wire signed [`OutBus]		out_8_21_r;
wire signed [`OutBus]		out_8_21_i;
wire signed [`OutBus]		out_8_22_r;
wire signed [`OutBus]		out_8_22_i;
wire signed [`OutBus]		out_8_23_r;
wire signed [`OutBus]		out_8_23_i;
wire signed [`OutBus]		out_8_24_r;
wire signed [`OutBus]		out_8_24_i;
wire signed [`OutBus]		out_8_25_r;
wire signed [`OutBus]		out_8_25_i;
wire signed [`OutBus]		out_8_26_r;
wire signed [`OutBus]		out_8_26_i;
wire signed [`OutBus]		out_8_27_r;
wire signed [`OutBus]		out_8_27_i;
wire signed [`OutBus]		out_8_28_r;
wire signed [`OutBus]		out_8_28_i;
wire signed [`OutBus]		out_8_29_r;
wire signed [`OutBus]		out_8_29_i;
wire signed [`OutBus]		out_8_30_r;
wire signed [`OutBus]		out_8_30_i;
wire signed [`OutBus]		out_8_31_r;
wire signed [`OutBus]		out_8_31_i;
wire signed [`OutBus]		out_8_32_r;
wire signed [`OutBus]		out_8_32_i;
wire signed [`OutBus]		out_9_1_r;
wire signed [`OutBus]		out_9_1_i;
wire signed [`OutBus]		out_9_2_r;
wire signed [`OutBus]		out_9_2_i;
wire signed [`OutBus]		out_9_3_r;
wire signed [`OutBus]		out_9_3_i;
wire signed [`OutBus]		out_9_4_r;
wire signed [`OutBus]		out_9_4_i;
wire signed [`OutBus]		out_9_5_r;
wire signed [`OutBus]		out_9_5_i;
wire signed [`OutBus]		out_9_6_r;
wire signed [`OutBus]		out_9_6_i;
wire signed [`OutBus]		out_9_7_r;
wire signed [`OutBus]		out_9_7_i;
wire signed [`OutBus]		out_9_8_r;
wire signed [`OutBus]		out_9_8_i;
wire signed [`OutBus]		out_9_9_r;
wire signed [`OutBus]		out_9_9_i;
wire signed [`OutBus]		out_9_10_r;
wire signed [`OutBus]		out_9_10_i;
wire signed [`OutBus]		out_9_11_r;
wire signed [`OutBus]		out_9_11_i;
wire signed [`OutBus]		out_9_12_r;
wire signed [`OutBus]		out_9_12_i;
wire signed [`OutBus]		out_9_13_r;
wire signed [`OutBus]		out_9_13_i;
wire signed [`OutBus]		out_9_14_r;
wire signed [`OutBus]		out_9_14_i;
wire signed [`OutBus]		out_9_15_r;
wire signed [`OutBus]		out_9_15_i;
wire signed [`OutBus]		out_9_16_r;
wire signed [`OutBus]		out_9_16_i;
wire signed [`OutBus]		out_9_17_r;
wire signed [`OutBus]		out_9_17_i;
wire signed [`OutBus]		out_9_18_r;
wire signed [`OutBus]		out_9_18_i;
wire signed [`OutBus]		out_9_19_r;
wire signed [`OutBus]		out_9_19_i;
wire signed [`OutBus]		out_9_20_r;
wire signed [`OutBus]		out_9_20_i;
wire signed [`OutBus]		out_9_21_r;
wire signed [`OutBus]		out_9_21_i;
wire signed [`OutBus]		out_9_22_r;
wire signed [`OutBus]		out_9_22_i;
wire signed [`OutBus]		out_9_23_r;
wire signed [`OutBus]		out_9_23_i;
wire signed [`OutBus]		out_9_24_r;
wire signed [`OutBus]		out_9_24_i;
wire signed [`OutBus]		out_9_25_r;
wire signed [`OutBus]		out_9_25_i;
wire signed [`OutBus]		out_9_26_r;
wire signed [`OutBus]		out_9_26_i;
wire signed [`OutBus]		out_9_27_r;
wire signed [`OutBus]		out_9_27_i;
wire signed [`OutBus]		out_9_28_r;
wire signed [`OutBus]		out_9_28_i;
wire signed [`OutBus]		out_9_29_r;
wire signed [`OutBus]		out_9_29_i;
wire signed [`OutBus]		out_9_30_r;
wire signed [`OutBus]		out_9_30_i;
wire signed [`OutBus]		out_9_31_r;
wire signed [`OutBus]		out_9_31_i;
wire signed [`OutBus]		out_9_32_r;
wire signed [`OutBus]		out_9_32_i;
wire signed [`OutBus]		out_10_1_r;
wire signed [`OutBus]		out_10_1_i;
wire signed [`OutBus]		out_10_2_r;
wire signed [`OutBus]		out_10_2_i;
wire signed [`OutBus]		out_10_3_r;
wire signed [`OutBus]		out_10_3_i;
wire signed [`OutBus]		out_10_4_r;
wire signed [`OutBus]		out_10_4_i;
wire signed [`OutBus]		out_10_5_r;
wire signed [`OutBus]		out_10_5_i;
wire signed [`OutBus]		out_10_6_r;
wire signed [`OutBus]		out_10_6_i;
wire signed [`OutBus]		out_10_7_r;
wire signed [`OutBus]		out_10_7_i;
wire signed [`OutBus]		out_10_8_r;
wire signed [`OutBus]		out_10_8_i;
wire signed [`OutBus]		out_10_9_r;
wire signed [`OutBus]		out_10_9_i;
wire signed [`OutBus]		out_10_10_r;
wire signed [`OutBus]		out_10_10_i;
wire signed [`OutBus]		out_10_11_r;
wire signed [`OutBus]		out_10_11_i;
wire signed [`OutBus]		out_10_12_r;
wire signed [`OutBus]		out_10_12_i;
wire signed [`OutBus]		out_10_13_r;
wire signed [`OutBus]		out_10_13_i;
wire signed [`OutBus]		out_10_14_r;
wire signed [`OutBus]		out_10_14_i;
wire signed [`OutBus]		out_10_15_r;
wire signed [`OutBus]		out_10_15_i;
wire signed [`OutBus]		out_10_16_r;
wire signed [`OutBus]		out_10_16_i;
wire signed [`OutBus]		out_10_17_r;
wire signed [`OutBus]		out_10_17_i;
wire signed [`OutBus]		out_10_18_r;
wire signed [`OutBus]		out_10_18_i;
wire signed [`OutBus]		out_10_19_r;
wire signed [`OutBus]		out_10_19_i;
wire signed [`OutBus]		out_10_20_r;
wire signed [`OutBus]		out_10_20_i;
wire signed [`OutBus]		out_10_21_r;
wire signed [`OutBus]		out_10_21_i;
wire signed [`OutBus]		out_10_22_r;
wire signed [`OutBus]		out_10_22_i;
wire signed [`OutBus]		out_10_23_r;
wire signed [`OutBus]		out_10_23_i;
wire signed [`OutBus]		out_10_24_r;
wire signed [`OutBus]		out_10_24_i;
wire signed [`OutBus]		out_10_25_r;
wire signed [`OutBus]		out_10_25_i;
wire signed [`OutBus]		out_10_26_r;
wire signed [`OutBus]		out_10_26_i;
wire signed [`OutBus]		out_10_27_r;
wire signed [`OutBus]		out_10_27_i;
wire signed [`OutBus]		out_10_28_r;
wire signed [`OutBus]		out_10_28_i;
wire signed [`OutBus]		out_10_29_r;
wire signed [`OutBus]		out_10_29_i;
wire signed [`OutBus]		out_10_30_r;
wire signed [`OutBus]		out_10_30_i;
wire signed [`OutBus]		out_10_31_r;
wire signed [`OutBus]		out_10_31_i;
wire signed [`OutBus]		out_10_32_r;
wire signed [`OutBus]		out_10_32_i;
wire signed [`OutBus]		out_11_1_r;
wire signed [`OutBus]		out_11_1_i;
wire signed [`OutBus]		out_11_2_r;
wire signed [`OutBus]		out_11_2_i;
wire signed [`OutBus]		out_11_3_r;
wire signed [`OutBus]		out_11_3_i;
wire signed [`OutBus]		out_11_4_r;
wire signed [`OutBus]		out_11_4_i;
wire signed [`OutBus]		out_11_5_r;
wire signed [`OutBus]		out_11_5_i;
wire signed [`OutBus]		out_11_6_r;
wire signed [`OutBus]		out_11_6_i;
wire signed [`OutBus]		out_11_7_r;
wire signed [`OutBus]		out_11_7_i;
wire signed [`OutBus]		out_11_8_r;
wire signed [`OutBus]		out_11_8_i;
wire signed [`OutBus]		out_11_9_r;
wire signed [`OutBus]		out_11_9_i;
wire signed [`OutBus]		out_11_10_r;
wire signed [`OutBus]		out_11_10_i;
wire signed [`OutBus]		out_11_11_r;
wire signed [`OutBus]		out_11_11_i;
wire signed [`OutBus]		out_11_12_r;
wire signed [`OutBus]		out_11_12_i;
wire signed [`OutBus]		out_11_13_r;
wire signed [`OutBus]		out_11_13_i;
wire signed [`OutBus]		out_11_14_r;
wire signed [`OutBus]		out_11_14_i;
wire signed [`OutBus]		out_11_15_r;
wire signed [`OutBus]		out_11_15_i;
wire signed [`OutBus]		out_11_16_r;
wire signed [`OutBus]		out_11_16_i;
wire signed [`OutBus]		out_11_17_r;
wire signed [`OutBus]		out_11_17_i;
wire signed [`OutBus]		out_11_18_r;
wire signed [`OutBus]		out_11_18_i;
wire signed [`OutBus]		out_11_19_r;
wire signed [`OutBus]		out_11_19_i;
wire signed [`OutBus]		out_11_20_r;
wire signed [`OutBus]		out_11_20_i;
wire signed [`OutBus]		out_11_21_r;
wire signed [`OutBus]		out_11_21_i;
wire signed [`OutBus]		out_11_22_r;
wire signed [`OutBus]		out_11_22_i;
wire signed [`OutBus]		out_11_23_r;
wire signed [`OutBus]		out_11_23_i;
wire signed [`OutBus]		out_11_24_r;
wire signed [`OutBus]		out_11_24_i;
wire signed [`OutBus]		out_11_25_r;
wire signed [`OutBus]		out_11_25_i;
wire signed [`OutBus]		out_11_26_r;
wire signed [`OutBus]		out_11_26_i;
wire signed [`OutBus]		out_11_27_r;
wire signed [`OutBus]		out_11_27_i;
wire signed [`OutBus]		out_11_28_r;
wire signed [`OutBus]		out_11_28_i;
wire signed [`OutBus]		out_11_29_r;
wire signed [`OutBus]		out_11_29_i;
wire signed [`OutBus]		out_11_30_r;
wire signed [`OutBus]		out_11_30_i;
wire signed [`OutBus]		out_11_31_r;
wire signed [`OutBus]		out_11_31_i;
wire signed [`OutBus]		out_11_32_r;
wire signed [`OutBus]		out_11_32_i;
wire signed [`OutBus]		out_12_1_r;
wire signed [`OutBus]		out_12_1_i;
wire signed [`OutBus]		out_12_2_r;
wire signed [`OutBus]		out_12_2_i;
wire signed [`OutBus]		out_12_3_r;
wire signed [`OutBus]		out_12_3_i;
wire signed [`OutBus]		out_12_4_r;
wire signed [`OutBus]		out_12_4_i;
wire signed [`OutBus]		out_12_5_r;
wire signed [`OutBus]		out_12_5_i;
wire signed [`OutBus]		out_12_6_r;
wire signed [`OutBus]		out_12_6_i;
wire signed [`OutBus]		out_12_7_r;
wire signed [`OutBus]		out_12_7_i;
wire signed [`OutBus]		out_12_8_r;
wire signed [`OutBus]		out_12_8_i;
wire signed [`OutBus]		out_12_9_r;
wire signed [`OutBus]		out_12_9_i;
wire signed [`OutBus]		out_12_10_r;
wire signed [`OutBus]		out_12_10_i;
wire signed [`OutBus]		out_12_11_r;
wire signed [`OutBus]		out_12_11_i;
wire signed [`OutBus]		out_12_12_r;
wire signed [`OutBus]		out_12_12_i;
wire signed [`OutBus]		out_12_13_r;
wire signed [`OutBus]		out_12_13_i;
wire signed [`OutBus]		out_12_14_r;
wire signed [`OutBus]		out_12_14_i;
wire signed [`OutBus]		out_12_15_r;
wire signed [`OutBus]		out_12_15_i;
wire signed [`OutBus]		out_12_16_r;
wire signed [`OutBus]		out_12_16_i;
wire signed [`OutBus]		out_12_17_r;
wire signed [`OutBus]		out_12_17_i;
wire signed [`OutBus]		out_12_18_r;
wire signed [`OutBus]		out_12_18_i;
wire signed [`OutBus]		out_12_19_r;
wire signed [`OutBus]		out_12_19_i;
wire signed [`OutBus]		out_12_20_r;
wire signed [`OutBus]		out_12_20_i;
wire signed [`OutBus]		out_12_21_r;
wire signed [`OutBus]		out_12_21_i;
wire signed [`OutBus]		out_12_22_r;
wire signed [`OutBus]		out_12_22_i;
wire signed [`OutBus]		out_12_23_r;
wire signed [`OutBus]		out_12_23_i;
wire signed [`OutBus]		out_12_24_r;
wire signed [`OutBus]		out_12_24_i;
wire signed [`OutBus]		out_12_25_r;
wire signed [`OutBus]		out_12_25_i;
wire signed [`OutBus]		out_12_26_r;
wire signed [`OutBus]		out_12_26_i;
wire signed [`OutBus]		out_12_27_r;
wire signed [`OutBus]		out_12_27_i;
wire signed [`OutBus]		out_12_28_r;
wire signed [`OutBus]		out_12_28_i;
wire signed [`OutBus]		out_12_29_r;
wire signed [`OutBus]		out_12_29_i;
wire signed [`OutBus]		out_12_30_r;
wire signed [`OutBus]		out_12_30_i;
wire signed [`OutBus]		out_12_31_r;
wire signed [`OutBus]		out_12_31_i;
wire signed [`OutBus]		out_12_32_r;
wire signed [`OutBus]		out_12_32_i;
wire signed [`OutBus]		out_13_1_r;
wire signed [`OutBus]		out_13_1_i;
wire signed [`OutBus]		out_13_2_r;
wire signed [`OutBus]		out_13_2_i;
wire signed [`OutBus]		out_13_3_r;
wire signed [`OutBus]		out_13_3_i;
wire signed [`OutBus]		out_13_4_r;
wire signed [`OutBus]		out_13_4_i;
wire signed [`OutBus]		out_13_5_r;
wire signed [`OutBus]		out_13_5_i;
wire signed [`OutBus]		out_13_6_r;
wire signed [`OutBus]		out_13_6_i;
wire signed [`OutBus]		out_13_7_r;
wire signed [`OutBus]		out_13_7_i;
wire signed [`OutBus]		out_13_8_r;
wire signed [`OutBus]		out_13_8_i;
wire signed [`OutBus]		out_13_9_r;
wire signed [`OutBus]		out_13_9_i;
wire signed [`OutBus]		out_13_10_r;
wire signed [`OutBus]		out_13_10_i;
wire signed [`OutBus]		out_13_11_r;
wire signed [`OutBus]		out_13_11_i;
wire signed [`OutBus]		out_13_12_r;
wire signed [`OutBus]		out_13_12_i;
wire signed [`OutBus]		out_13_13_r;
wire signed [`OutBus]		out_13_13_i;
wire signed [`OutBus]		out_13_14_r;
wire signed [`OutBus]		out_13_14_i;
wire signed [`OutBus]		out_13_15_r;
wire signed [`OutBus]		out_13_15_i;
wire signed [`OutBus]		out_13_16_r;
wire signed [`OutBus]		out_13_16_i;
wire signed [`OutBus]		out_13_17_r;
wire signed [`OutBus]		out_13_17_i;
wire signed [`OutBus]		out_13_18_r;
wire signed [`OutBus]		out_13_18_i;
wire signed [`OutBus]		out_13_19_r;
wire signed [`OutBus]		out_13_19_i;
wire signed [`OutBus]		out_13_20_r;
wire signed [`OutBus]		out_13_20_i;
wire signed [`OutBus]		out_13_21_r;
wire signed [`OutBus]		out_13_21_i;
wire signed [`OutBus]		out_13_22_r;
wire signed [`OutBus]		out_13_22_i;
wire signed [`OutBus]		out_13_23_r;
wire signed [`OutBus]		out_13_23_i;
wire signed [`OutBus]		out_13_24_r;
wire signed [`OutBus]		out_13_24_i;
wire signed [`OutBus]		out_13_25_r;
wire signed [`OutBus]		out_13_25_i;
wire signed [`OutBus]		out_13_26_r;
wire signed [`OutBus]		out_13_26_i;
wire signed [`OutBus]		out_13_27_r;
wire signed [`OutBus]		out_13_27_i;
wire signed [`OutBus]		out_13_28_r;
wire signed [`OutBus]		out_13_28_i;
wire signed [`OutBus]		out_13_29_r;
wire signed [`OutBus]		out_13_29_i;
wire signed [`OutBus]		out_13_30_r;
wire signed [`OutBus]		out_13_30_i;
wire signed [`OutBus]		out_13_31_r;
wire signed [`OutBus]		out_13_31_i;
wire signed [`OutBus]		out_13_32_r;
wire signed [`OutBus]		out_13_32_i;
wire signed [`OutBus]		out_14_1_r;
wire signed [`OutBus]		out_14_1_i;
wire signed [`OutBus]		out_14_2_r;
wire signed [`OutBus]		out_14_2_i;
wire signed [`OutBus]		out_14_3_r;
wire signed [`OutBus]		out_14_3_i;
wire signed [`OutBus]		out_14_4_r;
wire signed [`OutBus]		out_14_4_i;
wire signed [`OutBus]		out_14_5_r;
wire signed [`OutBus]		out_14_5_i;
wire signed [`OutBus]		out_14_6_r;
wire signed [`OutBus]		out_14_6_i;
wire signed [`OutBus]		out_14_7_r;
wire signed [`OutBus]		out_14_7_i;
wire signed [`OutBus]		out_14_8_r;
wire signed [`OutBus]		out_14_8_i;
wire signed [`OutBus]		out_14_9_r;
wire signed [`OutBus]		out_14_9_i;
wire signed [`OutBus]		out_14_10_r;
wire signed [`OutBus]		out_14_10_i;
wire signed [`OutBus]		out_14_11_r;
wire signed [`OutBus]		out_14_11_i;
wire signed [`OutBus]		out_14_12_r;
wire signed [`OutBus]		out_14_12_i;
wire signed [`OutBus]		out_14_13_r;
wire signed [`OutBus]		out_14_13_i;
wire signed [`OutBus]		out_14_14_r;
wire signed [`OutBus]		out_14_14_i;
wire signed [`OutBus]		out_14_15_r;
wire signed [`OutBus]		out_14_15_i;
wire signed [`OutBus]		out_14_16_r;
wire signed [`OutBus]		out_14_16_i;
wire signed [`OutBus]		out_14_17_r;
wire signed [`OutBus]		out_14_17_i;
wire signed [`OutBus]		out_14_18_r;
wire signed [`OutBus]		out_14_18_i;
wire signed [`OutBus]		out_14_19_r;
wire signed [`OutBus]		out_14_19_i;
wire signed [`OutBus]		out_14_20_r;
wire signed [`OutBus]		out_14_20_i;
wire signed [`OutBus]		out_14_21_r;
wire signed [`OutBus]		out_14_21_i;
wire signed [`OutBus]		out_14_22_r;
wire signed [`OutBus]		out_14_22_i;
wire signed [`OutBus]		out_14_23_r;
wire signed [`OutBus]		out_14_23_i;
wire signed [`OutBus]		out_14_24_r;
wire signed [`OutBus]		out_14_24_i;
wire signed [`OutBus]		out_14_25_r;
wire signed [`OutBus]		out_14_25_i;
wire signed [`OutBus]		out_14_26_r;
wire signed [`OutBus]		out_14_26_i;
wire signed [`OutBus]		out_14_27_r;
wire signed [`OutBus]		out_14_27_i;
wire signed [`OutBus]		out_14_28_r;
wire signed [`OutBus]		out_14_28_i;
wire signed [`OutBus]		out_14_29_r;
wire signed [`OutBus]		out_14_29_i;
wire signed [`OutBus]		out_14_30_r;
wire signed [`OutBus]		out_14_30_i;
wire signed [`OutBus]		out_14_31_r;
wire signed [`OutBus]		out_14_31_i;
wire signed [`OutBus]		out_14_32_r;
wire signed [`OutBus]		out_14_32_i;
wire signed [`OutBus]		out_15_1_r;
wire signed [`OutBus]		out_15_1_i;
wire signed [`OutBus]		out_15_2_r;
wire signed [`OutBus]		out_15_2_i;
wire signed [`OutBus]		out_15_3_r;
wire signed [`OutBus]		out_15_3_i;
wire signed [`OutBus]		out_15_4_r;
wire signed [`OutBus]		out_15_4_i;
wire signed [`OutBus]		out_15_5_r;
wire signed [`OutBus]		out_15_5_i;
wire signed [`OutBus]		out_15_6_r;
wire signed [`OutBus]		out_15_6_i;
wire signed [`OutBus]		out_15_7_r;
wire signed [`OutBus]		out_15_7_i;
wire signed [`OutBus]		out_15_8_r;
wire signed [`OutBus]		out_15_8_i;
wire signed [`OutBus]		out_15_9_r;
wire signed [`OutBus]		out_15_9_i;
wire signed [`OutBus]		out_15_10_r;
wire signed [`OutBus]		out_15_10_i;
wire signed [`OutBus]		out_15_11_r;
wire signed [`OutBus]		out_15_11_i;
wire signed [`OutBus]		out_15_12_r;
wire signed [`OutBus]		out_15_12_i;
wire signed [`OutBus]		out_15_13_r;
wire signed [`OutBus]		out_15_13_i;
wire signed [`OutBus]		out_15_14_r;
wire signed [`OutBus]		out_15_14_i;
wire signed [`OutBus]		out_15_15_r;
wire signed [`OutBus]		out_15_15_i;
wire signed [`OutBus]		out_15_16_r;
wire signed [`OutBus]		out_15_16_i;
wire signed [`OutBus]		out_15_17_r;
wire signed [`OutBus]		out_15_17_i;
wire signed [`OutBus]		out_15_18_r;
wire signed [`OutBus]		out_15_18_i;
wire signed [`OutBus]		out_15_19_r;
wire signed [`OutBus]		out_15_19_i;
wire signed [`OutBus]		out_15_20_r;
wire signed [`OutBus]		out_15_20_i;
wire signed [`OutBus]		out_15_21_r;
wire signed [`OutBus]		out_15_21_i;
wire signed [`OutBus]		out_15_22_r;
wire signed [`OutBus]		out_15_22_i;
wire signed [`OutBus]		out_15_23_r;
wire signed [`OutBus]		out_15_23_i;
wire signed [`OutBus]		out_15_24_r;
wire signed [`OutBus]		out_15_24_i;
wire signed [`OutBus]		out_15_25_r;
wire signed [`OutBus]		out_15_25_i;
wire signed [`OutBus]		out_15_26_r;
wire signed [`OutBus]		out_15_26_i;
wire signed [`OutBus]		out_15_27_r;
wire signed [`OutBus]		out_15_27_i;
wire signed [`OutBus]		out_15_28_r;
wire signed [`OutBus]		out_15_28_i;
wire signed [`OutBus]		out_15_29_r;
wire signed [`OutBus]		out_15_29_i;
wire signed [`OutBus]		out_15_30_r;
wire signed [`OutBus]		out_15_30_i;
wire signed [`OutBus]		out_15_31_r;
wire signed [`OutBus]		out_15_31_i;
wire signed [`OutBus]		out_15_32_r;
wire signed [`OutBus]		out_15_32_i;
wire signed [`OutBus]		out_16_1_r;
wire signed [`OutBus]		out_16_1_i;
wire signed [`OutBus]		out_16_2_r;
wire signed [`OutBus]		out_16_2_i;
wire signed [`OutBus]		out_16_3_r;
wire signed [`OutBus]		out_16_3_i;
wire signed [`OutBus]		out_16_4_r;
wire signed [`OutBus]		out_16_4_i;
wire signed [`OutBus]		out_16_5_r;
wire signed [`OutBus]		out_16_5_i;
wire signed [`OutBus]		out_16_6_r;
wire signed [`OutBus]		out_16_6_i;
wire signed [`OutBus]		out_16_7_r;
wire signed [`OutBus]		out_16_7_i;
wire signed [`OutBus]		out_16_8_r;
wire signed [`OutBus]		out_16_8_i;
wire signed [`OutBus]		out_16_9_r;
wire signed [`OutBus]		out_16_9_i;
wire signed [`OutBus]		out_16_10_r;
wire signed [`OutBus]		out_16_10_i;
wire signed [`OutBus]		out_16_11_r;
wire signed [`OutBus]		out_16_11_i;
wire signed [`OutBus]		out_16_12_r;
wire signed [`OutBus]		out_16_12_i;
wire signed [`OutBus]		out_16_13_r;
wire signed [`OutBus]		out_16_13_i;
wire signed [`OutBus]		out_16_14_r;
wire signed [`OutBus]		out_16_14_i;
wire signed [`OutBus]		out_16_15_r;
wire signed [`OutBus]		out_16_15_i;
wire signed [`OutBus]		out_16_16_r;
wire signed [`OutBus]		out_16_16_i;
wire signed [`OutBus]		out_16_17_r;
wire signed [`OutBus]		out_16_17_i;
wire signed [`OutBus]		out_16_18_r;
wire signed [`OutBus]		out_16_18_i;
wire signed [`OutBus]		out_16_19_r;
wire signed [`OutBus]		out_16_19_i;
wire signed [`OutBus]		out_16_20_r;
wire signed [`OutBus]		out_16_20_i;
wire signed [`OutBus]		out_16_21_r;
wire signed [`OutBus]		out_16_21_i;
wire signed [`OutBus]		out_16_22_r;
wire signed [`OutBus]		out_16_22_i;
wire signed [`OutBus]		out_16_23_r;
wire signed [`OutBus]		out_16_23_i;
wire signed [`OutBus]		out_16_24_r;
wire signed [`OutBus]		out_16_24_i;
wire signed [`OutBus]		out_16_25_r;
wire signed [`OutBus]		out_16_25_i;
wire signed [`OutBus]		out_16_26_r;
wire signed [`OutBus]		out_16_26_i;
wire signed [`OutBus]		out_16_27_r;
wire signed [`OutBus]		out_16_27_i;
wire signed [`OutBus]		out_16_28_r;
wire signed [`OutBus]		out_16_28_i;
wire signed [`OutBus]		out_16_29_r;
wire signed [`OutBus]		out_16_29_i;
wire signed [`OutBus]		out_16_30_r;
wire signed [`OutBus]		out_16_30_i;
wire signed [`OutBus]		out_16_31_r;
wire signed [`OutBus]		out_16_31_i;
wire signed [`OutBus]		out_16_32_r;
wire signed [`OutBus]		out_16_32_i;
wire signed [`OutBus]		out_17_1_r;
wire signed [`OutBus]		out_17_1_i;
wire signed [`OutBus]		out_17_2_r;
wire signed [`OutBus]		out_17_2_i;
wire signed [`OutBus]		out_17_3_r;
wire signed [`OutBus]		out_17_3_i;
wire signed [`OutBus]		out_17_4_r;
wire signed [`OutBus]		out_17_4_i;
wire signed [`OutBus]		out_17_5_r;
wire signed [`OutBus]		out_17_5_i;
wire signed [`OutBus]		out_17_6_r;
wire signed [`OutBus]		out_17_6_i;
wire signed [`OutBus]		out_17_7_r;
wire signed [`OutBus]		out_17_7_i;
wire signed [`OutBus]		out_17_8_r;
wire signed [`OutBus]		out_17_8_i;
wire signed [`OutBus]		out_17_9_r;
wire signed [`OutBus]		out_17_9_i;
wire signed [`OutBus]		out_17_10_r;
wire signed [`OutBus]		out_17_10_i;
wire signed [`OutBus]		out_17_11_r;
wire signed [`OutBus]		out_17_11_i;
wire signed [`OutBus]		out_17_12_r;
wire signed [`OutBus]		out_17_12_i;
wire signed [`OutBus]		out_17_13_r;
wire signed [`OutBus]		out_17_13_i;
wire signed [`OutBus]		out_17_14_r;
wire signed [`OutBus]		out_17_14_i;
wire signed [`OutBus]		out_17_15_r;
wire signed [`OutBus]		out_17_15_i;
wire signed [`OutBus]		out_17_16_r;
wire signed [`OutBus]		out_17_16_i;
wire signed [`OutBus]		out_17_17_r;
wire signed [`OutBus]		out_17_17_i;
wire signed [`OutBus]		out_17_18_r;
wire signed [`OutBus]		out_17_18_i;
wire signed [`OutBus]		out_17_19_r;
wire signed [`OutBus]		out_17_19_i;
wire signed [`OutBus]		out_17_20_r;
wire signed [`OutBus]		out_17_20_i;
wire signed [`OutBus]		out_17_21_r;
wire signed [`OutBus]		out_17_21_i;
wire signed [`OutBus]		out_17_22_r;
wire signed [`OutBus]		out_17_22_i;
wire signed [`OutBus]		out_17_23_r;
wire signed [`OutBus]		out_17_23_i;
wire signed [`OutBus]		out_17_24_r;
wire signed [`OutBus]		out_17_24_i;
wire signed [`OutBus]		out_17_25_r;
wire signed [`OutBus]		out_17_25_i;
wire signed [`OutBus]		out_17_26_r;
wire signed [`OutBus]		out_17_26_i;
wire signed [`OutBus]		out_17_27_r;
wire signed [`OutBus]		out_17_27_i;
wire signed [`OutBus]		out_17_28_r;
wire signed [`OutBus]		out_17_28_i;
wire signed [`OutBus]		out_17_29_r;
wire signed [`OutBus]		out_17_29_i;
wire signed [`OutBus]		out_17_30_r;
wire signed [`OutBus]		out_17_30_i;
wire signed [`OutBus]		out_17_31_r;
wire signed [`OutBus]		out_17_31_i;
wire signed [`OutBus]		out_17_32_r;
wire signed [`OutBus]		out_17_32_i;
wire signed [`OutBus]		out_18_1_r;
wire signed [`OutBus]		out_18_1_i;
wire signed [`OutBus]		out_18_2_r;
wire signed [`OutBus]		out_18_2_i;
wire signed [`OutBus]		out_18_3_r;
wire signed [`OutBus]		out_18_3_i;
wire signed [`OutBus]		out_18_4_r;
wire signed [`OutBus]		out_18_4_i;
wire signed [`OutBus]		out_18_5_r;
wire signed [`OutBus]		out_18_5_i;
wire signed [`OutBus]		out_18_6_r;
wire signed [`OutBus]		out_18_6_i;
wire signed [`OutBus]		out_18_7_r;
wire signed [`OutBus]		out_18_7_i;
wire signed [`OutBus]		out_18_8_r;
wire signed [`OutBus]		out_18_8_i;
wire signed [`OutBus]		out_18_9_r;
wire signed [`OutBus]		out_18_9_i;
wire signed [`OutBus]		out_18_10_r;
wire signed [`OutBus]		out_18_10_i;
wire signed [`OutBus]		out_18_11_r;
wire signed [`OutBus]		out_18_11_i;
wire signed [`OutBus]		out_18_12_r;
wire signed [`OutBus]		out_18_12_i;
wire signed [`OutBus]		out_18_13_r;
wire signed [`OutBus]		out_18_13_i;
wire signed [`OutBus]		out_18_14_r;
wire signed [`OutBus]		out_18_14_i;
wire signed [`OutBus]		out_18_15_r;
wire signed [`OutBus]		out_18_15_i;
wire signed [`OutBus]		out_18_16_r;
wire signed [`OutBus]		out_18_16_i;
wire signed [`OutBus]		out_18_17_r;
wire signed [`OutBus]		out_18_17_i;
wire signed [`OutBus]		out_18_18_r;
wire signed [`OutBus]		out_18_18_i;
wire signed [`OutBus]		out_18_19_r;
wire signed [`OutBus]		out_18_19_i;
wire signed [`OutBus]		out_18_20_r;
wire signed [`OutBus]		out_18_20_i;
wire signed [`OutBus]		out_18_21_r;
wire signed [`OutBus]		out_18_21_i;
wire signed [`OutBus]		out_18_22_r;
wire signed [`OutBus]		out_18_22_i;
wire signed [`OutBus]		out_18_23_r;
wire signed [`OutBus]		out_18_23_i;
wire signed [`OutBus]		out_18_24_r;
wire signed [`OutBus]		out_18_24_i;
wire signed [`OutBus]		out_18_25_r;
wire signed [`OutBus]		out_18_25_i;
wire signed [`OutBus]		out_18_26_r;
wire signed [`OutBus]		out_18_26_i;
wire signed [`OutBus]		out_18_27_r;
wire signed [`OutBus]		out_18_27_i;
wire signed [`OutBus]		out_18_28_r;
wire signed [`OutBus]		out_18_28_i;
wire signed [`OutBus]		out_18_29_r;
wire signed [`OutBus]		out_18_29_i;
wire signed [`OutBus]		out_18_30_r;
wire signed [`OutBus]		out_18_30_i;
wire signed [`OutBus]		out_18_31_r;
wire signed [`OutBus]		out_18_31_i;
wire signed [`OutBus]		out_18_32_r;
wire signed [`OutBus]		out_18_32_i;
wire signed [`OutBus]		out_19_1_r;
wire signed [`OutBus]		out_19_1_i;
wire signed [`OutBus]		out_19_2_r;
wire signed [`OutBus]		out_19_2_i;
wire signed [`OutBus]		out_19_3_r;
wire signed [`OutBus]		out_19_3_i;
wire signed [`OutBus]		out_19_4_r;
wire signed [`OutBus]		out_19_4_i;
wire signed [`OutBus]		out_19_5_r;
wire signed [`OutBus]		out_19_5_i;
wire signed [`OutBus]		out_19_6_r;
wire signed [`OutBus]		out_19_6_i;
wire signed [`OutBus]		out_19_7_r;
wire signed [`OutBus]		out_19_7_i;
wire signed [`OutBus]		out_19_8_r;
wire signed [`OutBus]		out_19_8_i;
wire signed [`OutBus]		out_19_9_r;
wire signed [`OutBus]		out_19_9_i;
wire signed [`OutBus]		out_19_10_r;
wire signed [`OutBus]		out_19_10_i;
wire signed [`OutBus]		out_19_11_r;
wire signed [`OutBus]		out_19_11_i;
wire signed [`OutBus]		out_19_12_r;
wire signed [`OutBus]		out_19_12_i;
wire signed [`OutBus]		out_19_13_r;
wire signed [`OutBus]		out_19_13_i;
wire signed [`OutBus]		out_19_14_r;
wire signed [`OutBus]		out_19_14_i;
wire signed [`OutBus]		out_19_15_r;
wire signed [`OutBus]		out_19_15_i;
wire signed [`OutBus]		out_19_16_r;
wire signed [`OutBus]		out_19_16_i;
wire signed [`OutBus]		out_19_17_r;
wire signed [`OutBus]		out_19_17_i;
wire signed [`OutBus]		out_19_18_r;
wire signed [`OutBus]		out_19_18_i;
wire signed [`OutBus]		out_19_19_r;
wire signed [`OutBus]		out_19_19_i;
wire signed [`OutBus]		out_19_20_r;
wire signed [`OutBus]		out_19_20_i;
wire signed [`OutBus]		out_19_21_r;
wire signed [`OutBus]		out_19_21_i;
wire signed [`OutBus]		out_19_22_r;
wire signed [`OutBus]		out_19_22_i;
wire signed [`OutBus]		out_19_23_r;
wire signed [`OutBus]		out_19_23_i;
wire signed [`OutBus]		out_19_24_r;
wire signed [`OutBus]		out_19_24_i;
wire signed [`OutBus]		out_19_25_r;
wire signed [`OutBus]		out_19_25_i;
wire signed [`OutBus]		out_19_26_r;
wire signed [`OutBus]		out_19_26_i;
wire signed [`OutBus]		out_19_27_r;
wire signed [`OutBus]		out_19_27_i;
wire signed [`OutBus]		out_19_28_r;
wire signed [`OutBus]		out_19_28_i;
wire signed [`OutBus]		out_19_29_r;
wire signed [`OutBus]		out_19_29_i;
wire signed [`OutBus]		out_19_30_r;
wire signed [`OutBus]		out_19_30_i;
wire signed [`OutBus]		out_19_31_r;
wire signed [`OutBus]		out_19_31_i;
wire signed [`OutBus]		out_19_32_r;
wire signed [`OutBus]		out_19_32_i;
wire signed [`OutBus]		out_20_1_r;
wire signed [`OutBus]		out_20_1_i;
wire signed [`OutBus]		out_20_2_r;
wire signed [`OutBus]		out_20_2_i;
wire signed [`OutBus]		out_20_3_r;
wire signed [`OutBus]		out_20_3_i;
wire signed [`OutBus]		out_20_4_r;
wire signed [`OutBus]		out_20_4_i;
wire signed [`OutBus]		out_20_5_r;
wire signed [`OutBus]		out_20_5_i;
wire signed [`OutBus]		out_20_6_r;
wire signed [`OutBus]		out_20_6_i;
wire signed [`OutBus]		out_20_7_r;
wire signed [`OutBus]		out_20_7_i;
wire signed [`OutBus]		out_20_8_r;
wire signed [`OutBus]		out_20_8_i;
wire signed [`OutBus]		out_20_9_r;
wire signed [`OutBus]		out_20_9_i;
wire signed [`OutBus]		out_20_10_r;
wire signed [`OutBus]		out_20_10_i;
wire signed [`OutBus]		out_20_11_r;
wire signed [`OutBus]		out_20_11_i;
wire signed [`OutBus]		out_20_12_r;
wire signed [`OutBus]		out_20_12_i;
wire signed [`OutBus]		out_20_13_r;
wire signed [`OutBus]		out_20_13_i;
wire signed [`OutBus]		out_20_14_r;
wire signed [`OutBus]		out_20_14_i;
wire signed [`OutBus]		out_20_15_r;
wire signed [`OutBus]		out_20_15_i;
wire signed [`OutBus]		out_20_16_r;
wire signed [`OutBus]		out_20_16_i;
wire signed [`OutBus]		out_20_17_r;
wire signed [`OutBus]		out_20_17_i;
wire signed [`OutBus]		out_20_18_r;
wire signed [`OutBus]		out_20_18_i;
wire signed [`OutBus]		out_20_19_r;
wire signed [`OutBus]		out_20_19_i;
wire signed [`OutBus]		out_20_20_r;
wire signed [`OutBus]		out_20_20_i;
wire signed [`OutBus]		out_20_21_r;
wire signed [`OutBus]		out_20_21_i;
wire signed [`OutBus]		out_20_22_r;
wire signed [`OutBus]		out_20_22_i;
wire signed [`OutBus]		out_20_23_r;
wire signed [`OutBus]		out_20_23_i;
wire signed [`OutBus]		out_20_24_r;
wire signed [`OutBus]		out_20_24_i;
wire signed [`OutBus]		out_20_25_r;
wire signed [`OutBus]		out_20_25_i;
wire signed [`OutBus]		out_20_26_r;
wire signed [`OutBus]		out_20_26_i;
wire signed [`OutBus]		out_20_27_r;
wire signed [`OutBus]		out_20_27_i;
wire signed [`OutBus]		out_20_28_r;
wire signed [`OutBus]		out_20_28_i;
wire signed [`OutBus]		out_20_29_r;
wire signed [`OutBus]		out_20_29_i;
wire signed [`OutBus]		out_20_30_r;
wire signed [`OutBus]		out_20_30_i;
wire signed [`OutBus]		out_20_31_r;
wire signed [`OutBus]		out_20_31_i;
wire signed [`OutBus]		out_20_32_r;
wire signed [`OutBus]		out_20_32_i;
wire signed [`OutBus]		out_21_1_r;
wire signed [`OutBus]		out_21_1_i;
wire signed [`OutBus]		out_21_2_r;
wire signed [`OutBus]		out_21_2_i;
wire signed [`OutBus]		out_21_3_r;
wire signed [`OutBus]		out_21_3_i;
wire signed [`OutBus]		out_21_4_r;
wire signed [`OutBus]		out_21_4_i;
wire signed [`OutBus]		out_21_5_r;
wire signed [`OutBus]		out_21_5_i;
wire signed [`OutBus]		out_21_6_r;
wire signed [`OutBus]		out_21_6_i;
wire signed [`OutBus]		out_21_7_r;
wire signed [`OutBus]		out_21_7_i;
wire signed [`OutBus]		out_21_8_r;
wire signed [`OutBus]		out_21_8_i;
wire signed [`OutBus]		out_21_9_r;
wire signed [`OutBus]		out_21_9_i;
wire signed [`OutBus]		out_21_10_r;
wire signed [`OutBus]		out_21_10_i;
wire signed [`OutBus]		out_21_11_r;
wire signed [`OutBus]		out_21_11_i;
wire signed [`OutBus]		out_21_12_r;
wire signed [`OutBus]		out_21_12_i;
wire signed [`OutBus]		out_21_13_r;
wire signed [`OutBus]		out_21_13_i;
wire signed [`OutBus]		out_21_14_r;
wire signed [`OutBus]		out_21_14_i;
wire signed [`OutBus]		out_21_15_r;
wire signed [`OutBus]		out_21_15_i;
wire signed [`OutBus]		out_21_16_r;
wire signed [`OutBus]		out_21_16_i;
wire signed [`OutBus]		out_21_17_r;
wire signed [`OutBus]		out_21_17_i;
wire signed [`OutBus]		out_21_18_r;
wire signed [`OutBus]		out_21_18_i;
wire signed [`OutBus]		out_21_19_r;
wire signed [`OutBus]		out_21_19_i;
wire signed [`OutBus]		out_21_20_r;
wire signed [`OutBus]		out_21_20_i;
wire signed [`OutBus]		out_21_21_r;
wire signed [`OutBus]		out_21_21_i;
wire signed [`OutBus]		out_21_22_r;
wire signed [`OutBus]		out_21_22_i;
wire signed [`OutBus]		out_21_23_r;
wire signed [`OutBus]		out_21_23_i;
wire signed [`OutBus]		out_21_24_r;
wire signed [`OutBus]		out_21_24_i;
wire signed [`OutBus]		out_21_25_r;
wire signed [`OutBus]		out_21_25_i;
wire signed [`OutBus]		out_21_26_r;
wire signed [`OutBus]		out_21_26_i;
wire signed [`OutBus]		out_21_27_r;
wire signed [`OutBus]		out_21_27_i;
wire signed [`OutBus]		out_21_28_r;
wire signed [`OutBus]		out_21_28_i;
wire signed [`OutBus]		out_21_29_r;
wire signed [`OutBus]		out_21_29_i;
wire signed [`OutBus]		out_21_30_r;
wire signed [`OutBus]		out_21_30_i;
wire signed [`OutBus]		out_21_31_r;
wire signed [`OutBus]		out_21_31_i;
wire signed [`OutBus]		out_21_32_r;
wire signed [`OutBus]		out_21_32_i;
wire signed [`OutBus]		out_22_1_r;
wire signed [`OutBus]		out_22_1_i;
wire signed [`OutBus]		out_22_2_r;
wire signed [`OutBus]		out_22_2_i;
wire signed [`OutBus]		out_22_3_r;
wire signed [`OutBus]		out_22_3_i;
wire signed [`OutBus]		out_22_4_r;
wire signed [`OutBus]		out_22_4_i;
wire signed [`OutBus]		out_22_5_r;
wire signed [`OutBus]		out_22_5_i;
wire signed [`OutBus]		out_22_6_r;
wire signed [`OutBus]		out_22_6_i;
wire signed [`OutBus]		out_22_7_r;
wire signed [`OutBus]		out_22_7_i;
wire signed [`OutBus]		out_22_8_r;
wire signed [`OutBus]		out_22_8_i;
wire signed [`OutBus]		out_22_9_r;
wire signed [`OutBus]		out_22_9_i;
wire signed [`OutBus]		out_22_10_r;
wire signed [`OutBus]		out_22_10_i;
wire signed [`OutBus]		out_22_11_r;
wire signed [`OutBus]		out_22_11_i;
wire signed [`OutBus]		out_22_12_r;
wire signed [`OutBus]		out_22_12_i;
wire signed [`OutBus]		out_22_13_r;
wire signed [`OutBus]		out_22_13_i;
wire signed [`OutBus]		out_22_14_r;
wire signed [`OutBus]		out_22_14_i;
wire signed [`OutBus]		out_22_15_r;
wire signed [`OutBus]		out_22_15_i;
wire signed [`OutBus]		out_22_16_r;
wire signed [`OutBus]		out_22_16_i;
wire signed [`OutBus]		out_22_17_r;
wire signed [`OutBus]		out_22_17_i;
wire signed [`OutBus]		out_22_18_r;
wire signed [`OutBus]		out_22_18_i;
wire signed [`OutBus]		out_22_19_r;
wire signed [`OutBus]		out_22_19_i;
wire signed [`OutBus]		out_22_20_r;
wire signed [`OutBus]		out_22_20_i;
wire signed [`OutBus]		out_22_21_r;
wire signed [`OutBus]		out_22_21_i;
wire signed [`OutBus]		out_22_22_r;
wire signed [`OutBus]		out_22_22_i;
wire signed [`OutBus]		out_22_23_r;
wire signed [`OutBus]		out_22_23_i;
wire signed [`OutBus]		out_22_24_r;
wire signed [`OutBus]		out_22_24_i;
wire signed [`OutBus]		out_22_25_r;
wire signed [`OutBus]		out_22_25_i;
wire signed [`OutBus]		out_22_26_r;
wire signed [`OutBus]		out_22_26_i;
wire signed [`OutBus]		out_22_27_r;
wire signed [`OutBus]		out_22_27_i;
wire signed [`OutBus]		out_22_28_r;
wire signed [`OutBus]		out_22_28_i;
wire signed [`OutBus]		out_22_29_r;
wire signed [`OutBus]		out_22_29_i;
wire signed [`OutBus]		out_22_30_r;
wire signed [`OutBus]		out_22_30_i;
wire signed [`OutBus]		out_22_31_r;
wire signed [`OutBus]		out_22_31_i;
wire signed [`OutBus]		out_22_32_r;
wire signed [`OutBus]		out_22_32_i;
wire signed [`OutBus]		out_23_1_r;
wire signed [`OutBus]		out_23_1_i;
wire signed [`OutBus]		out_23_2_r;
wire signed [`OutBus]		out_23_2_i;
wire signed [`OutBus]		out_23_3_r;
wire signed [`OutBus]		out_23_3_i;
wire signed [`OutBus]		out_23_4_r;
wire signed [`OutBus]		out_23_4_i;
wire signed [`OutBus]		out_23_5_r;
wire signed [`OutBus]		out_23_5_i;
wire signed [`OutBus]		out_23_6_r;
wire signed [`OutBus]		out_23_6_i;
wire signed [`OutBus]		out_23_7_r;
wire signed [`OutBus]		out_23_7_i;
wire signed [`OutBus]		out_23_8_r;
wire signed [`OutBus]		out_23_8_i;
wire signed [`OutBus]		out_23_9_r;
wire signed [`OutBus]		out_23_9_i;
wire signed [`OutBus]		out_23_10_r;
wire signed [`OutBus]		out_23_10_i;
wire signed [`OutBus]		out_23_11_r;
wire signed [`OutBus]		out_23_11_i;
wire signed [`OutBus]		out_23_12_r;
wire signed [`OutBus]		out_23_12_i;
wire signed [`OutBus]		out_23_13_r;
wire signed [`OutBus]		out_23_13_i;
wire signed [`OutBus]		out_23_14_r;
wire signed [`OutBus]		out_23_14_i;
wire signed [`OutBus]		out_23_15_r;
wire signed [`OutBus]		out_23_15_i;
wire signed [`OutBus]		out_23_16_r;
wire signed [`OutBus]		out_23_16_i;
wire signed [`OutBus]		out_23_17_r;
wire signed [`OutBus]		out_23_17_i;
wire signed [`OutBus]		out_23_18_r;
wire signed [`OutBus]		out_23_18_i;
wire signed [`OutBus]		out_23_19_r;
wire signed [`OutBus]		out_23_19_i;
wire signed [`OutBus]		out_23_20_r;
wire signed [`OutBus]		out_23_20_i;
wire signed [`OutBus]		out_23_21_r;
wire signed [`OutBus]		out_23_21_i;
wire signed [`OutBus]		out_23_22_r;
wire signed [`OutBus]		out_23_22_i;
wire signed [`OutBus]		out_23_23_r;
wire signed [`OutBus]		out_23_23_i;
wire signed [`OutBus]		out_23_24_r;
wire signed [`OutBus]		out_23_24_i;
wire signed [`OutBus]		out_23_25_r;
wire signed [`OutBus]		out_23_25_i;
wire signed [`OutBus]		out_23_26_r;
wire signed [`OutBus]		out_23_26_i;
wire signed [`OutBus]		out_23_27_r;
wire signed [`OutBus]		out_23_27_i;
wire signed [`OutBus]		out_23_28_r;
wire signed [`OutBus]		out_23_28_i;
wire signed [`OutBus]		out_23_29_r;
wire signed [`OutBus]		out_23_29_i;
wire signed [`OutBus]		out_23_30_r;
wire signed [`OutBus]		out_23_30_i;
wire signed [`OutBus]		out_23_31_r;
wire signed [`OutBus]		out_23_31_i;
wire signed [`OutBus]		out_23_32_r;
wire signed [`OutBus]		out_23_32_i;
wire signed [`OutBus]		out_24_1_r;
wire signed [`OutBus]		out_24_1_i;
wire signed [`OutBus]		out_24_2_r;
wire signed [`OutBus]		out_24_2_i;
wire signed [`OutBus]		out_24_3_r;
wire signed [`OutBus]		out_24_3_i;
wire signed [`OutBus]		out_24_4_r;
wire signed [`OutBus]		out_24_4_i;
wire signed [`OutBus]		out_24_5_r;
wire signed [`OutBus]		out_24_5_i;
wire signed [`OutBus]		out_24_6_r;
wire signed [`OutBus]		out_24_6_i;
wire signed [`OutBus]		out_24_7_r;
wire signed [`OutBus]		out_24_7_i;
wire signed [`OutBus]		out_24_8_r;
wire signed [`OutBus]		out_24_8_i;
wire signed [`OutBus]		out_24_9_r;
wire signed [`OutBus]		out_24_9_i;
wire signed [`OutBus]		out_24_10_r;
wire signed [`OutBus]		out_24_10_i;
wire signed [`OutBus]		out_24_11_r;
wire signed [`OutBus]		out_24_11_i;
wire signed [`OutBus]		out_24_12_r;
wire signed [`OutBus]		out_24_12_i;
wire signed [`OutBus]		out_24_13_r;
wire signed [`OutBus]		out_24_13_i;
wire signed [`OutBus]		out_24_14_r;
wire signed [`OutBus]		out_24_14_i;
wire signed [`OutBus]		out_24_15_r;
wire signed [`OutBus]		out_24_15_i;
wire signed [`OutBus]		out_24_16_r;
wire signed [`OutBus]		out_24_16_i;
wire signed [`OutBus]		out_24_17_r;
wire signed [`OutBus]		out_24_17_i;
wire signed [`OutBus]		out_24_18_r;
wire signed [`OutBus]		out_24_18_i;
wire signed [`OutBus]		out_24_19_r;
wire signed [`OutBus]		out_24_19_i;
wire signed [`OutBus]		out_24_20_r;
wire signed [`OutBus]		out_24_20_i;
wire signed [`OutBus]		out_24_21_r;
wire signed [`OutBus]		out_24_21_i;
wire signed [`OutBus]		out_24_22_r;
wire signed [`OutBus]		out_24_22_i;
wire signed [`OutBus]		out_24_23_r;
wire signed [`OutBus]		out_24_23_i;
wire signed [`OutBus]		out_24_24_r;
wire signed [`OutBus]		out_24_24_i;
wire signed [`OutBus]		out_24_25_r;
wire signed [`OutBus]		out_24_25_i;
wire signed [`OutBus]		out_24_26_r;
wire signed [`OutBus]		out_24_26_i;
wire signed [`OutBus]		out_24_27_r;
wire signed [`OutBus]		out_24_27_i;
wire signed [`OutBus]		out_24_28_r;
wire signed [`OutBus]		out_24_28_i;
wire signed [`OutBus]		out_24_29_r;
wire signed [`OutBus]		out_24_29_i;
wire signed [`OutBus]		out_24_30_r;
wire signed [`OutBus]		out_24_30_i;
wire signed [`OutBus]		out_24_31_r;
wire signed [`OutBus]		out_24_31_i;
wire signed [`OutBus]		out_24_32_r;
wire signed [`OutBus]		out_24_32_i;
wire signed [`OutBus]		out_25_1_r;
wire signed [`OutBus]		out_25_1_i;
wire signed [`OutBus]		out_25_2_r;
wire signed [`OutBus]		out_25_2_i;
wire signed [`OutBus]		out_25_3_r;
wire signed [`OutBus]		out_25_3_i;
wire signed [`OutBus]		out_25_4_r;
wire signed [`OutBus]		out_25_4_i;
wire signed [`OutBus]		out_25_5_r;
wire signed [`OutBus]		out_25_5_i;
wire signed [`OutBus]		out_25_6_r;
wire signed [`OutBus]		out_25_6_i;
wire signed [`OutBus]		out_25_7_r;
wire signed [`OutBus]		out_25_7_i;
wire signed [`OutBus]		out_25_8_r;
wire signed [`OutBus]		out_25_8_i;
wire signed [`OutBus]		out_25_9_r;
wire signed [`OutBus]		out_25_9_i;
wire signed [`OutBus]		out_25_10_r;
wire signed [`OutBus]		out_25_10_i;
wire signed [`OutBus]		out_25_11_r;
wire signed [`OutBus]		out_25_11_i;
wire signed [`OutBus]		out_25_12_r;
wire signed [`OutBus]		out_25_12_i;
wire signed [`OutBus]		out_25_13_r;
wire signed [`OutBus]		out_25_13_i;
wire signed [`OutBus]		out_25_14_r;
wire signed [`OutBus]		out_25_14_i;
wire signed [`OutBus]		out_25_15_r;
wire signed [`OutBus]		out_25_15_i;
wire signed [`OutBus]		out_25_16_r;
wire signed [`OutBus]		out_25_16_i;
wire signed [`OutBus]		out_25_17_r;
wire signed [`OutBus]		out_25_17_i;
wire signed [`OutBus]		out_25_18_r;
wire signed [`OutBus]		out_25_18_i;
wire signed [`OutBus]		out_25_19_r;
wire signed [`OutBus]		out_25_19_i;
wire signed [`OutBus]		out_25_20_r;
wire signed [`OutBus]		out_25_20_i;
wire signed [`OutBus]		out_25_21_r;
wire signed [`OutBus]		out_25_21_i;
wire signed [`OutBus]		out_25_22_r;
wire signed [`OutBus]		out_25_22_i;
wire signed [`OutBus]		out_25_23_r;
wire signed [`OutBus]		out_25_23_i;
wire signed [`OutBus]		out_25_24_r;
wire signed [`OutBus]		out_25_24_i;
wire signed [`OutBus]		out_25_25_r;
wire signed [`OutBus]		out_25_25_i;
wire signed [`OutBus]		out_25_26_r;
wire signed [`OutBus]		out_25_26_i;
wire signed [`OutBus]		out_25_27_r;
wire signed [`OutBus]		out_25_27_i;
wire signed [`OutBus]		out_25_28_r;
wire signed [`OutBus]		out_25_28_i;
wire signed [`OutBus]		out_25_29_r;
wire signed [`OutBus]		out_25_29_i;
wire signed [`OutBus]		out_25_30_r;
wire signed [`OutBus]		out_25_30_i;
wire signed [`OutBus]		out_25_31_r;
wire signed [`OutBus]		out_25_31_i;
wire signed [`OutBus]		out_25_32_r;
wire signed [`OutBus]		out_25_32_i;
wire signed [`OutBus]		out_26_1_r;
wire signed [`OutBus]		out_26_1_i;
wire signed [`OutBus]		out_26_2_r;
wire signed [`OutBus]		out_26_2_i;
wire signed [`OutBus]		out_26_3_r;
wire signed [`OutBus]		out_26_3_i;
wire signed [`OutBus]		out_26_4_r;
wire signed [`OutBus]		out_26_4_i;
wire signed [`OutBus]		out_26_5_r;
wire signed [`OutBus]		out_26_5_i;
wire signed [`OutBus]		out_26_6_r;
wire signed [`OutBus]		out_26_6_i;
wire signed [`OutBus]		out_26_7_r;
wire signed [`OutBus]		out_26_7_i;
wire signed [`OutBus]		out_26_8_r;
wire signed [`OutBus]		out_26_8_i;
wire signed [`OutBus]		out_26_9_r;
wire signed [`OutBus]		out_26_9_i;
wire signed [`OutBus]		out_26_10_r;
wire signed [`OutBus]		out_26_10_i;
wire signed [`OutBus]		out_26_11_r;
wire signed [`OutBus]		out_26_11_i;
wire signed [`OutBus]		out_26_12_r;
wire signed [`OutBus]		out_26_12_i;
wire signed [`OutBus]		out_26_13_r;
wire signed [`OutBus]		out_26_13_i;
wire signed [`OutBus]		out_26_14_r;
wire signed [`OutBus]		out_26_14_i;
wire signed [`OutBus]		out_26_15_r;
wire signed [`OutBus]		out_26_15_i;
wire signed [`OutBus]		out_26_16_r;
wire signed [`OutBus]		out_26_16_i;
wire signed [`OutBus]		out_26_17_r;
wire signed [`OutBus]		out_26_17_i;
wire signed [`OutBus]		out_26_18_r;
wire signed [`OutBus]		out_26_18_i;
wire signed [`OutBus]		out_26_19_r;
wire signed [`OutBus]		out_26_19_i;
wire signed [`OutBus]		out_26_20_r;
wire signed [`OutBus]		out_26_20_i;
wire signed [`OutBus]		out_26_21_r;
wire signed [`OutBus]		out_26_21_i;
wire signed [`OutBus]		out_26_22_r;
wire signed [`OutBus]		out_26_22_i;
wire signed [`OutBus]		out_26_23_r;
wire signed [`OutBus]		out_26_23_i;
wire signed [`OutBus]		out_26_24_r;
wire signed [`OutBus]		out_26_24_i;
wire signed [`OutBus]		out_26_25_r;
wire signed [`OutBus]		out_26_25_i;
wire signed [`OutBus]		out_26_26_r;
wire signed [`OutBus]		out_26_26_i;
wire signed [`OutBus]		out_26_27_r;
wire signed [`OutBus]		out_26_27_i;
wire signed [`OutBus]		out_26_28_r;
wire signed [`OutBus]		out_26_28_i;
wire signed [`OutBus]		out_26_29_r;
wire signed [`OutBus]		out_26_29_i;
wire signed [`OutBus]		out_26_30_r;
wire signed [`OutBus]		out_26_30_i;
wire signed [`OutBus]		out_26_31_r;
wire signed [`OutBus]		out_26_31_i;
wire signed [`OutBus]		out_26_32_r;
wire signed [`OutBus]		out_26_32_i;
wire signed [`OutBus]		out_27_1_r;
wire signed [`OutBus]		out_27_1_i;
wire signed [`OutBus]		out_27_2_r;
wire signed [`OutBus]		out_27_2_i;
wire signed [`OutBus]		out_27_3_r;
wire signed [`OutBus]		out_27_3_i;
wire signed [`OutBus]		out_27_4_r;
wire signed [`OutBus]		out_27_4_i;
wire signed [`OutBus]		out_27_5_r;
wire signed [`OutBus]		out_27_5_i;
wire signed [`OutBus]		out_27_6_r;
wire signed [`OutBus]		out_27_6_i;
wire signed [`OutBus]		out_27_7_r;
wire signed [`OutBus]		out_27_7_i;
wire signed [`OutBus]		out_27_8_r;
wire signed [`OutBus]		out_27_8_i;
wire signed [`OutBus]		out_27_9_r;
wire signed [`OutBus]		out_27_9_i;
wire signed [`OutBus]		out_27_10_r;
wire signed [`OutBus]		out_27_10_i;
wire signed [`OutBus]		out_27_11_r;
wire signed [`OutBus]		out_27_11_i;
wire signed [`OutBus]		out_27_12_r;
wire signed [`OutBus]		out_27_12_i;
wire signed [`OutBus]		out_27_13_r;
wire signed [`OutBus]		out_27_13_i;
wire signed [`OutBus]		out_27_14_r;
wire signed [`OutBus]		out_27_14_i;
wire signed [`OutBus]		out_27_15_r;
wire signed [`OutBus]		out_27_15_i;
wire signed [`OutBus]		out_27_16_r;
wire signed [`OutBus]		out_27_16_i;
wire signed [`OutBus]		out_27_17_r;
wire signed [`OutBus]		out_27_17_i;
wire signed [`OutBus]		out_27_18_r;
wire signed [`OutBus]		out_27_18_i;
wire signed [`OutBus]		out_27_19_r;
wire signed [`OutBus]		out_27_19_i;
wire signed [`OutBus]		out_27_20_r;
wire signed [`OutBus]		out_27_20_i;
wire signed [`OutBus]		out_27_21_r;
wire signed [`OutBus]		out_27_21_i;
wire signed [`OutBus]		out_27_22_r;
wire signed [`OutBus]		out_27_22_i;
wire signed [`OutBus]		out_27_23_r;
wire signed [`OutBus]		out_27_23_i;
wire signed [`OutBus]		out_27_24_r;
wire signed [`OutBus]		out_27_24_i;
wire signed [`OutBus]		out_27_25_r;
wire signed [`OutBus]		out_27_25_i;
wire signed [`OutBus]		out_27_26_r;
wire signed [`OutBus]		out_27_26_i;
wire signed [`OutBus]		out_27_27_r;
wire signed [`OutBus]		out_27_27_i;
wire signed [`OutBus]		out_27_28_r;
wire signed [`OutBus]		out_27_28_i;
wire signed [`OutBus]		out_27_29_r;
wire signed [`OutBus]		out_27_29_i;
wire signed [`OutBus]		out_27_30_r;
wire signed [`OutBus]		out_27_30_i;
wire signed [`OutBus]		out_27_31_r;
wire signed [`OutBus]		out_27_31_i;
wire signed [`OutBus]		out_27_32_r;
wire signed [`OutBus]		out_27_32_i;
wire signed [`OutBus]		out_28_1_r;
wire signed [`OutBus]		out_28_1_i;
wire signed [`OutBus]		out_28_2_r;
wire signed [`OutBus]		out_28_2_i;
wire signed [`OutBus]		out_28_3_r;
wire signed [`OutBus]		out_28_3_i;
wire signed [`OutBus]		out_28_4_r;
wire signed [`OutBus]		out_28_4_i;
wire signed [`OutBus]		out_28_5_r;
wire signed [`OutBus]		out_28_5_i;
wire signed [`OutBus]		out_28_6_r;
wire signed [`OutBus]		out_28_6_i;
wire signed [`OutBus]		out_28_7_r;
wire signed [`OutBus]		out_28_7_i;
wire signed [`OutBus]		out_28_8_r;
wire signed [`OutBus]		out_28_8_i;
wire signed [`OutBus]		out_28_9_r;
wire signed [`OutBus]		out_28_9_i;
wire signed [`OutBus]		out_28_10_r;
wire signed [`OutBus]		out_28_10_i;
wire signed [`OutBus]		out_28_11_r;
wire signed [`OutBus]		out_28_11_i;
wire signed [`OutBus]		out_28_12_r;
wire signed [`OutBus]		out_28_12_i;
wire signed [`OutBus]		out_28_13_r;
wire signed [`OutBus]		out_28_13_i;
wire signed [`OutBus]		out_28_14_r;
wire signed [`OutBus]		out_28_14_i;
wire signed [`OutBus]		out_28_15_r;
wire signed [`OutBus]		out_28_15_i;
wire signed [`OutBus]		out_28_16_r;
wire signed [`OutBus]		out_28_16_i;
wire signed [`OutBus]		out_28_17_r;
wire signed [`OutBus]		out_28_17_i;
wire signed [`OutBus]		out_28_18_r;
wire signed [`OutBus]		out_28_18_i;
wire signed [`OutBus]		out_28_19_r;
wire signed [`OutBus]		out_28_19_i;
wire signed [`OutBus]		out_28_20_r;
wire signed [`OutBus]		out_28_20_i;
wire signed [`OutBus]		out_28_21_r;
wire signed [`OutBus]		out_28_21_i;
wire signed [`OutBus]		out_28_22_r;
wire signed [`OutBus]		out_28_22_i;
wire signed [`OutBus]		out_28_23_r;
wire signed [`OutBus]		out_28_23_i;
wire signed [`OutBus]		out_28_24_r;
wire signed [`OutBus]		out_28_24_i;
wire signed [`OutBus]		out_28_25_r;
wire signed [`OutBus]		out_28_25_i;
wire signed [`OutBus]		out_28_26_r;
wire signed [`OutBus]		out_28_26_i;
wire signed [`OutBus]		out_28_27_r;
wire signed [`OutBus]		out_28_27_i;
wire signed [`OutBus]		out_28_28_r;
wire signed [`OutBus]		out_28_28_i;
wire signed [`OutBus]		out_28_29_r;
wire signed [`OutBus]		out_28_29_i;
wire signed [`OutBus]		out_28_30_r;
wire signed [`OutBus]		out_28_30_i;
wire signed [`OutBus]		out_28_31_r;
wire signed [`OutBus]		out_28_31_i;
wire signed [`OutBus]		out_28_32_r;
wire signed [`OutBus]		out_28_32_i;
wire signed [`OutBus]		out_29_1_r;
wire signed [`OutBus]		out_29_1_i;
wire signed [`OutBus]		out_29_2_r;
wire signed [`OutBus]		out_29_2_i;
wire signed [`OutBus]		out_29_3_r;
wire signed [`OutBus]		out_29_3_i;
wire signed [`OutBus]		out_29_4_r;
wire signed [`OutBus]		out_29_4_i;
wire signed [`OutBus]		out_29_5_r;
wire signed [`OutBus]		out_29_5_i;
wire signed [`OutBus]		out_29_6_r;
wire signed [`OutBus]		out_29_6_i;
wire signed [`OutBus]		out_29_7_r;
wire signed [`OutBus]		out_29_7_i;
wire signed [`OutBus]		out_29_8_r;
wire signed [`OutBus]		out_29_8_i;
wire signed [`OutBus]		out_29_9_r;
wire signed [`OutBus]		out_29_9_i;
wire signed [`OutBus]		out_29_10_r;
wire signed [`OutBus]		out_29_10_i;
wire signed [`OutBus]		out_29_11_r;
wire signed [`OutBus]		out_29_11_i;
wire signed [`OutBus]		out_29_12_r;
wire signed [`OutBus]		out_29_12_i;
wire signed [`OutBus]		out_29_13_r;
wire signed [`OutBus]		out_29_13_i;
wire signed [`OutBus]		out_29_14_r;
wire signed [`OutBus]		out_29_14_i;
wire signed [`OutBus]		out_29_15_r;
wire signed [`OutBus]		out_29_15_i;
wire signed [`OutBus]		out_29_16_r;
wire signed [`OutBus]		out_29_16_i;
wire signed [`OutBus]		out_29_17_r;
wire signed [`OutBus]		out_29_17_i;
wire signed [`OutBus]		out_29_18_r;
wire signed [`OutBus]		out_29_18_i;
wire signed [`OutBus]		out_29_19_r;
wire signed [`OutBus]		out_29_19_i;
wire signed [`OutBus]		out_29_20_r;
wire signed [`OutBus]		out_29_20_i;
wire signed [`OutBus]		out_29_21_r;
wire signed [`OutBus]		out_29_21_i;
wire signed [`OutBus]		out_29_22_r;
wire signed [`OutBus]		out_29_22_i;
wire signed [`OutBus]		out_29_23_r;
wire signed [`OutBus]		out_29_23_i;
wire signed [`OutBus]		out_29_24_r;
wire signed [`OutBus]		out_29_24_i;
wire signed [`OutBus]		out_29_25_r;
wire signed [`OutBus]		out_29_25_i;
wire signed [`OutBus]		out_29_26_r;
wire signed [`OutBus]		out_29_26_i;
wire signed [`OutBus]		out_29_27_r;
wire signed [`OutBus]		out_29_27_i;
wire signed [`OutBus]		out_29_28_r;
wire signed [`OutBus]		out_29_28_i;
wire signed [`OutBus]		out_29_29_r;
wire signed [`OutBus]		out_29_29_i;
wire signed [`OutBus]		out_29_30_r;
wire signed [`OutBus]		out_29_30_i;
wire signed [`OutBus]		out_29_31_r;
wire signed [`OutBus]		out_29_31_i;
wire signed [`OutBus]		out_29_32_r;
wire signed [`OutBus]		out_29_32_i;
wire signed [`OutBus]		out_30_1_r;
wire signed [`OutBus]		out_30_1_i;
wire signed [`OutBus]		out_30_2_r;
wire signed [`OutBus]		out_30_2_i;
wire signed [`OutBus]		out_30_3_r;
wire signed [`OutBus]		out_30_3_i;
wire signed [`OutBus]		out_30_4_r;
wire signed [`OutBus]		out_30_4_i;
wire signed [`OutBus]		out_30_5_r;
wire signed [`OutBus]		out_30_5_i;
wire signed [`OutBus]		out_30_6_r;
wire signed [`OutBus]		out_30_6_i;
wire signed [`OutBus]		out_30_7_r;
wire signed [`OutBus]		out_30_7_i;
wire signed [`OutBus]		out_30_8_r;
wire signed [`OutBus]		out_30_8_i;
wire signed [`OutBus]		out_30_9_r;
wire signed [`OutBus]		out_30_9_i;
wire signed [`OutBus]		out_30_10_r;
wire signed [`OutBus]		out_30_10_i;
wire signed [`OutBus]		out_30_11_r;
wire signed [`OutBus]		out_30_11_i;
wire signed [`OutBus]		out_30_12_r;
wire signed [`OutBus]		out_30_12_i;
wire signed [`OutBus]		out_30_13_r;
wire signed [`OutBus]		out_30_13_i;
wire signed [`OutBus]		out_30_14_r;
wire signed [`OutBus]		out_30_14_i;
wire signed [`OutBus]		out_30_15_r;
wire signed [`OutBus]		out_30_15_i;
wire signed [`OutBus]		out_30_16_r;
wire signed [`OutBus]		out_30_16_i;
wire signed [`OutBus]		out_30_17_r;
wire signed [`OutBus]		out_30_17_i;
wire signed [`OutBus]		out_30_18_r;
wire signed [`OutBus]		out_30_18_i;
wire signed [`OutBus]		out_30_19_r;
wire signed [`OutBus]		out_30_19_i;
wire signed [`OutBus]		out_30_20_r;
wire signed [`OutBus]		out_30_20_i;
wire signed [`OutBus]		out_30_21_r;
wire signed [`OutBus]		out_30_21_i;
wire signed [`OutBus]		out_30_22_r;
wire signed [`OutBus]		out_30_22_i;
wire signed [`OutBus]		out_30_23_r;
wire signed [`OutBus]		out_30_23_i;
wire signed [`OutBus]		out_30_24_r;
wire signed [`OutBus]		out_30_24_i;
wire signed [`OutBus]		out_30_25_r;
wire signed [`OutBus]		out_30_25_i;
wire signed [`OutBus]		out_30_26_r;
wire signed [`OutBus]		out_30_26_i;
wire signed [`OutBus]		out_30_27_r;
wire signed [`OutBus]		out_30_27_i;
wire signed [`OutBus]		out_30_28_r;
wire signed [`OutBus]		out_30_28_i;
wire signed [`OutBus]		out_30_29_r;
wire signed [`OutBus]		out_30_29_i;
wire signed [`OutBus]		out_30_30_r;
wire signed [`OutBus]		out_30_30_i;
wire signed [`OutBus]		out_30_31_r;
wire signed [`OutBus]		out_30_31_i;
wire signed [`OutBus]		out_30_32_r;
wire signed [`OutBus]		out_30_32_i;
wire signed [`OutBus]		out_31_1_r;
wire signed [`OutBus]		out_31_1_i;
wire signed [`OutBus]		out_31_2_r;
wire signed [`OutBus]		out_31_2_i;
wire signed [`OutBus]		out_31_3_r;
wire signed [`OutBus]		out_31_3_i;
wire signed [`OutBus]		out_31_4_r;
wire signed [`OutBus]		out_31_4_i;
wire signed [`OutBus]		out_31_5_r;
wire signed [`OutBus]		out_31_5_i;
wire signed [`OutBus]		out_31_6_r;
wire signed [`OutBus]		out_31_6_i;
wire signed [`OutBus]		out_31_7_r;
wire signed [`OutBus]		out_31_7_i;
wire signed [`OutBus]		out_31_8_r;
wire signed [`OutBus]		out_31_8_i;
wire signed [`OutBus]		out_31_9_r;
wire signed [`OutBus]		out_31_9_i;
wire signed [`OutBus]		out_31_10_r;
wire signed [`OutBus]		out_31_10_i;
wire signed [`OutBus]		out_31_11_r;
wire signed [`OutBus]		out_31_11_i;
wire signed [`OutBus]		out_31_12_r;
wire signed [`OutBus]		out_31_12_i;
wire signed [`OutBus]		out_31_13_r;
wire signed [`OutBus]		out_31_13_i;
wire signed [`OutBus]		out_31_14_r;
wire signed [`OutBus]		out_31_14_i;
wire signed [`OutBus]		out_31_15_r;
wire signed [`OutBus]		out_31_15_i;
wire signed [`OutBus]		out_31_16_r;
wire signed [`OutBus]		out_31_16_i;
wire signed [`OutBus]		out_31_17_r;
wire signed [`OutBus]		out_31_17_i;
wire signed [`OutBus]		out_31_18_r;
wire signed [`OutBus]		out_31_18_i;
wire signed [`OutBus]		out_31_19_r;
wire signed [`OutBus]		out_31_19_i;
wire signed [`OutBus]		out_31_20_r;
wire signed [`OutBus]		out_31_20_i;
wire signed [`OutBus]		out_31_21_r;
wire signed [`OutBus]		out_31_21_i;
wire signed [`OutBus]		out_31_22_r;
wire signed [`OutBus]		out_31_22_i;
wire signed [`OutBus]		out_31_23_r;
wire signed [`OutBus]		out_31_23_i;
wire signed [`OutBus]		out_31_24_r;
wire signed [`OutBus]		out_31_24_i;
wire signed [`OutBus]		out_31_25_r;
wire signed [`OutBus]		out_31_25_i;
wire signed [`OutBus]		out_31_26_r;
wire signed [`OutBus]		out_31_26_i;
wire signed [`OutBus]		out_31_27_r;
wire signed [`OutBus]		out_31_27_i;
wire signed [`OutBus]		out_31_28_r;
wire signed [`OutBus]		out_31_28_i;
wire signed [`OutBus]		out_31_29_r;
wire signed [`OutBus]		out_31_29_i;
wire signed [`OutBus]		out_31_30_r;
wire signed [`OutBus]		out_31_30_i;
wire signed [`OutBus]		out_31_31_r;
wire signed [`OutBus]		out_31_31_i;
wire signed [`OutBus]		out_31_32_r;
wire signed [`OutBus]		out_31_32_i;
wire signed [`OutBus]		out_32_1_r;
wire signed [`OutBus]		out_32_1_i;
wire signed [`OutBus]		out_32_2_r;
wire signed [`OutBus]		out_32_2_i;
wire signed [`OutBus]		out_32_3_r;
wire signed [`OutBus]		out_32_3_i;
wire signed [`OutBus]		out_32_4_r;
wire signed [`OutBus]		out_32_4_i;
wire signed [`OutBus]		out_32_5_r;
wire signed [`OutBus]		out_32_5_i;
wire signed [`OutBus]		out_32_6_r;
wire signed [`OutBus]		out_32_6_i;
wire signed [`OutBus]		out_32_7_r;
wire signed [`OutBus]		out_32_7_i;
wire signed [`OutBus]		out_32_8_r;
wire signed [`OutBus]		out_32_8_i;
wire signed [`OutBus]		out_32_9_r;
wire signed [`OutBus]		out_32_9_i;
wire signed [`OutBus]		out_32_10_r;
wire signed [`OutBus]		out_32_10_i;
wire signed [`OutBus]		out_32_11_r;
wire signed [`OutBus]		out_32_11_i;
wire signed [`OutBus]		out_32_12_r;
wire signed [`OutBus]		out_32_12_i;
wire signed [`OutBus]		out_32_13_r;
wire signed [`OutBus]		out_32_13_i;
wire signed [`OutBus]		out_32_14_r;
wire signed [`OutBus]		out_32_14_i;
wire signed [`OutBus]		out_32_15_r;
wire signed [`OutBus]		out_32_15_i;
wire signed [`OutBus]		out_32_16_r;
wire signed [`OutBus]		out_32_16_i;
wire signed [`OutBus]		out_32_17_r;
wire signed [`OutBus]		out_32_17_i;
wire signed [`OutBus]		out_32_18_r;
wire signed [`OutBus]		out_32_18_i;
wire signed [`OutBus]		out_32_19_r;
wire signed [`OutBus]		out_32_19_i;
wire signed [`OutBus]		out_32_20_r;
wire signed [`OutBus]		out_32_20_i;
wire signed [`OutBus]		out_32_21_r;
wire signed [`OutBus]		out_32_21_i;
wire signed [`OutBus]		out_32_22_r;
wire signed [`OutBus]		out_32_22_i;
wire signed [`OutBus]		out_32_23_r;
wire signed [`OutBus]		out_32_23_i;
wire signed [`OutBus]		out_32_24_r;
wire signed [`OutBus]		out_32_24_i;
wire signed [`OutBus]		out_32_25_r;
wire signed [`OutBus]		out_32_25_i;
wire signed [`OutBus]		out_32_26_r;
wire signed [`OutBus]		out_32_26_i;
wire signed [`OutBus]		out_32_27_r;
wire signed [`OutBus]		out_32_27_i;
wire signed [`OutBus]		out_32_28_r;
wire signed [`OutBus]		out_32_28_i;
wire signed [`OutBus]		out_32_29_r;
wire signed [`OutBus]		out_32_29_i;
wire signed [`OutBus]		out_32_30_r;
wire signed [`OutBus]		out_32_30_i;
wire signed [`OutBus]		out_32_31_r;
wire signed [`OutBus]		out_32_31_i;
wire signed [`OutBus]		out_32_32_r;
wire signed [`OutBus]		out_32_32_i;

top sim (clk,in_1_1_r,in_1_1_i,in_1_2_r,in_1_2_i,in_1_3_r,in_1_3_i,in_1_4_r,in_1_4_i,in_1_5_r,in_1_5_i,in_1_6_r,in_1_6_i,in_1_7_r,in_1_7_i,in_1_8_r,in_1_8_i,in_1_9_r,in_1_9_i,in_1_10_r,in_1_10_i,in_1_11_r,in_1_11_i,in_1_12_r,in_1_12_i,in_1_13_r,in_1_13_i,in_1_14_r,in_1_14_i,in_1_15_r,in_1_15_i,in_1_16_r,in_1_16_i,in_1_17_r,in_1_17_i,in_1_18_r,in_1_18_i,in_1_19_r,in_1_19_i,in_1_20_r,in_1_20_i,in_1_21_r,in_1_21_i,in_1_22_r,in_1_22_i,in_1_23_r,in_1_23_i,in_1_24_r,in_1_24_i,in_1_25_r,in_1_25_i,in_1_26_r,in_1_26_i,in_1_27_r,in_1_27_i,in_1_28_r,in_1_28_i,in_1_29_r,in_1_29_i,in_1_30_r,in_1_30_i,in_1_31_r,in_1_31_i,in_1_32_r,in_1_32_i,in_2_1_r,in_2_1_i,in_2_2_r,in_2_2_i,in_2_3_r,in_2_3_i,in_2_4_r,in_2_4_i,in_2_5_r,in_2_5_i,in_2_6_r,in_2_6_i,in_2_7_r,in_2_7_i,in_2_8_r,in_2_8_i,in_2_9_r,in_2_9_i,in_2_10_r,in_2_10_i,in_2_11_r,in_2_11_i,in_2_12_r,in_2_12_i,in_2_13_r,in_2_13_i,in_2_14_r,in_2_14_i,in_2_15_r,in_2_15_i,in_2_16_r,in_2_16_i,in_2_17_r,in_2_17_i,in_2_18_r,in_2_18_i,in_2_19_r,in_2_19_i,in_2_20_r,in_2_20_i,in_2_21_r,in_2_21_i,in_2_22_r,in_2_22_i,in_2_23_r,in_2_23_i,in_2_24_r,in_2_24_i,in_2_25_r,in_2_25_i,in_2_26_r,in_2_26_i,in_2_27_r,in_2_27_i,in_2_28_r,in_2_28_i,in_2_29_r,in_2_29_i,in_2_30_r,in_2_30_i,in_2_31_r,in_2_31_i,in_2_32_r,in_2_32_i,in_3_1_r,in_3_1_i,in_3_2_r,in_3_2_i,in_3_3_r,in_3_3_i,in_3_4_r,in_3_4_i,in_3_5_r,in_3_5_i,in_3_6_r,in_3_6_i,in_3_7_r,in_3_7_i,in_3_8_r,in_3_8_i,in_3_9_r,in_3_9_i,in_3_10_r,in_3_10_i,in_3_11_r,in_3_11_i,in_3_12_r,in_3_12_i,in_3_13_r,in_3_13_i,in_3_14_r,in_3_14_i,in_3_15_r,in_3_15_i,in_3_16_r,in_3_16_i,in_3_17_r,in_3_17_i,in_3_18_r,in_3_18_i,in_3_19_r,in_3_19_i,in_3_20_r,in_3_20_i,in_3_21_r,in_3_21_i,in_3_22_r,in_3_22_i,in_3_23_r,in_3_23_i,in_3_24_r,in_3_24_i,in_3_25_r,in_3_25_i,in_3_26_r,in_3_26_i,in_3_27_r,in_3_27_i,in_3_28_r,in_3_28_i,in_3_29_r,in_3_29_i,in_3_30_r,in_3_30_i,in_3_31_r,in_3_31_i,in_3_32_r,in_3_32_i,in_4_1_r,in_4_1_i,in_4_2_r,in_4_2_i,in_4_3_r,in_4_3_i,in_4_4_r,in_4_4_i,in_4_5_r,in_4_5_i,in_4_6_r,in_4_6_i,in_4_7_r,in_4_7_i,in_4_8_r,in_4_8_i,in_4_9_r,in_4_9_i,in_4_10_r,in_4_10_i,in_4_11_r,in_4_11_i,in_4_12_r,in_4_12_i,in_4_13_r,in_4_13_i,in_4_14_r,in_4_14_i,in_4_15_r,in_4_15_i,in_4_16_r,in_4_16_i,in_4_17_r,in_4_17_i,in_4_18_r,in_4_18_i,in_4_19_r,in_4_19_i,in_4_20_r,in_4_20_i,in_4_21_r,in_4_21_i,in_4_22_r,in_4_22_i,in_4_23_r,in_4_23_i,in_4_24_r,in_4_24_i,in_4_25_r,in_4_25_i,in_4_26_r,in_4_26_i,in_4_27_r,in_4_27_i,in_4_28_r,in_4_28_i,in_4_29_r,in_4_29_i,in_4_30_r,in_4_30_i,in_4_31_r,in_4_31_i,in_4_32_r,in_4_32_i,in_5_1_r,in_5_1_i,in_5_2_r,in_5_2_i,in_5_3_r,in_5_3_i,in_5_4_r,in_5_4_i,in_5_5_r,in_5_5_i,in_5_6_r,in_5_6_i,in_5_7_r,in_5_7_i,in_5_8_r,in_5_8_i,in_5_9_r,in_5_9_i,in_5_10_r,in_5_10_i,in_5_11_r,in_5_11_i,in_5_12_r,in_5_12_i,in_5_13_r,in_5_13_i,in_5_14_r,in_5_14_i,in_5_15_r,in_5_15_i,in_5_16_r,in_5_16_i,in_5_17_r,in_5_17_i,in_5_18_r,in_5_18_i,in_5_19_r,in_5_19_i,in_5_20_r,in_5_20_i,in_5_21_r,in_5_21_i,in_5_22_r,in_5_22_i,in_5_23_r,in_5_23_i,in_5_24_r,in_5_24_i,in_5_25_r,in_5_25_i,in_5_26_r,in_5_26_i,in_5_27_r,in_5_27_i,in_5_28_r,in_5_28_i,in_5_29_r,in_5_29_i,in_5_30_r,in_5_30_i,in_5_31_r,in_5_31_i,in_5_32_r,in_5_32_i,in_6_1_r,in_6_1_i,in_6_2_r,in_6_2_i,in_6_3_r,in_6_3_i,in_6_4_r,in_6_4_i,in_6_5_r,in_6_5_i,in_6_6_r,in_6_6_i,in_6_7_r,in_6_7_i,in_6_8_r,in_6_8_i,in_6_9_r,in_6_9_i,in_6_10_r,in_6_10_i,in_6_11_r,in_6_11_i,in_6_12_r,in_6_12_i,in_6_13_r,in_6_13_i,in_6_14_r,in_6_14_i,in_6_15_r,in_6_15_i,in_6_16_r,in_6_16_i,in_6_17_r,in_6_17_i,in_6_18_r,in_6_18_i,in_6_19_r,in_6_19_i,in_6_20_r,in_6_20_i,in_6_21_r,in_6_21_i,in_6_22_r,in_6_22_i,in_6_23_r,in_6_23_i,in_6_24_r,in_6_24_i,in_6_25_r,in_6_25_i,in_6_26_r,in_6_26_i,in_6_27_r,in_6_27_i,in_6_28_r,in_6_28_i,in_6_29_r,in_6_29_i,in_6_30_r,in_6_30_i,in_6_31_r,in_6_31_i,in_6_32_r,in_6_32_i,in_7_1_r,in_7_1_i,in_7_2_r,in_7_2_i,in_7_3_r,in_7_3_i,in_7_4_r,in_7_4_i,in_7_5_r,in_7_5_i,in_7_6_r,in_7_6_i,in_7_7_r,in_7_7_i,in_7_8_r,in_7_8_i,in_7_9_r,in_7_9_i,in_7_10_r,in_7_10_i,in_7_11_r,in_7_11_i,in_7_12_r,in_7_12_i,in_7_13_r,in_7_13_i,in_7_14_r,in_7_14_i,in_7_15_r,in_7_15_i,in_7_16_r,in_7_16_i,in_7_17_r,in_7_17_i,in_7_18_r,in_7_18_i,in_7_19_r,in_7_19_i,in_7_20_r,in_7_20_i,in_7_21_r,in_7_21_i,in_7_22_r,in_7_22_i,in_7_23_r,in_7_23_i,in_7_24_r,in_7_24_i,in_7_25_r,in_7_25_i,in_7_26_r,in_7_26_i,in_7_27_r,in_7_27_i,in_7_28_r,in_7_28_i,in_7_29_r,in_7_29_i,in_7_30_r,in_7_30_i,in_7_31_r,in_7_31_i,in_7_32_r,in_7_32_i,in_8_1_r,in_8_1_i,in_8_2_r,in_8_2_i,in_8_3_r,in_8_3_i,in_8_4_r,in_8_4_i,in_8_5_r,in_8_5_i,in_8_6_r,in_8_6_i,in_8_7_r,in_8_7_i,in_8_8_r,in_8_8_i,in_8_9_r,in_8_9_i,in_8_10_r,in_8_10_i,in_8_11_r,in_8_11_i,in_8_12_r,in_8_12_i,in_8_13_r,in_8_13_i,in_8_14_r,in_8_14_i,in_8_15_r,in_8_15_i,in_8_16_r,in_8_16_i,in_8_17_r,in_8_17_i,in_8_18_r,in_8_18_i,in_8_19_r,in_8_19_i,in_8_20_r,in_8_20_i,in_8_21_r,in_8_21_i,in_8_22_r,in_8_22_i,in_8_23_r,in_8_23_i,in_8_24_r,in_8_24_i,in_8_25_r,in_8_25_i,in_8_26_r,in_8_26_i,in_8_27_r,in_8_27_i,in_8_28_r,in_8_28_i,in_8_29_r,in_8_29_i,in_8_30_r,in_8_30_i,in_8_31_r,in_8_31_i,in_8_32_r,in_8_32_i,in_9_1_r,in_9_1_i,in_9_2_r,in_9_2_i,in_9_3_r,in_9_3_i,in_9_4_r,in_9_4_i,in_9_5_r,in_9_5_i,in_9_6_r,in_9_6_i,in_9_7_r,in_9_7_i,in_9_8_r,in_9_8_i,in_9_9_r,in_9_9_i,in_9_10_r,in_9_10_i,in_9_11_r,in_9_11_i,in_9_12_r,in_9_12_i,in_9_13_r,in_9_13_i,in_9_14_r,in_9_14_i,in_9_15_r,in_9_15_i,in_9_16_r,in_9_16_i,in_9_17_r,in_9_17_i,in_9_18_r,in_9_18_i,in_9_19_r,in_9_19_i,in_9_20_r,in_9_20_i,in_9_21_r,in_9_21_i,in_9_22_r,in_9_22_i,in_9_23_r,in_9_23_i,in_9_24_r,in_9_24_i,in_9_25_r,in_9_25_i,in_9_26_r,in_9_26_i,in_9_27_r,in_9_27_i,in_9_28_r,in_9_28_i,in_9_29_r,in_9_29_i,in_9_30_r,in_9_30_i,in_9_31_r,in_9_31_i,in_9_32_r,in_9_32_i,in_10_1_r,in_10_1_i,in_10_2_r,in_10_2_i,in_10_3_r,in_10_3_i,in_10_4_r,in_10_4_i,in_10_5_r,in_10_5_i,in_10_6_r,in_10_6_i,in_10_7_r,in_10_7_i,in_10_8_r,in_10_8_i,in_10_9_r,in_10_9_i,in_10_10_r,in_10_10_i,in_10_11_r,in_10_11_i,in_10_12_r,in_10_12_i,in_10_13_r,in_10_13_i,in_10_14_r,in_10_14_i,in_10_15_r,in_10_15_i,in_10_16_r,in_10_16_i,in_10_17_r,in_10_17_i,in_10_18_r,in_10_18_i,in_10_19_r,in_10_19_i,in_10_20_r,in_10_20_i,in_10_21_r,in_10_21_i,in_10_22_r,in_10_22_i,in_10_23_r,in_10_23_i,in_10_24_r,in_10_24_i,in_10_25_r,in_10_25_i,in_10_26_r,in_10_26_i,in_10_27_r,in_10_27_i,in_10_28_r,in_10_28_i,in_10_29_r,in_10_29_i,in_10_30_r,in_10_30_i,in_10_31_r,in_10_31_i,in_10_32_r,in_10_32_i,in_11_1_r,in_11_1_i,in_11_2_r,in_11_2_i,in_11_3_r,in_11_3_i,in_11_4_r,in_11_4_i,in_11_5_r,in_11_5_i,in_11_6_r,in_11_6_i,in_11_7_r,in_11_7_i,in_11_8_r,in_11_8_i,in_11_9_r,in_11_9_i,in_11_10_r,in_11_10_i,in_11_11_r,in_11_11_i,in_11_12_r,in_11_12_i,in_11_13_r,in_11_13_i,in_11_14_r,in_11_14_i,in_11_15_r,in_11_15_i,in_11_16_r,in_11_16_i,in_11_17_r,in_11_17_i,in_11_18_r,in_11_18_i,in_11_19_r,in_11_19_i,in_11_20_r,in_11_20_i,in_11_21_r,in_11_21_i,in_11_22_r,in_11_22_i,in_11_23_r,in_11_23_i,in_11_24_r,in_11_24_i,in_11_25_r,in_11_25_i,in_11_26_r,in_11_26_i,in_11_27_r,in_11_27_i,in_11_28_r,in_11_28_i,in_11_29_r,in_11_29_i,in_11_30_r,in_11_30_i,in_11_31_r,in_11_31_i,in_11_32_r,in_11_32_i,in_12_1_r,in_12_1_i,in_12_2_r,in_12_2_i,in_12_3_r,in_12_3_i,in_12_4_r,in_12_4_i,in_12_5_r,in_12_5_i,in_12_6_r,in_12_6_i,in_12_7_r,in_12_7_i,in_12_8_r,in_12_8_i,in_12_9_r,in_12_9_i,in_12_10_r,in_12_10_i,in_12_11_r,in_12_11_i,in_12_12_r,in_12_12_i,in_12_13_r,in_12_13_i,in_12_14_r,in_12_14_i,in_12_15_r,in_12_15_i,in_12_16_r,in_12_16_i,in_12_17_r,in_12_17_i,in_12_18_r,in_12_18_i,in_12_19_r,in_12_19_i,in_12_20_r,in_12_20_i,in_12_21_r,in_12_21_i,in_12_22_r,in_12_22_i,in_12_23_r,in_12_23_i,in_12_24_r,in_12_24_i,in_12_25_r,in_12_25_i,in_12_26_r,in_12_26_i,in_12_27_r,in_12_27_i,in_12_28_r,in_12_28_i,in_12_29_r,in_12_29_i,in_12_30_r,in_12_30_i,in_12_31_r,in_12_31_i,in_12_32_r,in_12_32_i,in_13_1_r,in_13_1_i,in_13_2_r,in_13_2_i,in_13_3_r,in_13_3_i,in_13_4_r,in_13_4_i,in_13_5_r,in_13_5_i,in_13_6_r,in_13_6_i,in_13_7_r,in_13_7_i,in_13_8_r,in_13_8_i,in_13_9_r,in_13_9_i,in_13_10_r,in_13_10_i,in_13_11_r,in_13_11_i,in_13_12_r,in_13_12_i,in_13_13_r,in_13_13_i,in_13_14_r,in_13_14_i,in_13_15_r,in_13_15_i,in_13_16_r,in_13_16_i,in_13_17_r,in_13_17_i,in_13_18_r,in_13_18_i,in_13_19_r,in_13_19_i,in_13_20_r,in_13_20_i,in_13_21_r,in_13_21_i,in_13_22_r,in_13_22_i,in_13_23_r,in_13_23_i,in_13_24_r,in_13_24_i,in_13_25_r,in_13_25_i,in_13_26_r,in_13_26_i,in_13_27_r,in_13_27_i,in_13_28_r,in_13_28_i,in_13_29_r,in_13_29_i,in_13_30_r,in_13_30_i,in_13_31_r,in_13_31_i,in_13_32_r,in_13_32_i,in_14_1_r,in_14_1_i,in_14_2_r,in_14_2_i,in_14_3_r,in_14_3_i,in_14_4_r,in_14_4_i,in_14_5_r,in_14_5_i,in_14_6_r,in_14_6_i,in_14_7_r,in_14_7_i,in_14_8_r,in_14_8_i,in_14_9_r,in_14_9_i,in_14_10_r,in_14_10_i,in_14_11_r,in_14_11_i,in_14_12_r,in_14_12_i,in_14_13_r,in_14_13_i,in_14_14_r,in_14_14_i,in_14_15_r,in_14_15_i,in_14_16_r,in_14_16_i,in_14_17_r,in_14_17_i,in_14_18_r,in_14_18_i,in_14_19_r,in_14_19_i,in_14_20_r,in_14_20_i,in_14_21_r,in_14_21_i,in_14_22_r,in_14_22_i,in_14_23_r,in_14_23_i,in_14_24_r,in_14_24_i,in_14_25_r,in_14_25_i,in_14_26_r,in_14_26_i,in_14_27_r,in_14_27_i,in_14_28_r,in_14_28_i,in_14_29_r,in_14_29_i,in_14_30_r,in_14_30_i,in_14_31_r,in_14_31_i,in_14_32_r,in_14_32_i,in_15_1_r,in_15_1_i,in_15_2_r,in_15_2_i,in_15_3_r,in_15_3_i,in_15_4_r,in_15_4_i,in_15_5_r,in_15_5_i,in_15_6_r,in_15_6_i,in_15_7_r,in_15_7_i,in_15_8_r,in_15_8_i,in_15_9_r,in_15_9_i,in_15_10_r,in_15_10_i,in_15_11_r,in_15_11_i,in_15_12_r,in_15_12_i,in_15_13_r,in_15_13_i,in_15_14_r,in_15_14_i,in_15_15_r,in_15_15_i,in_15_16_r,in_15_16_i,in_15_17_r,in_15_17_i,in_15_18_r,in_15_18_i,in_15_19_r,in_15_19_i,in_15_20_r,in_15_20_i,in_15_21_r,in_15_21_i,in_15_22_r,in_15_22_i,in_15_23_r,in_15_23_i,in_15_24_r,in_15_24_i,in_15_25_r,in_15_25_i,in_15_26_r,in_15_26_i,in_15_27_r,in_15_27_i,in_15_28_r,in_15_28_i,in_15_29_r,in_15_29_i,in_15_30_r,in_15_30_i,in_15_31_r,in_15_31_i,in_15_32_r,in_15_32_i,in_16_1_r,in_16_1_i,in_16_2_r,in_16_2_i,in_16_3_r,in_16_3_i,in_16_4_r,in_16_4_i,in_16_5_r,in_16_5_i,in_16_6_r,in_16_6_i,in_16_7_r,in_16_7_i,in_16_8_r,in_16_8_i,in_16_9_r,in_16_9_i,in_16_10_r,in_16_10_i,in_16_11_r,in_16_11_i,in_16_12_r,in_16_12_i,in_16_13_r,in_16_13_i,in_16_14_r,in_16_14_i,in_16_15_r,in_16_15_i,in_16_16_r,in_16_16_i,in_16_17_r,in_16_17_i,in_16_18_r,in_16_18_i,in_16_19_r,in_16_19_i,in_16_20_r,in_16_20_i,in_16_21_r,in_16_21_i,in_16_22_r,in_16_22_i,in_16_23_r,in_16_23_i,in_16_24_r,in_16_24_i,in_16_25_r,in_16_25_i,in_16_26_r,in_16_26_i,in_16_27_r,in_16_27_i,in_16_28_r,in_16_28_i,in_16_29_r,in_16_29_i,in_16_30_r,in_16_30_i,in_16_31_r,in_16_31_i,in_16_32_r,in_16_32_i,in_17_1_r,in_17_1_i,in_17_2_r,in_17_2_i,in_17_3_r,in_17_3_i,in_17_4_r,in_17_4_i,in_17_5_r,in_17_5_i,in_17_6_r,in_17_6_i,in_17_7_r,in_17_7_i,in_17_8_r,in_17_8_i,in_17_9_r,in_17_9_i,in_17_10_r,in_17_10_i,in_17_11_r,in_17_11_i,in_17_12_r,in_17_12_i,in_17_13_r,in_17_13_i,in_17_14_r,in_17_14_i,in_17_15_r,in_17_15_i,in_17_16_r,in_17_16_i,in_17_17_r,in_17_17_i,in_17_18_r,in_17_18_i,in_17_19_r,in_17_19_i,in_17_20_r,in_17_20_i,in_17_21_r,in_17_21_i,in_17_22_r,in_17_22_i,in_17_23_r,in_17_23_i,in_17_24_r,in_17_24_i,in_17_25_r,in_17_25_i,in_17_26_r,in_17_26_i,in_17_27_r,in_17_27_i,in_17_28_r,in_17_28_i,in_17_29_r,in_17_29_i,in_17_30_r,in_17_30_i,in_17_31_r,in_17_31_i,in_17_32_r,in_17_32_i,in_18_1_r,in_18_1_i,in_18_2_r,in_18_2_i,in_18_3_r,in_18_3_i,in_18_4_r,in_18_4_i,in_18_5_r,in_18_5_i,in_18_6_r,in_18_6_i,in_18_7_r,in_18_7_i,in_18_8_r,in_18_8_i,in_18_9_r,in_18_9_i,in_18_10_r,in_18_10_i,in_18_11_r,in_18_11_i,in_18_12_r,in_18_12_i,in_18_13_r,in_18_13_i,in_18_14_r,in_18_14_i,in_18_15_r,in_18_15_i,in_18_16_r,in_18_16_i,in_18_17_r,in_18_17_i,in_18_18_r,in_18_18_i,in_18_19_r,in_18_19_i,in_18_20_r,in_18_20_i,in_18_21_r,in_18_21_i,in_18_22_r,in_18_22_i,in_18_23_r,in_18_23_i,in_18_24_r,in_18_24_i,in_18_25_r,in_18_25_i,in_18_26_r,in_18_26_i,in_18_27_r,in_18_27_i,in_18_28_r,in_18_28_i,in_18_29_r,in_18_29_i,in_18_30_r,in_18_30_i,in_18_31_r,in_18_31_i,in_18_32_r,in_18_32_i,in_19_1_r,in_19_1_i,in_19_2_r,in_19_2_i,in_19_3_r,in_19_3_i,in_19_4_r,in_19_4_i,in_19_5_r,in_19_5_i,in_19_6_r,in_19_6_i,in_19_7_r,in_19_7_i,in_19_8_r,in_19_8_i,in_19_9_r,in_19_9_i,in_19_10_r,in_19_10_i,in_19_11_r,in_19_11_i,in_19_12_r,in_19_12_i,in_19_13_r,in_19_13_i,in_19_14_r,in_19_14_i,in_19_15_r,in_19_15_i,in_19_16_r,in_19_16_i,in_19_17_r,in_19_17_i,in_19_18_r,in_19_18_i,in_19_19_r,in_19_19_i,in_19_20_r,in_19_20_i,in_19_21_r,in_19_21_i,in_19_22_r,in_19_22_i,in_19_23_r,in_19_23_i,in_19_24_r,in_19_24_i,in_19_25_r,in_19_25_i,in_19_26_r,in_19_26_i,in_19_27_r,in_19_27_i,in_19_28_r,in_19_28_i,in_19_29_r,in_19_29_i,in_19_30_r,in_19_30_i,in_19_31_r,in_19_31_i,in_19_32_r,in_19_32_i,in_20_1_r,in_20_1_i,in_20_2_r,in_20_2_i,in_20_3_r,in_20_3_i,in_20_4_r,in_20_4_i,in_20_5_r,in_20_5_i,in_20_6_r,in_20_6_i,in_20_7_r,in_20_7_i,in_20_8_r,in_20_8_i,in_20_9_r,in_20_9_i,in_20_10_r,in_20_10_i,in_20_11_r,in_20_11_i,in_20_12_r,in_20_12_i,in_20_13_r,in_20_13_i,in_20_14_r,in_20_14_i,in_20_15_r,in_20_15_i,in_20_16_r,in_20_16_i,in_20_17_r,in_20_17_i,in_20_18_r,in_20_18_i,in_20_19_r,in_20_19_i,in_20_20_r,in_20_20_i,in_20_21_r,in_20_21_i,in_20_22_r,in_20_22_i,in_20_23_r,in_20_23_i,in_20_24_r,in_20_24_i,in_20_25_r,in_20_25_i,in_20_26_r,in_20_26_i,in_20_27_r,in_20_27_i,in_20_28_r,in_20_28_i,in_20_29_r,in_20_29_i,in_20_30_r,in_20_30_i,in_20_31_r,in_20_31_i,in_20_32_r,in_20_32_i,in_21_1_r,in_21_1_i,in_21_2_r,in_21_2_i,in_21_3_r,in_21_3_i,in_21_4_r,in_21_4_i,in_21_5_r,in_21_5_i,in_21_6_r,in_21_6_i,in_21_7_r,in_21_7_i,in_21_8_r,in_21_8_i,in_21_9_r,in_21_9_i,in_21_10_r,in_21_10_i,in_21_11_r,in_21_11_i,in_21_12_r,in_21_12_i,in_21_13_r,in_21_13_i,in_21_14_r,in_21_14_i,in_21_15_r,in_21_15_i,in_21_16_r,in_21_16_i,in_21_17_r,in_21_17_i,in_21_18_r,in_21_18_i,in_21_19_r,in_21_19_i,in_21_20_r,in_21_20_i,in_21_21_r,in_21_21_i,in_21_22_r,in_21_22_i,in_21_23_r,in_21_23_i,in_21_24_r,in_21_24_i,in_21_25_r,in_21_25_i,in_21_26_r,in_21_26_i,in_21_27_r,in_21_27_i,in_21_28_r,in_21_28_i,in_21_29_r,in_21_29_i,in_21_30_r,in_21_30_i,in_21_31_r,in_21_31_i,in_21_32_r,in_21_32_i,in_22_1_r,in_22_1_i,in_22_2_r,in_22_2_i,in_22_3_r,in_22_3_i,in_22_4_r,in_22_4_i,in_22_5_r,in_22_5_i,in_22_6_r,in_22_6_i,in_22_7_r,in_22_7_i,in_22_8_r,in_22_8_i,in_22_9_r,in_22_9_i,in_22_10_r,in_22_10_i,in_22_11_r,in_22_11_i,in_22_12_r,in_22_12_i,in_22_13_r,in_22_13_i,in_22_14_r,in_22_14_i,in_22_15_r,in_22_15_i,in_22_16_r,in_22_16_i,in_22_17_r,in_22_17_i,in_22_18_r,in_22_18_i,in_22_19_r,in_22_19_i,in_22_20_r,in_22_20_i,in_22_21_r,in_22_21_i,in_22_22_r,in_22_22_i,in_22_23_r,in_22_23_i,in_22_24_r,in_22_24_i,in_22_25_r,in_22_25_i,in_22_26_r,in_22_26_i,in_22_27_r,in_22_27_i,in_22_28_r,in_22_28_i,in_22_29_r,in_22_29_i,in_22_30_r,in_22_30_i,in_22_31_r,in_22_31_i,in_22_32_r,in_22_32_i,in_23_1_r,in_23_1_i,in_23_2_r,in_23_2_i,in_23_3_r,in_23_3_i,in_23_4_r,in_23_4_i,in_23_5_r,in_23_5_i,in_23_6_r,in_23_6_i,in_23_7_r,in_23_7_i,in_23_8_r,in_23_8_i,in_23_9_r,in_23_9_i,in_23_10_r,in_23_10_i,in_23_11_r,in_23_11_i,in_23_12_r,in_23_12_i,in_23_13_r,in_23_13_i,in_23_14_r,in_23_14_i,in_23_15_r,in_23_15_i,in_23_16_r,in_23_16_i,in_23_17_r,in_23_17_i,in_23_18_r,in_23_18_i,in_23_19_r,in_23_19_i,in_23_20_r,in_23_20_i,in_23_21_r,in_23_21_i,in_23_22_r,in_23_22_i,in_23_23_r,in_23_23_i,in_23_24_r,in_23_24_i,in_23_25_r,in_23_25_i,in_23_26_r,in_23_26_i,in_23_27_r,in_23_27_i,in_23_28_r,in_23_28_i,in_23_29_r,in_23_29_i,in_23_30_r,in_23_30_i,in_23_31_r,in_23_31_i,in_23_32_r,in_23_32_i,in_24_1_r,in_24_1_i,in_24_2_r,in_24_2_i,in_24_3_r,in_24_3_i,in_24_4_r,in_24_4_i,in_24_5_r,in_24_5_i,in_24_6_r,in_24_6_i,in_24_7_r,in_24_7_i,in_24_8_r,in_24_8_i,in_24_9_r,in_24_9_i,in_24_10_r,in_24_10_i,in_24_11_r,in_24_11_i,in_24_12_r,in_24_12_i,in_24_13_r,in_24_13_i,in_24_14_r,in_24_14_i,in_24_15_r,in_24_15_i,in_24_16_r,in_24_16_i,in_24_17_r,in_24_17_i,in_24_18_r,in_24_18_i,in_24_19_r,in_24_19_i,in_24_20_r,in_24_20_i,in_24_21_r,in_24_21_i,in_24_22_r,in_24_22_i,in_24_23_r,in_24_23_i,in_24_24_r,in_24_24_i,in_24_25_r,in_24_25_i,in_24_26_r,in_24_26_i,in_24_27_r,in_24_27_i,in_24_28_r,in_24_28_i,in_24_29_r,in_24_29_i,in_24_30_r,in_24_30_i,in_24_31_r,in_24_31_i,in_24_32_r,in_24_32_i,in_25_1_r,in_25_1_i,in_25_2_r,in_25_2_i,in_25_3_r,in_25_3_i,in_25_4_r,in_25_4_i,in_25_5_r,in_25_5_i,in_25_6_r,in_25_6_i,in_25_7_r,in_25_7_i,in_25_8_r,in_25_8_i,in_25_9_r,in_25_9_i,in_25_10_r,in_25_10_i,in_25_11_r,in_25_11_i,in_25_12_r,in_25_12_i,in_25_13_r,in_25_13_i,in_25_14_r,in_25_14_i,in_25_15_r,in_25_15_i,in_25_16_r,in_25_16_i,in_25_17_r,in_25_17_i,in_25_18_r,in_25_18_i,in_25_19_r,in_25_19_i,in_25_20_r,in_25_20_i,in_25_21_r,in_25_21_i,in_25_22_r,in_25_22_i,in_25_23_r,in_25_23_i,in_25_24_r,in_25_24_i,in_25_25_r,in_25_25_i,in_25_26_r,in_25_26_i,in_25_27_r,in_25_27_i,in_25_28_r,in_25_28_i,in_25_29_r,in_25_29_i,in_25_30_r,in_25_30_i,in_25_31_r,in_25_31_i,in_25_32_r,in_25_32_i,in_26_1_r,in_26_1_i,in_26_2_r,in_26_2_i,in_26_3_r,in_26_3_i,in_26_4_r,in_26_4_i,in_26_5_r,in_26_5_i,in_26_6_r,in_26_6_i,in_26_7_r,in_26_7_i,in_26_8_r,in_26_8_i,in_26_9_r,in_26_9_i,in_26_10_r,in_26_10_i,in_26_11_r,in_26_11_i,in_26_12_r,in_26_12_i,in_26_13_r,in_26_13_i,in_26_14_r,in_26_14_i,in_26_15_r,in_26_15_i,in_26_16_r,in_26_16_i,in_26_17_r,in_26_17_i,in_26_18_r,in_26_18_i,in_26_19_r,in_26_19_i,in_26_20_r,in_26_20_i,in_26_21_r,in_26_21_i,in_26_22_r,in_26_22_i,in_26_23_r,in_26_23_i,in_26_24_r,in_26_24_i,in_26_25_r,in_26_25_i,in_26_26_r,in_26_26_i,in_26_27_r,in_26_27_i,in_26_28_r,in_26_28_i,in_26_29_r,in_26_29_i,in_26_30_r,in_26_30_i,in_26_31_r,in_26_31_i,in_26_32_r,in_26_32_i,in_27_1_r,in_27_1_i,in_27_2_r,in_27_2_i,in_27_3_r,in_27_3_i,in_27_4_r,in_27_4_i,in_27_5_r,in_27_5_i,in_27_6_r,in_27_6_i,in_27_7_r,in_27_7_i,in_27_8_r,in_27_8_i,in_27_9_r,in_27_9_i,in_27_10_r,in_27_10_i,in_27_11_r,in_27_11_i,in_27_12_r,in_27_12_i,in_27_13_r,in_27_13_i,in_27_14_r,in_27_14_i,in_27_15_r,in_27_15_i,in_27_16_r,in_27_16_i,in_27_17_r,in_27_17_i,in_27_18_r,in_27_18_i,in_27_19_r,in_27_19_i,in_27_20_r,in_27_20_i,in_27_21_r,in_27_21_i,in_27_22_r,in_27_22_i,in_27_23_r,in_27_23_i,in_27_24_r,in_27_24_i,in_27_25_r,in_27_25_i,in_27_26_r,in_27_26_i,in_27_27_r,in_27_27_i,in_27_28_r,in_27_28_i,in_27_29_r,in_27_29_i,in_27_30_r,in_27_30_i,in_27_31_r,in_27_31_i,in_27_32_r,in_27_32_i,in_28_1_r,in_28_1_i,in_28_2_r,in_28_2_i,in_28_3_r,in_28_3_i,in_28_4_r,in_28_4_i,in_28_5_r,in_28_5_i,in_28_6_r,in_28_6_i,in_28_7_r,in_28_7_i,in_28_8_r,in_28_8_i,in_28_9_r,in_28_9_i,in_28_10_r,in_28_10_i,in_28_11_r,in_28_11_i,in_28_12_r,in_28_12_i,in_28_13_r,in_28_13_i,in_28_14_r,in_28_14_i,in_28_15_r,in_28_15_i,in_28_16_r,in_28_16_i,in_28_17_r,in_28_17_i,in_28_18_r,in_28_18_i,in_28_19_r,in_28_19_i,in_28_20_r,in_28_20_i,in_28_21_r,in_28_21_i,in_28_22_r,in_28_22_i,in_28_23_r,in_28_23_i,in_28_24_r,in_28_24_i,in_28_25_r,in_28_25_i,in_28_26_r,in_28_26_i,in_28_27_r,in_28_27_i,in_28_28_r,in_28_28_i,in_28_29_r,in_28_29_i,in_28_30_r,in_28_30_i,in_28_31_r,in_28_31_i,in_28_32_r,in_28_32_i,in_29_1_r,in_29_1_i,in_29_2_r,in_29_2_i,in_29_3_r,in_29_3_i,in_29_4_r,in_29_4_i,in_29_5_r,in_29_5_i,in_29_6_r,in_29_6_i,in_29_7_r,in_29_7_i,in_29_8_r,in_29_8_i,in_29_9_r,in_29_9_i,in_29_10_r,in_29_10_i,in_29_11_r,in_29_11_i,in_29_12_r,in_29_12_i,in_29_13_r,in_29_13_i,in_29_14_r,in_29_14_i,in_29_15_r,in_29_15_i,in_29_16_r,in_29_16_i,in_29_17_r,in_29_17_i,in_29_18_r,in_29_18_i,in_29_19_r,in_29_19_i,in_29_20_r,in_29_20_i,in_29_21_r,in_29_21_i,in_29_22_r,in_29_22_i,in_29_23_r,in_29_23_i,in_29_24_r,in_29_24_i,in_29_25_r,in_29_25_i,in_29_26_r,in_29_26_i,in_29_27_r,in_29_27_i,in_29_28_r,in_29_28_i,in_29_29_r,in_29_29_i,in_29_30_r,in_29_30_i,in_29_31_r,in_29_31_i,in_29_32_r,in_29_32_i,in_30_1_r,in_30_1_i,in_30_2_r,in_30_2_i,in_30_3_r,in_30_3_i,in_30_4_r,in_30_4_i,in_30_5_r,in_30_5_i,in_30_6_r,in_30_6_i,in_30_7_r,in_30_7_i,in_30_8_r,in_30_8_i,in_30_9_r,in_30_9_i,in_30_10_r,in_30_10_i,in_30_11_r,in_30_11_i,in_30_12_r,in_30_12_i,in_30_13_r,in_30_13_i,in_30_14_r,in_30_14_i,in_30_15_r,in_30_15_i,in_30_16_r,in_30_16_i,in_30_17_r,in_30_17_i,in_30_18_r,in_30_18_i,in_30_19_r,in_30_19_i,in_30_20_r,in_30_20_i,in_30_21_r,in_30_21_i,in_30_22_r,in_30_22_i,in_30_23_r,in_30_23_i,in_30_24_r,in_30_24_i,in_30_25_r,in_30_25_i,in_30_26_r,in_30_26_i,in_30_27_r,in_30_27_i,in_30_28_r,in_30_28_i,in_30_29_r,in_30_29_i,in_30_30_r,in_30_30_i,in_30_31_r,in_30_31_i,in_30_32_r,in_30_32_i,in_31_1_r,in_31_1_i,in_31_2_r,in_31_2_i,in_31_3_r,in_31_3_i,in_31_4_r,in_31_4_i,in_31_5_r,in_31_5_i,in_31_6_r,in_31_6_i,in_31_7_r,in_31_7_i,in_31_8_r,in_31_8_i,in_31_9_r,in_31_9_i,in_31_10_r,in_31_10_i,in_31_11_r,in_31_11_i,in_31_12_r,in_31_12_i,in_31_13_r,in_31_13_i,in_31_14_r,in_31_14_i,in_31_15_r,in_31_15_i,in_31_16_r,in_31_16_i,in_31_17_r,in_31_17_i,in_31_18_r,in_31_18_i,in_31_19_r,in_31_19_i,in_31_20_r,in_31_20_i,in_31_21_r,in_31_21_i,in_31_22_r,in_31_22_i,in_31_23_r,in_31_23_i,in_31_24_r,in_31_24_i,in_31_25_r,in_31_25_i,in_31_26_r,in_31_26_i,in_31_27_r,in_31_27_i,in_31_28_r,in_31_28_i,in_31_29_r,in_31_29_i,in_31_30_r,in_31_30_i,in_31_31_r,in_31_31_i,in_31_32_r,in_31_32_i,in_32_1_r,in_32_1_i,in_32_2_r,in_32_2_i,in_32_3_r,in_32_3_i,in_32_4_r,in_32_4_i,in_32_5_r,in_32_5_i,in_32_6_r,in_32_6_i,in_32_7_r,in_32_7_i,in_32_8_r,in_32_8_i,in_32_9_r,in_32_9_i,in_32_10_r,in_32_10_i,in_32_11_r,in_32_11_i,in_32_12_r,in_32_12_i,in_32_13_r,in_32_13_i,in_32_14_r,in_32_14_i,in_32_15_r,in_32_15_i,in_32_16_r,in_32_16_i,in_32_17_r,in_32_17_i,in_32_18_r,in_32_18_i,in_32_19_r,in_32_19_i,in_32_20_r,in_32_20_i,in_32_21_r,in_32_21_i,in_32_22_r,in_32_22_i,in_32_23_r,in_32_23_i,in_32_24_r,in_32_24_i,in_32_25_r,in_32_25_i,in_32_26_r,in_32_26_i,in_32_27_r,in_32_27_i,in_32_28_r,in_32_28_i,in_32_29_r,in_32_29_i,in_32_30_r,in_32_30_i,in_32_31_r,in_32_31_i,in_32_32_r,in_32_32_i,out_1_1_r,out_1_1_i,out_1_2_r,out_1_2_i,out_1_3_r,out_1_3_i,out_1_4_r,out_1_4_i,out_1_5_r,out_1_5_i,out_1_6_r,out_1_6_i,out_1_7_r,out_1_7_i,out_1_8_r,out_1_8_i,out_1_9_r,out_1_9_i,out_1_10_r,out_1_10_i,out_1_11_r,out_1_11_i,out_1_12_r,out_1_12_i,out_1_13_r,out_1_13_i,out_1_14_r,out_1_14_i,out_1_15_r,out_1_15_i,out_1_16_r,out_1_16_i,out_1_17_r,out_1_17_i,out_1_18_r,out_1_18_i,out_1_19_r,out_1_19_i,out_1_20_r,out_1_20_i,out_1_21_r,out_1_21_i,out_1_22_r,out_1_22_i,out_1_23_r,out_1_23_i,out_1_24_r,out_1_24_i,out_1_25_r,out_1_25_i,out_1_26_r,out_1_26_i,out_1_27_r,out_1_27_i,out_1_28_r,out_1_28_i,out_1_29_r,out_1_29_i,out_1_30_r,out_1_30_i,out_1_31_r,out_1_31_i,out_1_32_r,out_1_32_i,out_2_1_r,out_2_1_i,out_2_2_r,out_2_2_i,out_2_3_r,out_2_3_i,out_2_4_r,out_2_4_i,out_2_5_r,out_2_5_i,out_2_6_r,out_2_6_i,out_2_7_r,out_2_7_i,out_2_8_r,out_2_8_i,out_2_9_r,out_2_9_i,out_2_10_r,out_2_10_i,out_2_11_r,out_2_11_i,out_2_12_r,out_2_12_i,out_2_13_r,out_2_13_i,out_2_14_r,out_2_14_i,out_2_15_r,out_2_15_i,out_2_16_r,out_2_16_i,out_2_17_r,out_2_17_i,out_2_18_r,out_2_18_i,out_2_19_r,out_2_19_i,out_2_20_r,out_2_20_i,out_2_21_r,out_2_21_i,out_2_22_r,out_2_22_i,out_2_23_r,out_2_23_i,out_2_24_r,out_2_24_i,out_2_25_r,out_2_25_i,out_2_26_r,out_2_26_i,out_2_27_r,out_2_27_i,out_2_28_r,out_2_28_i,out_2_29_r,out_2_29_i,out_2_30_r,out_2_30_i,out_2_31_r,out_2_31_i,out_2_32_r,out_2_32_i,out_3_1_r,out_3_1_i,out_3_2_r,out_3_2_i,out_3_3_r,out_3_3_i,out_3_4_r,out_3_4_i,out_3_5_r,out_3_5_i,out_3_6_r,out_3_6_i,out_3_7_r,out_3_7_i,out_3_8_r,out_3_8_i,out_3_9_r,out_3_9_i,out_3_10_r,out_3_10_i,out_3_11_r,out_3_11_i,out_3_12_r,out_3_12_i,out_3_13_r,out_3_13_i,out_3_14_r,out_3_14_i,out_3_15_r,out_3_15_i,out_3_16_r,out_3_16_i,out_3_17_r,out_3_17_i,out_3_18_r,out_3_18_i,out_3_19_r,out_3_19_i,out_3_20_r,out_3_20_i,out_3_21_r,out_3_21_i,out_3_22_r,out_3_22_i,out_3_23_r,out_3_23_i,out_3_24_r,out_3_24_i,out_3_25_r,out_3_25_i,out_3_26_r,out_3_26_i,out_3_27_r,out_3_27_i,out_3_28_r,out_3_28_i,out_3_29_r,out_3_29_i,out_3_30_r,out_3_30_i,out_3_31_r,out_3_31_i,out_3_32_r,out_3_32_i,out_4_1_r,out_4_1_i,out_4_2_r,out_4_2_i,out_4_3_r,out_4_3_i,out_4_4_r,out_4_4_i,out_4_5_r,out_4_5_i,out_4_6_r,out_4_6_i,out_4_7_r,out_4_7_i,out_4_8_r,out_4_8_i,out_4_9_r,out_4_9_i,out_4_10_r,out_4_10_i,out_4_11_r,out_4_11_i,out_4_12_r,out_4_12_i,out_4_13_r,out_4_13_i,out_4_14_r,out_4_14_i,out_4_15_r,out_4_15_i,out_4_16_r,out_4_16_i,out_4_17_r,out_4_17_i,out_4_18_r,out_4_18_i,out_4_19_r,out_4_19_i,out_4_20_r,out_4_20_i,out_4_21_r,out_4_21_i,out_4_22_r,out_4_22_i,out_4_23_r,out_4_23_i,out_4_24_r,out_4_24_i,out_4_25_r,out_4_25_i,out_4_26_r,out_4_26_i,out_4_27_r,out_4_27_i,out_4_28_r,out_4_28_i,out_4_29_r,out_4_29_i,out_4_30_r,out_4_30_i,out_4_31_r,out_4_31_i,out_4_32_r,out_4_32_i,out_5_1_r,out_5_1_i,out_5_2_r,out_5_2_i,out_5_3_r,out_5_3_i,out_5_4_r,out_5_4_i,out_5_5_r,out_5_5_i,out_5_6_r,out_5_6_i,out_5_7_r,out_5_7_i,out_5_8_r,out_5_8_i,out_5_9_r,out_5_9_i,out_5_10_r,out_5_10_i,out_5_11_r,out_5_11_i,out_5_12_r,out_5_12_i,out_5_13_r,out_5_13_i,out_5_14_r,out_5_14_i,out_5_15_r,out_5_15_i,out_5_16_r,out_5_16_i,out_5_17_r,out_5_17_i,out_5_18_r,out_5_18_i,out_5_19_r,out_5_19_i,out_5_20_r,out_5_20_i,out_5_21_r,out_5_21_i,out_5_22_r,out_5_22_i,out_5_23_r,out_5_23_i,out_5_24_r,out_5_24_i,out_5_25_r,out_5_25_i,out_5_26_r,out_5_26_i,out_5_27_r,out_5_27_i,out_5_28_r,out_5_28_i,out_5_29_r,out_5_29_i,out_5_30_r,out_5_30_i,out_5_31_r,out_5_31_i,out_5_32_r,out_5_32_i,out_6_1_r,out_6_1_i,out_6_2_r,out_6_2_i,out_6_3_r,out_6_3_i,out_6_4_r,out_6_4_i,out_6_5_r,out_6_5_i,out_6_6_r,out_6_6_i,out_6_7_r,out_6_7_i,out_6_8_r,out_6_8_i,out_6_9_r,out_6_9_i,out_6_10_r,out_6_10_i,out_6_11_r,out_6_11_i,out_6_12_r,out_6_12_i,out_6_13_r,out_6_13_i,out_6_14_r,out_6_14_i,out_6_15_r,out_6_15_i,out_6_16_r,out_6_16_i,out_6_17_r,out_6_17_i,out_6_18_r,out_6_18_i,out_6_19_r,out_6_19_i,out_6_20_r,out_6_20_i,out_6_21_r,out_6_21_i,out_6_22_r,out_6_22_i,out_6_23_r,out_6_23_i,out_6_24_r,out_6_24_i,out_6_25_r,out_6_25_i,out_6_26_r,out_6_26_i,out_6_27_r,out_6_27_i,out_6_28_r,out_6_28_i,out_6_29_r,out_6_29_i,out_6_30_r,out_6_30_i,out_6_31_r,out_6_31_i,out_6_32_r,out_6_32_i,out_7_1_r,out_7_1_i,out_7_2_r,out_7_2_i,out_7_3_r,out_7_3_i,out_7_4_r,out_7_4_i,out_7_5_r,out_7_5_i,out_7_6_r,out_7_6_i,out_7_7_r,out_7_7_i,out_7_8_r,out_7_8_i,out_7_9_r,out_7_9_i,out_7_10_r,out_7_10_i,out_7_11_r,out_7_11_i,out_7_12_r,out_7_12_i,out_7_13_r,out_7_13_i,out_7_14_r,out_7_14_i,out_7_15_r,out_7_15_i,out_7_16_r,out_7_16_i,out_7_17_r,out_7_17_i,out_7_18_r,out_7_18_i,out_7_19_r,out_7_19_i,out_7_20_r,out_7_20_i,out_7_21_r,out_7_21_i,out_7_22_r,out_7_22_i,out_7_23_r,out_7_23_i,out_7_24_r,out_7_24_i,out_7_25_r,out_7_25_i,out_7_26_r,out_7_26_i,out_7_27_r,out_7_27_i,out_7_28_r,out_7_28_i,out_7_29_r,out_7_29_i,out_7_30_r,out_7_30_i,out_7_31_r,out_7_31_i,out_7_32_r,out_7_32_i,out_8_1_r,out_8_1_i,out_8_2_r,out_8_2_i,out_8_3_r,out_8_3_i,out_8_4_r,out_8_4_i,out_8_5_r,out_8_5_i,out_8_6_r,out_8_6_i,out_8_7_r,out_8_7_i,out_8_8_r,out_8_8_i,out_8_9_r,out_8_9_i,out_8_10_r,out_8_10_i,out_8_11_r,out_8_11_i,out_8_12_r,out_8_12_i,out_8_13_r,out_8_13_i,out_8_14_r,out_8_14_i,out_8_15_r,out_8_15_i,out_8_16_r,out_8_16_i,out_8_17_r,out_8_17_i,out_8_18_r,out_8_18_i,out_8_19_r,out_8_19_i,out_8_20_r,out_8_20_i,out_8_21_r,out_8_21_i,out_8_22_r,out_8_22_i,out_8_23_r,out_8_23_i,out_8_24_r,out_8_24_i,out_8_25_r,out_8_25_i,out_8_26_r,out_8_26_i,out_8_27_r,out_8_27_i,out_8_28_r,out_8_28_i,out_8_29_r,out_8_29_i,out_8_30_r,out_8_30_i,out_8_31_r,out_8_31_i,out_8_32_r,out_8_32_i,out_9_1_r,out_9_1_i,out_9_2_r,out_9_2_i,out_9_3_r,out_9_3_i,out_9_4_r,out_9_4_i,out_9_5_r,out_9_5_i,out_9_6_r,out_9_6_i,out_9_7_r,out_9_7_i,out_9_8_r,out_9_8_i,out_9_9_r,out_9_9_i,out_9_10_r,out_9_10_i,out_9_11_r,out_9_11_i,out_9_12_r,out_9_12_i,out_9_13_r,out_9_13_i,out_9_14_r,out_9_14_i,out_9_15_r,out_9_15_i,out_9_16_r,out_9_16_i,out_9_17_r,out_9_17_i,out_9_18_r,out_9_18_i,out_9_19_r,out_9_19_i,out_9_20_r,out_9_20_i,out_9_21_r,out_9_21_i,out_9_22_r,out_9_22_i,out_9_23_r,out_9_23_i,out_9_24_r,out_9_24_i,out_9_25_r,out_9_25_i,out_9_26_r,out_9_26_i,out_9_27_r,out_9_27_i,out_9_28_r,out_9_28_i,out_9_29_r,out_9_29_i,out_9_30_r,out_9_30_i,out_9_31_r,out_9_31_i,out_9_32_r,out_9_32_i,out_10_1_r,out_10_1_i,out_10_2_r,out_10_2_i,out_10_3_r,out_10_3_i,out_10_4_r,out_10_4_i,out_10_5_r,out_10_5_i,out_10_6_r,out_10_6_i,out_10_7_r,out_10_7_i,out_10_8_r,out_10_8_i,out_10_9_r,out_10_9_i,out_10_10_r,out_10_10_i,out_10_11_r,out_10_11_i,out_10_12_r,out_10_12_i,out_10_13_r,out_10_13_i,out_10_14_r,out_10_14_i,out_10_15_r,out_10_15_i,out_10_16_r,out_10_16_i,out_10_17_r,out_10_17_i,out_10_18_r,out_10_18_i,out_10_19_r,out_10_19_i,out_10_20_r,out_10_20_i,out_10_21_r,out_10_21_i,out_10_22_r,out_10_22_i,out_10_23_r,out_10_23_i,out_10_24_r,out_10_24_i,out_10_25_r,out_10_25_i,out_10_26_r,out_10_26_i,out_10_27_r,out_10_27_i,out_10_28_r,out_10_28_i,out_10_29_r,out_10_29_i,out_10_30_r,out_10_30_i,out_10_31_r,out_10_31_i,out_10_32_r,out_10_32_i,out_11_1_r,out_11_1_i,out_11_2_r,out_11_2_i,out_11_3_r,out_11_3_i,out_11_4_r,out_11_4_i,out_11_5_r,out_11_5_i,out_11_6_r,out_11_6_i,out_11_7_r,out_11_7_i,out_11_8_r,out_11_8_i,out_11_9_r,out_11_9_i,out_11_10_r,out_11_10_i,out_11_11_r,out_11_11_i,out_11_12_r,out_11_12_i,out_11_13_r,out_11_13_i,out_11_14_r,out_11_14_i,out_11_15_r,out_11_15_i,out_11_16_r,out_11_16_i,out_11_17_r,out_11_17_i,out_11_18_r,out_11_18_i,out_11_19_r,out_11_19_i,out_11_20_r,out_11_20_i,out_11_21_r,out_11_21_i,out_11_22_r,out_11_22_i,out_11_23_r,out_11_23_i,out_11_24_r,out_11_24_i,out_11_25_r,out_11_25_i,out_11_26_r,out_11_26_i,out_11_27_r,out_11_27_i,out_11_28_r,out_11_28_i,out_11_29_r,out_11_29_i,out_11_30_r,out_11_30_i,out_11_31_r,out_11_31_i,out_11_32_r,out_11_32_i,out_12_1_r,out_12_1_i,out_12_2_r,out_12_2_i,out_12_3_r,out_12_3_i,out_12_4_r,out_12_4_i,out_12_5_r,out_12_5_i,out_12_6_r,out_12_6_i,out_12_7_r,out_12_7_i,out_12_8_r,out_12_8_i,out_12_9_r,out_12_9_i,out_12_10_r,out_12_10_i,out_12_11_r,out_12_11_i,out_12_12_r,out_12_12_i,out_12_13_r,out_12_13_i,out_12_14_r,out_12_14_i,out_12_15_r,out_12_15_i,out_12_16_r,out_12_16_i,out_12_17_r,out_12_17_i,out_12_18_r,out_12_18_i,out_12_19_r,out_12_19_i,out_12_20_r,out_12_20_i,out_12_21_r,out_12_21_i,out_12_22_r,out_12_22_i,out_12_23_r,out_12_23_i,out_12_24_r,out_12_24_i,out_12_25_r,out_12_25_i,out_12_26_r,out_12_26_i,out_12_27_r,out_12_27_i,out_12_28_r,out_12_28_i,out_12_29_r,out_12_29_i,out_12_30_r,out_12_30_i,out_12_31_r,out_12_31_i,out_12_32_r,out_12_32_i,out_13_1_r,out_13_1_i,out_13_2_r,out_13_2_i,out_13_3_r,out_13_3_i,out_13_4_r,out_13_4_i,out_13_5_r,out_13_5_i,out_13_6_r,out_13_6_i,out_13_7_r,out_13_7_i,out_13_8_r,out_13_8_i,out_13_9_r,out_13_9_i,out_13_10_r,out_13_10_i,out_13_11_r,out_13_11_i,out_13_12_r,out_13_12_i,out_13_13_r,out_13_13_i,out_13_14_r,out_13_14_i,out_13_15_r,out_13_15_i,out_13_16_r,out_13_16_i,out_13_17_r,out_13_17_i,out_13_18_r,out_13_18_i,out_13_19_r,out_13_19_i,out_13_20_r,out_13_20_i,out_13_21_r,out_13_21_i,out_13_22_r,out_13_22_i,out_13_23_r,out_13_23_i,out_13_24_r,out_13_24_i,out_13_25_r,out_13_25_i,out_13_26_r,out_13_26_i,out_13_27_r,out_13_27_i,out_13_28_r,out_13_28_i,out_13_29_r,out_13_29_i,out_13_30_r,out_13_30_i,out_13_31_r,out_13_31_i,out_13_32_r,out_13_32_i,out_14_1_r,out_14_1_i,out_14_2_r,out_14_2_i,out_14_3_r,out_14_3_i,out_14_4_r,out_14_4_i,out_14_5_r,out_14_5_i,out_14_6_r,out_14_6_i,out_14_7_r,out_14_7_i,out_14_8_r,out_14_8_i,out_14_9_r,out_14_9_i,out_14_10_r,out_14_10_i,out_14_11_r,out_14_11_i,out_14_12_r,out_14_12_i,out_14_13_r,out_14_13_i,out_14_14_r,out_14_14_i,out_14_15_r,out_14_15_i,out_14_16_r,out_14_16_i,out_14_17_r,out_14_17_i,out_14_18_r,out_14_18_i,out_14_19_r,out_14_19_i,out_14_20_r,out_14_20_i,out_14_21_r,out_14_21_i,out_14_22_r,out_14_22_i,out_14_23_r,out_14_23_i,out_14_24_r,out_14_24_i,out_14_25_r,out_14_25_i,out_14_26_r,out_14_26_i,out_14_27_r,out_14_27_i,out_14_28_r,out_14_28_i,out_14_29_r,out_14_29_i,out_14_30_r,out_14_30_i,out_14_31_r,out_14_31_i,out_14_32_r,out_14_32_i,out_15_1_r,out_15_1_i,out_15_2_r,out_15_2_i,out_15_3_r,out_15_3_i,out_15_4_r,out_15_4_i,out_15_5_r,out_15_5_i,out_15_6_r,out_15_6_i,out_15_7_r,out_15_7_i,out_15_8_r,out_15_8_i,out_15_9_r,out_15_9_i,out_15_10_r,out_15_10_i,out_15_11_r,out_15_11_i,out_15_12_r,out_15_12_i,out_15_13_r,out_15_13_i,out_15_14_r,out_15_14_i,out_15_15_r,out_15_15_i,out_15_16_r,out_15_16_i,out_15_17_r,out_15_17_i,out_15_18_r,out_15_18_i,out_15_19_r,out_15_19_i,out_15_20_r,out_15_20_i,out_15_21_r,out_15_21_i,out_15_22_r,out_15_22_i,out_15_23_r,out_15_23_i,out_15_24_r,out_15_24_i,out_15_25_r,out_15_25_i,out_15_26_r,out_15_26_i,out_15_27_r,out_15_27_i,out_15_28_r,out_15_28_i,out_15_29_r,out_15_29_i,out_15_30_r,out_15_30_i,out_15_31_r,out_15_31_i,out_15_32_r,out_15_32_i,out_16_1_r,out_16_1_i,out_16_2_r,out_16_2_i,out_16_3_r,out_16_3_i,out_16_4_r,out_16_4_i,out_16_5_r,out_16_5_i,out_16_6_r,out_16_6_i,out_16_7_r,out_16_7_i,out_16_8_r,out_16_8_i,out_16_9_r,out_16_9_i,out_16_10_r,out_16_10_i,out_16_11_r,out_16_11_i,out_16_12_r,out_16_12_i,out_16_13_r,out_16_13_i,out_16_14_r,out_16_14_i,out_16_15_r,out_16_15_i,out_16_16_r,out_16_16_i,out_16_17_r,out_16_17_i,out_16_18_r,out_16_18_i,out_16_19_r,out_16_19_i,out_16_20_r,out_16_20_i,out_16_21_r,out_16_21_i,out_16_22_r,out_16_22_i,out_16_23_r,out_16_23_i,out_16_24_r,out_16_24_i,out_16_25_r,out_16_25_i,out_16_26_r,out_16_26_i,out_16_27_r,out_16_27_i,out_16_28_r,out_16_28_i,out_16_29_r,out_16_29_i,out_16_30_r,out_16_30_i,out_16_31_r,out_16_31_i,out_16_32_r,out_16_32_i,out_17_1_r,out_17_1_i,out_17_2_r,out_17_2_i,out_17_3_r,out_17_3_i,out_17_4_r,out_17_4_i,out_17_5_r,out_17_5_i,out_17_6_r,out_17_6_i,out_17_7_r,out_17_7_i,out_17_8_r,out_17_8_i,out_17_9_r,out_17_9_i,out_17_10_r,out_17_10_i,out_17_11_r,out_17_11_i,out_17_12_r,out_17_12_i,out_17_13_r,out_17_13_i,out_17_14_r,out_17_14_i,out_17_15_r,out_17_15_i,out_17_16_r,out_17_16_i,out_17_17_r,out_17_17_i,out_17_18_r,out_17_18_i,out_17_19_r,out_17_19_i,out_17_20_r,out_17_20_i,out_17_21_r,out_17_21_i,out_17_22_r,out_17_22_i,out_17_23_r,out_17_23_i,out_17_24_r,out_17_24_i,out_17_25_r,out_17_25_i,out_17_26_r,out_17_26_i,out_17_27_r,out_17_27_i,out_17_28_r,out_17_28_i,out_17_29_r,out_17_29_i,out_17_30_r,out_17_30_i,out_17_31_r,out_17_31_i,out_17_32_r,out_17_32_i,out_18_1_r,out_18_1_i,out_18_2_r,out_18_2_i,out_18_3_r,out_18_3_i,out_18_4_r,out_18_4_i,out_18_5_r,out_18_5_i,out_18_6_r,out_18_6_i,out_18_7_r,out_18_7_i,out_18_8_r,out_18_8_i,out_18_9_r,out_18_9_i,out_18_10_r,out_18_10_i,out_18_11_r,out_18_11_i,out_18_12_r,out_18_12_i,out_18_13_r,out_18_13_i,out_18_14_r,out_18_14_i,out_18_15_r,out_18_15_i,out_18_16_r,out_18_16_i,out_18_17_r,out_18_17_i,out_18_18_r,out_18_18_i,out_18_19_r,out_18_19_i,out_18_20_r,out_18_20_i,out_18_21_r,out_18_21_i,out_18_22_r,out_18_22_i,out_18_23_r,out_18_23_i,out_18_24_r,out_18_24_i,out_18_25_r,out_18_25_i,out_18_26_r,out_18_26_i,out_18_27_r,out_18_27_i,out_18_28_r,out_18_28_i,out_18_29_r,out_18_29_i,out_18_30_r,out_18_30_i,out_18_31_r,out_18_31_i,out_18_32_r,out_18_32_i,out_19_1_r,out_19_1_i,out_19_2_r,out_19_2_i,out_19_3_r,out_19_3_i,out_19_4_r,out_19_4_i,out_19_5_r,out_19_5_i,out_19_6_r,out_19_6_i,out_19_7_r,out_19_7_i,out_19_8_r,out_19_8_i,out_19_9_r,out_19_9_i,out_19_10_r,out_19_10_i,out_19_11_r,out_19_11_i,out_19_12_r,out_19_12_i,out_19_13_r,out_19_13_i,out_19_14_r,out_19_14_i,out_19_15_r,out_19_15_i,out_19_16_r,out_19_16_i,out_19_17_r,out_19_17_i,out_19_18_r,out_19_18_i,out_19_19_r,out_19_19_i,out_19_20_r,out_19_20_i,out_19_21_r,out_19_21_i,out_19_22_r,out_19_22_i,out_19_23_r,out_19_23_i,out_19_24_r,out_19_24_i,out_19_25_r,out_19_25_i,out_19_26_r,out_19_26_i,out_19_27_r,out_19_27_i,out_19_28_r,out_19_28_i,out_19_29_r,out_19_29_i,out_19_30_r,out_19_30_i,out_19_31_r,out_19_31_i,out_19_32_r,out_19_32_i,out_20_1_r,out_20_1_i,out_20_2_r,out_20_2_i,out_20_3_r,out_20_3_i,out_20_4_r,out_20_4_i,out_20_5_r,out_20_5_i,out_20_6_r,out_20_6_i,out_20_7_r,out_20_7_i,out_20_8_r,out_20_8_i,out_20_9_r,out_20_9_i,out_20_10_r,out_20_10_i,out_20_11_r,out_20_11_i,out_20_12_r,out_20_12_i,out_20_13_r,out_20_13_i,out_20_14_r,out_20_14_i,out_20_15_r,out_20_15_i,out_20_16_r,out_20_16_i,out_20_17_r,out_20_17_i,out_20_18_r,out_20_18_i,out_20_19_r,out_20_19_i,out_20_20_r,out_20_20_i,out_20_21_r,out_20_21_i,out_20_22_r,out_20_22_i,out_20_23_r,out_20_23_i,out_20_24_r,out_20_24_i,out_20_25_r,out_20_25_i,out_20_26_r,out_20_26_i,out_20_27_r,out_20_27_i,out_20_28_r,out_20_28_i,out_20_29_r,out_20_29_i,out_20_30_r,out_20_30_i,out_20_31_r,out_20_31_i,out_20_32_r,out_20_32_i,out_21_1_r,out_21_1_i,out_21_2_r,out_21_2_i,out_21_3_r,out_21_3_i,out_21_4_r,out_21_4_i,out_21_5_r,out_21_5_i,out_21_6_r,out_21_6_i,out_21_7_r,out_21_7_i,out_21_8_r,out_21_8_i,out_21_9_r,out_21_9_i,out_21_10_r,out_21_10_i,out_21_11_r,out_21_11_i,out_21_12_r,out_21_12_i,out_21_13_r,out_21_13_i,out_21_14_r,out_21_14_i,out_21_15_r,out_21_15_i,out_21_16_r,out_21_16_i,out_21_17_r,out_21_17_i,out_21_18_r,out_21_18_i,out_21_19_r,out_21_19_i,out_21_20_r,out_21_20_i,out_21_21_r,out_21_21_i,out_21_22_r,out_21_22_i,out_21_23_r,out_21_23_i,out_21_24_r,out_21_24_i,out_21_25_r,out_21_25_i,out_21_26_r,out_21_26_i,out_21_27_r,out_21_27_i,out_21_28_r,out_21_28_i,out_21_29_r,out_21_29_i,out_21_30_r,out_21_30_i,out_21_31_r,out_21_31_i,out_21_32_r,out_21_32_i,out_22_1_r,out_22_1_i,out_22_2_r,out_22_2_i,out_22_3_r,out_22_3_i,out_22_4_r,out_22_4_i,out_22_5_r,out_22_5_i,out_22_6_r,out_22_6_i,out_22_7_r,out_22_7_i,out_22_8_r,out_22_8_i,out_22_9_r,out_22_9_i,out_22_10_r,out_22_10_i,out_22_11_r,out_22_11_i,out_22_12_r,out_22_12_i,out_22_13_r,out_22_13_i,out_22_14_r,out_22_14_i,out_22_15_r,out_22_15_i,out_22_16_r,out_22_16_i,out_22_17_r,out_22_17_i,out_22_18_r,out_22_18_i,out_22_19_r,out_22_19_i,out_22_20_r,out_22_20_i,out_22_21_r,out_22_21_i,out_22_22_r,out_22_22_i,out_22_23_r,out_22_23_i,out_22_24_r,out_22_24_i,out_22_25_r,out_22_25_i,out_22_26_r,out_22_26_i,out_22_27_r,out_22_27_i,out_22_28_r,out_22_28_i,out_22_29_r,out_22_29_i,out_22_30_r,out_22_30_i,out_22_31_r,out_22_31_i,out_22_32_r,out_22_32_i,out_23_1_r,out_23_1_i,out_23_2_r,out_23_2_i,out_23_3_r,out_23_3_i,out_23_4_r,out_23_4_i,out_23_5_r,out_23_5_i,out_23_6_r,out_23_6_i,out_23_7_r,out_23_7_i,out_23_8_r,out_23_8_i,out_23_9_r,out_23_9_i,out_23_10_r,out_23_10_i,out_23_11_r,out_23_11_i,out_23_12_r,out_23_12_i,out_23_13_r,out_23_13_i,out_23_14_r,out_23_14_i,out_23_15_r,out_23_15_i,out_23_16_r,out_23_16_i,out_23_17_r,out_23_17_i,out_23_18_r,out_23_18_i,out_23_19_r,out_23_19_i,out_23_20_r,out_23_20_i,out_23_21_r,out_23_21_i,out_23_22_r,out_23_22_i,out_23_23_r,out_23_23_i,out_23_24_r,out_23_24_i,out_23_25_r,out_23_25_i,out_23_26_r,out_23_26_i,out_23_27_r,out_23_27_i,out_23_28_r,out_23_28_i,out_23_29_r,out_23_29_i,out_23_30_r,out_23_30_i,out_23_31_r,out_23_31_i,out_23_32_r,out_23_32_i,out_24_1_r,out_24_1_i,out_24_2_r,out_24_2_i,out_24_3_r,out_24_3_i,out_24_4_r,out_24_4_i,out_24_5_r,out_24_5_i,out_24_6_r,out_24_6_i,out_24_7_r,out_24_7_i,out_24_8_r,out_24_8_i,out_24_9_r,out_24_9_i,out_24_10_r,out_24_10_i,out_24_11_r,out_24_11_i,out_24_12_r,out_24_12_i,out_24_13_r,out_24_13_i,out_24_14_r,out_24_14_i,out_24_15_r,out_24_15_i,out_24_16_r,out_24_16_i,out_24_17_r,out_24_17_i,out_24_18_r,out_24_18_i,out_24_19_r,out_24_19_i,out_24_20_r,out_24_20_i,out_24_21_r,out_24_21_i,out_24_22_r,out_24_22_i,out_24_23_r,out_24_23_i,out_24_24_r,out_24_24_i,out_24_25_r,out_24_25_i,out_24_26_r,out_24_26_i,out_24_27_r,out_24_27_i,out_24_28_r,out_24_28_i,out_24_29_r,out_24_29_i,out_24_30_r,out_24_30_i,out_24_31_r,out_24_31_i,out_24_32_r,out_24_32_i,out_25_1_r,out_25_1_i,out_25_2_r,out_25_2_i,out_25_3_r,out_25_3_i,out_25_4_r,out_25_4_i,out_25_5_r,out_25_5_i,out_25_6_r,out_25_6_i,out_25_7_r,out_25_7_i,out_25_8_r,out_25_8_i,out_25_9_r,out_25_9_i,out_25_10_r,out_25_10_i,out_25_11_r,out_25_11_i,out_25_12_r,out_25_12_i,out_25_13_r,out_25_13_i,out_25_14_r,out_25_14_i,out_25_15_r,out_25_15_i,out_25_16_r,out_25_16_i,out_25_17_r,out_25_17_i,out_25_18_r,out_25_18_i,out_25_19_r,out_25_19_i,out_25_20_r,out_25_20_i,out_25_21_r,out_25_21_i,out_25_22_r,out_25_22_i,out_25_23_r,out_25_23_i,out_25_24_r,out_25_24_i,out_25_25_r,out_25_25_i,out_25_26_r,out_25_26_i,out_25_27_r,out_25_27_i,out_25_28_r,out_25_28_i,out_25_29_r,out_25_29_i,out_25_30_r,out_25_30_i,out_25_31_r,out_25_31_i,out_25_32_r,out_25_32_i,out_26_1_r,out_26_1_i,out_26_2_r,out_26_2_i,out_26_3_r,out_26_3_i,out_26_4_r,out_26_4_i,out_26_5_r,out_26_5_i,out_26_6_r,out_26_6_i,out_26_7_r,out_26_7_i,out_26_8_r,out_26_8_i,out_26_9_r,out_26_9_i,out_26_10_r,out_26_10_i,out_26_11_r,out_26_11_i,out_26_12_r,out_26_12_i,out_26_13_r,out_26_13_i,out_26_14_r,out_26_14_i,out_26_15_r,out_26_15_i,out_26_16_r,out_26_16_i,out_26_17_r,out_26_17_i,out_26_18_r,out_26_18_i,out_26_19_r,out_26_19_i,out_26_20_r,out_26_20_i,out_26_21_r,out_26_21_i,out_26_22_r,out_26_22_i,out_26_23_r,out_26_23_i,out_26_24_r,out_26_24_i,out_26_25_r,out_26_25_i,out_26_26_r,out_26_26_i,out_26_27_r,out_26_27_i,out_26_28_r,out_26_28_i,out_26_29_r,out_26_29_i,out_26_30_r,out_26_30_i,out_26_31_r,out_26_31_i,out_26_32_r,out_26_32_i,out_27_1_r,out_27_1_i,out_27_2_r,out_27_2_i,out_27_3_r,out_27_3_i,out_27_4_r,out_27_4_i,out_27_5_r,out_27_5_i,out_27_6_r,out_27_6_i,out_27_7_r,out_27_7_i,out_27_8_r,out_27_8_i,out_27_9_r,out_27_9_i,out_27_10_r,out_27_10_i,out_27_11_r,out_27_11_i,out_27_12_r,out_27_12_i,out_27_13_r,out_27_13_i,out_27_14_r,out_27_14_i,out_27_15_r,out_27_15_i,out_27_16_r,out_27_16_i,out_27_17_r,out_27_17_i,out_27_18_r,out_27_18_i,out_27_19_r,out_27_19_i,out_27_20_r,out_27_20_i,out_27_21_r,out_27_21_i,out_27_22_r,out_27_22_i,out_27_23_r,out_27_23_i,out_27_24_r,out_27_24_i,out_27_25_r,out_27_25_i,out_27_26_r,out_27_26_i,out_27_27_r,out_27_27_i,out_27_28_r,out_27_28_i,out_27_29_r,out_27_29_i,out_27_30_r,out_27_30_i,out_27_31_r,out_27_31_i,out_27_32_r,out_27_32_i,out_28_1_r,out_28_1_i,out_28_2_r,out_28_2_i,out_28_3_r,out_28_3_i,out_28_4_r,out_28_4_i,out_28_5_r,out_28_5_i,out_28_6_r,out_28_6_i,out_28_7_r,out_28_7_i,out_28_8_r,out_28_8_i,out_28_9_r,out_28_9_i,out_28_10_r,out_28_10_i,out_28_11_r,out_28_11_i,out_28_12_r,out_28_12_i,out_28_13_r,out_28_13_i,out_28_14_r,out_28_14_i,out_28_15_r,out_28_15_i,out_28_16_r,out_28_16_i,out_28_17_r,out_28_17_i,out_28_18_r,out_28_18_i,out_28_19_r,out_28_19_i,out_28_20_r,out_28_20_i,out_28_21_r,out_28_21_i,out_28_22_r,out_28_22_i,out_28_23_r,out_28_23_i,out_28_24_r,out_28_24_i,out_28_25_r,out_28_25_i,out_28_26_r,out_28_26_i,out_28_27_r,out_28_27_i,out_28_28_r,out_28_28_i,out_28_29_r,out_28_29_i,out_28_30_r,out_28_30_i,out_28_31_r,out_28_31_i,out_28_32_r,out_28_32_i,out_29_1_r,out_29_1_i,out_29_2_r,out_29_2_i,out_29_3_r,out_29_3_i,out_29_4_r,out_29_4_i,out_29_5_r,out_29_5_i,out_29_6_r,out_29_6_i,out_29_7_r,out_29_7_i,out_29_8_r,out_29_8_i,out_29_9_r,out_29_9_i,out_29_10_r,out_29_10_i,out_29_11_r,out_29_11_i,out_29_12_r,out_29_12_i,out_29_13_r,out_29_13_i,out_29_14_r,out_29_14_i,out_29_15_r,out_29_15_i,out_29_16_r,out_29_16_i,out_29_17_r,out_29_17_i,out_29_18_r,out_29_18_i,out_29_19_r,out_29_19_i,out_29_20_r,out_29_20_i,out_29_21_r,out_29_21_i,out_29_22_r,out_29_22_i,out_29_23_r,out_29_23_i,out_29_24_r,out_29_24_i,out_29_25_r,out_29_25_i,out_29_26_r,out_29_26_i,out_29_27_r,out_29_27_i,out_29_28_r,out_29_28_i,out_29_29_r,out_29_29_i,out_29_30_r,out_29_30_i,out_29_31_r,out_29_31_i,out_29_32_r,out_29_32_i,out_30_1_r,out_30_1_i,out_30_2_r,out_30_2_i,out_30_3_r,out_30_3_i,out_30_4_r,out_30_4_i,out_30_5_r,out_30_5_i,out_30_6_r,out_30_6_i,out_30_7_r,out_30_7_i,out_30_8_r,out_30_8_i,out_30_9_r,out_30_9_i,out_30_10_r,out_30_10_i,out_30_11_r,out_30_11_i,out_30_12_r,out_30_12_i,out_30_13_r,out_30_13_i,out_30_14_r,out_30_14_i,out_30_15_r,out_30_15_i,out_30_16_r,out_30_16_i,out_30_17_r,out_30_17_i,out_30_18_r,out_30_18_i,out_30_19_r,out_30_19_i,out_30_20_r,out_30_20_i,out_30_21_r,out_30_21_i,out_30_22_r,out_30_22_i,out_30_23_r,out_30_23_i,out_30_24_r,out_30_24_i,out_30_25_r,out_30_25_i,out_30_26_r,out_30_26_i,out_30_27_r,out_30_27_i,out_30_28_r,out_30_28_i,out_30_29_r,out_30_29_i,out_30_30_r,out_30_30_i,out_30_31_r,out_30_31_i,out_30_32_r,out_30_32_i,out_31_1_r,out_31_1_i,out_31_2_r,out_31_2_i,out_31_3_r,out_31_3_i,out_31_4_r,out_31_4_i,out_31_5_r,out_31_5_i,out_31_6_r,out_31_6_i,out_31_7_r,out_31_7_i,out_31_8_r,out_31_8_i,out_31_9_r,out_31_9_i,out_31_10_r,out_31_10_i,out_31_11_r,out_31_11_i,out_31_12_r,out_31_12_i,out_31_13_r,out_31_13_i,out_31_14_r,out_31_14_i,out_31_15_r,out_31_15_i,out_31_16_r,out_31_16_i,out_31_17_r,out_31_17_i,out_31_18_r,out_31_18_i,out_31_19_r,out_31_19_i,out_31_20_r,out_31_20_i,out_31_21_r,out_31_21_i,out_31_22_r,out_31_22_i,out_31_23_r,out_31_23_i,out_31_24_r,out_31_24_i,out_31_25_r,out_31_25_i,out_31_26_r,out_31_26_i,out_31_27_r,out_31_27_i,out_31_28_r,out_31_28_i,out_31_29_r,out_31_29_i,out_31_30_r,out_31_30_i,out_31_31_r,out_31_31_i,out_31_32_r,out_31_32_i,out_32_1_r,out_32_1_i,out_32_2_r,out_32_2_i,out_32_3_r,out_32_3_i,out_32_4_r,out_32_4_i,out_32_5_r,out_32_5_i,out_32_6_r,out_32_6_i,out_32_7_r,out_32_7_i,out_32_8_r,out_32_8_i,out_32_9_r,out_32_9_i,out_32_10_r,out_32_10_i,out_32_11_r,out_32_11_i,out_32_12_r,out_32_12_i,out_32_13_r,out_32_13_i,out_32_14_r,out_32_14_i,out_32_15_r,out_32_15_i,out_32_16_r,out_32_16_i,out_32_17_r,out_32_17_i,out_32_18_r,out_32_18_i,out_32_19_r,out_32_19_i,out_32_20_r,out_32_20_i,out_32_21_r,out_32_21_i,out_32_22_r,out_32_22_i,out_32_23_r,out_32_23_i,out_32_24_r,out_32_24_i,out_32_25_r,out_32_25_i,out_32_26_r,out_32_26_i,out_32_27_r,out_32_27_i,out_32_28_r,out_32_28_i,out_32_29_r,out_32_29_i,out_32_30_r,out_32_30_i,out_32_31_r,out_32_31_i,out_32_32_r,out_32_32_i);
initial begin
clk <= 1'b0;


in_1_1_r <= 16'sb0000000000000010;
in_1_1_i <= 16'sb0000000000000010;

in_1_2_r <= 16'sb0000000000000011;
in_1_2_i <= 16'sb0000000000000011;

in_1_3_r <= 16'sb0000000000000100;
in_1_3_i <= 16'sb0000000000000100;

in_1_4_r <= 16'sb0000000000000101;
in_1_4_i <= 16'sb0000000000000101;

in_1_5_r <= 16'sb0000000000000110;
in_1_5_i <= 16'sb0000000000000110;

in_1_6_r <= 16'sb0000000000000111;
in_1_6_i <= 16'sb0000000000000111;

in_1_7_r <= 16'sb0000000000001000;
in_1_7_i <= 16'sb0000000000001000;

in_1_8_r <= 16'sb0000000000001001;
in_1_8_i <= 16'sb0000000000001001;

in_1_9_r <= 16'sb0000000000001010;
in_1_9_i <= 16'sb0000000000001010;

in_1_10_r <= 16'sb0000000000001011;
in_1_10_i <= 16'sb0000000000001011;

in_1_11_r <= 16'sb0000000000001100;
in_1_11_i <= 16'sb0000000000001100;

in_1_12_r <= 16'sb0000000000001101;
in_1_12_i <= 16'sb0000000000001101;

in_1_13_r <= 16'sb0000000000001110;
in_1_13_i <= 16'sb0000000000001110;

in_1_14_r <= 16'sb0000000000001111;
in_1_14_i <= 16'sb0000000000001111;

in_1_15_r <= 16'sb0000000000010000;
in_1_15_i <= 16'sb0000000000010000;

in_1_16_r <= 16'sb0000000000010001;
in_1_16_i <= 16'sb0000000000010001;

in_1_17_r <= 16'sb0000000000010010;
in_1_17_i <= 16'sb0000000000010010;

in_1_18_r <= 16'sb0000000000010011;
in_1_18_i <= 16'sb0000000000010011;

in_1_19_r <= 16'sb0000000000010100;
in_1_19_i <= 16'sb0000000000010100;

in_1_20_r <= 16'sb0000000000010101;
in_1_20_i <= 16'sb0000000000010101;

in_1_21_r <= 16'sb0000000000010110;
in_1_21_i <= 16'sb0000000000010110;

in_1_22_r <= 16'sb0000000000010111;
in_1_22_i <= 16'sb0000000000010111;

in_1_23_r <= 16'sb0000000000011000;
in_1_23_i <= 16'sb0000000000011000;

in_1_24_r <= 16'sb0000000000011001;
in_1_24_i <= 16'sb0000000000011001;

in_1_25_r <= 16'sb0000000000011010;
in_1_25_i <= 16'sb0000000000011010;

in_1_26_r <= 16'sb0000000000011011;
in_1_26_i <= 16'sb0000000000011011;

in_1_27_r <= 16'sb0000000000011100;
in_1_27_i <= 16'sb0000000000011100;

in_1_28_r <= 16'sb0000000000011101;
in_1_28_i <= 16'sb0000000000011101;

in_1_29_r <= 16'sb0000000000011110;
in_1_29_i <= 16'sb0000000000011110;

in_1_30_r <= 16'sb0000000000011111;
in_1_30_i <= 16'sb0000000000011111;

in_1_31_r <= 16'sb0000000000100000;
in_1_31_i <= 16'sb0000000000100000;

in_1_32_r <= 16'sb0000000000100001;
in_1_32_i <= 16'sb0000000000100001;

in_2_1_r <= 16'sb0000000000000011;
in_2_1_i <= 16'sb0000000000000011;

in_2_2_r <= 16'sb0000000000000100;
in_2_2_i <= 16'sb0000000000000100;

in_2_3_r <= 16'sb0000000000000101;
in_2_3_i <= 16'sb0000000000000101;

in_2_4_r <= 16'sb0000000000000110;
in_2_4_i <= 16'sb0000000000000110;

in_2_5_r <= 16'sb0000000000000111;
in_2_5_i <= 16'sb0000000000000111;

in_2_6_r <= 16'sb0000000000001000;
in_2_6_i <= 16'sb0000000000001000;

in_2_7_r <= 16'sb0000000000001001;
in_2_7_i <= 16'sb0000000000001001;

in_2_8_r <= 16'sb0000000000001010;
in_2_8_i <= 16'sb0000000000001010;

in_2_9_r <= 16'sb0000000000001011;
in_2_9_i <= 16'sb0000000000001011;

in_2_10_r <= 16'sb0000000000001100;
in_2_10_i <= 16'sb0000000000001100;

in_2_11_r <= 16'sb0000000000001101;
in_2_11_i <= 16'sb0000000000001101;

in_2_12_r <= 16'sb0000000000001110;
in_2_12_i <= 16'sb0000000000001110;

in_2_13_r <= 16'sb0000000000001111;
in_2_13_i <= 16'sb0000000000001111;

in_2_14_r <= 16'sb0000000000010000;
in_2_14_i <= 16'sb0000000000010000;

in_2_15_r <= 16'sb0000000000010001;
in_2_15_i <= 16'sb0000000000010001;

in_2_16_r <= 16'sb0000000000010010;
in_2_16_i <= 16'sb0000000000010010;

in_2_17_r <= 16'sb0000000000010011;
in_2_17_i <= 16'sb0000000000010011;

in_2_18_r <= 16'sb0000000000010100;
in_2_18_i <= 16'sb0000000000010100;

in_2_19_r <= 16'sb0000000000010101;
in_2_19_i <= 16'sb0000000000010101;

in_2_20_r <= 16'sb0000000000010110;
in_2_20_i <= 16'sb0000000000010110;

in_2_21_r <= 16'sb0000000000010111;
in_2_21_i <= 16'sb0000000000010111;

in_2_22_r <= 16'sb0000000000011000;
in_2_22_i <= 16'sb0000000000011000;

in_2_23_r <= 16'sb0000000000011001;
in_2_23_i <= 16'sb0000000000011001;

in_2_24_r <= 16'sb0000000000011010;
in_2_24_i <= 16'sb0000000000011010;

in_2_25_r <= 16'sb0000000000011011;
in_2_25_i <= 16'sb0000000000011011;

in_2_26_r <= 16'sb0000000000011100;
in_2_26_i <= 16'sb0000000000011100;

in_2_27_r <= 16'sb0000000000011101;
in_2_27_i <= 16'sb0000000000011101;

in_2_28_r <= 16'sb0000000000011110;
in_2_28_i <= 16'sb0000000000011110;

in_2_29_r <= 16'sb0000000000011111;
in_2_29_i <= 16'sb0000000000011111;

in_2_30_r <= 16'sb0000000000100000;
in_2_30_i <= 16'sb0000000000100000;

in_2_31_r <= 16'sb0000000000100001;
in_2_31_i <= 16'sb0000000000100001;

in_2_32_r <= 16'sb0000000000100010;
in_2_32_i <= 16'sb0000000000100010;

in_3_1_r <= 16'sb0000000000000100;
in_3_1_i <= 16'sb0000000000000100;

in_3_2_r <= 16'sb0000000000000101;
in_3_2_i <= 16'sb0000000000000101;

in_3_3_r <= 16'sb0000000000000110;
in_3_3_i <= 16'sb0000000000000110;

in_3_4_r <= 16'sb0000000000000111;
in_3_4_i <= 16'sb0000000000000111;

in_3_5_r <= 16'sb0000000000001000;
in_3_5_i <= 16'sb0000000000001000;

in_3_6_r <= 16'sb0000000000001001;
in_3_6_i <= 16'sb0000000000001001;

in_3_7_r <= 16'sb0000000000001010;
in_3_7_i <= 16'sb0000000000001010;

in_3_8_r <= 16'sb0000000000001011;
in_3_8_i <= 16'sb0000000000001011;

in_3_9_r <= 16'sb0000000000001100;
in_3_9_i <= 16'sb0000000000001100;

in_3_10_r <= 16'sb0000000000001101;
in_3_10_i <= 16'sb0000000000001101;

in_3_11_r <= 16'sb0000000000001110;
in_3_11_i <= 16'sb0000000000001110;

in_3_12_r <= 16'sb0000000000001111;
in_3_12_i <= 16'sb0000000000001111;

in_3_13_r <= 16'sb0000000000010000;
in_3_13_i <= 16'sb0000000000010000;

in_3_14_r <= 16'sb0000000000010001;
in_3_14_i <= 16'sb0000000000010001;

in_3_15_r <= 16'sb0000000000010010;
in_3_15_i <= 16'sb0000000000010010;

in_3_16_r <= 16'sb0000000000010011;
in_3_16_i <= 16'sb0000000000010011;

in_3_17_r <= 16'sb0000000000010100;
in_3_17_i <= 16'sb0000000000010100;

in_3_18_r <= 16'sb0000000000010101;
in_3_18_i <= 16'sb0000000000010101;

in_3_19_r <= 16'sb0000000000010110;
in_3_19_i <= 16'sb0000000000010110;

in_3_20_r <= 16'sb0000000000010111;
in_3_20_i <= 16'sb0000000000010111;

in_3_21_r <= 16'sb0000000000011000;
in_3_21_i <= 16'sb0000000000011000;

in_3_22_r <= 16'sb0000000000011001;
in_3_22_i <= 16'sb0000000000011001;

in_3_23_r <= 16'sb0000000000011010;
in_3_23_i <= 16'sb0000000000011010;

in_3_24_r <= 16'sb0000000000011011;
in_3_24_i <= 16'sb0000000000011011;

in_3_25_r <= 16'sb0000000000011100;
in_3_25_i <= 16'sb0000000000011100;

in_3_26_r <= 16'sb0000000000011101;
in_3_26_i <= 16'sb0000000000011101;

in_3_27_r <= 16'sb0000000000011110;
in_3_27_i <= 16'sb0000000000011110;

in_3_28_r <= 16'sb0000000000011111;
in_3_28_i <= 16'sb0000000000011111;

in_3_29_r <= 16'sb0000000000100000;
in_3_29_i <= 16'sb0000000000100000;

in_3_30_r <= 16'sb0000000000100001;
in_3_30_i <= 16'sb0000000000100001;

in_3_31_r <= 16'sb0000000000100010;
in_3_31_i <= 16'sb0000000000100010;

in_3_32_r <= 16'sb0000000000100011;
in_3_32_i <= 16'sb0000000000100011;

in_4_1_r <= 16'sb0000000000000101;
in_4_1_i <= 16'sb0000000000000101;

in_4_2_r <= 16'sb0000000000000110;
in_4_2_i <= 16'sb0000000000000110;

in_4_3_r <= 16'sb0000000000000111;
in_4_3_i <= 16'sb0000000000000111;

in_4_4_r <= 16'sb0000000000001000;
in_4_4_i <= 16'sb0000000000001000;

in_4_5_r <= 16'sb0000000000001001;
in_4_5_i <= 16'sb0000000000001001;

in_4_6_r <= 16'sb0000000000001010;
in_4_6_i <= 16'sb0000000000001010;

in_4_7_r <= 16'sb0000000000001011;
in_4_7_i <= 16'sb0000000000001011;

in_4_8_r <= 16'sb0000000000001100;
in_4_8_i <= 16'sb0000000000001100;

in_4_9_r <= 16'sb0000000000001101;
in_4_9_i <= 16'sb0000000000001101;

in_4_10_r <= 16'sb0000000000001110;
in_4_10_i <= 16'sb0000000000001110;

in_4_11_r <= 16'sb0000000000001111;
in_4_11_i <= 16'sb0000000000001111;

in_4_12_r <= 16'sb0000000000010000;
in_4_12_i <= 16'sb0000000000010000;

in_4_13_r <= 16'sb0000000000010001;
in_4_13_i <= 16'sb0000000000010001;

in_4_14_r <= 16'sb0000000000010010;
in_4_14_i <= 16'sb0000000000010010;

in_4_15_r <= 16'sb0000000000010011;
in_4_15_i <= 16'sb0000000000010011;

in_4_16_r <= 16'sb0000000000010100;
in_4_16_i <= 16'sb0000000000010100;

in_4_17_r <= 16'sb0000000000010101;
in_4_17_i <= 16'sb0000000000010101;

in_4_18_r <= 16'sb0000000000010110;
in_4_18_i <= 16'sb0000000000010110;

in_4_19_r <= 16'sb0000000000010111;
in_4_19_i <= 16'sb0000000000010111;

in_4_20_r <= 16'sb0000000000011000;
in_4_20_i <= 16'sb0000000000011000;

in_4_21_r <= 16'sb0000000000011001;
in_4_21_i <= 16'sb0000000000011001;

in_4_22_r <= 16'sb0000000000011010;
in_4_22_i <= 16'sb0000000000011010;

in_4_23_r <= 16'sb0000000000011011;
in_4_23_i <= 16'sb0000000000011011;

in_4_24_r <= 16'sb0000000000011100;
in_4_24_i <= 16'sb0000000000011100;

in_4_25_r <= 16'sb0000000000011101;
in_4_25_i <= 16'sb0000000000011101;

in_4_26_r <= 16'sb0000000000011110;
in_4_26_i <= 16'sb0000000000011110;

in_4_27_r <= 16'sb0000000000011111;
in_4_27_i <= 16'sb0000000000011111;

in_4_28_r <= 16'sb0000000000100000;
in_4_28_i <= 16'sb0000000000100000;

in_4_29_r <= 16'sb0000000000100001;
in_4_29_i <= 16'sb0000000000100001;

in_4_30_r <= 16'sb0000000000100010;
in_4_30_i <= 16'sb0000000000100010;

in_4_31_r <= 16'sb0000000000100011;
in_4_31_i <= 16'sb0000000000100011;

in_4_32_r <= 16'sb0000000000100100;
in_4_32_i <= 16'sb0000000000100100;

in_5_1_r <= 16'sb0000000000000110;
in_5_1_i <= 16'sb0000000000000110;

in_5_2_r <= 16'sb0000000000000111;
in_5_2_i <= 16'sb0000000000000111;

in_5_3_r <= 16'sb0000000000001000;
in_5_3_i <= 16'sb0000000000001000;

in_5_4_r <= 16'sb0000000000001001;
in_5_4_i <= 16'sb0000000000001001;

in_5_5_r <= 16'sb0000000000001010;
in_5_5_i <= 16'sb0000000000001010;

in_5_6_r <= 16'sb0000000000001011;
in_5_6_i <= 16'sb0000000000001011;

in_5_7_r <= 16'sb0000000000001100;
in_5_7_i <= 16'sb0000000000001100;

in_5_8_r <= 16'sb0000000000001101;
in_5_8_i <= 16'sb0000000000001101;

in_5_9_r <= 16'sb0000000000001110;
in_5_9_i <= 16'sb0000000000001110;

in_5_10_r <= 16'sb0000000000001111;
in_5_10_i <= 16'sb0000000000001111;

in_5_11_r <= 16'sb0000000000010000;
in_5_11_i <= 16'sb0000000000010000;

in_5_12_r <= 16'sb0000000000010001;
in_5_12_i <= 16'sb0000000000010001;

in_5_13_r <= 16'sb0000000000010010;
in_5_13_i <= 16'sb0000000000010010;

in_5_14_r <= 16'sb0000000000010011;
in_5_14_i <= 16'sb0000000000010011;

in_5_15_r <= 16'sb0000000000010100;
in_5_15_i <= 16'sb0000000000010100;

in_5_16_r <= 16'sb0000000000010101;
in_5_16_i <= 16'sb0000000000010101;

in_5_17_r <= 16'sb0000000000010110;
in_5_17_i <= 16'sb0000000000010110;

in_5_18_r <= 16'sb0000000000010111;
in_5_18_i <= 16'sb0000000000010111;

in_5_19_r <= 16'sb0000000000011000;
in_5_19_i <= 16'sb0000000000011000;

in_5_20_r <= 16'sb0000000000011001;
in_5_20_i <= 16'sb0000000000011001;

in_5_21_r <= 16'sb0000000000011010;
in_5_21_i <= 16'sb0000000000011010;

in_5_22_r <= 16'sb0000000000011011;
in_5_22_i <= 16'sb0000000000011011;

in_5_23_r <= 16'sb0000000000011100;
in_5_23_i <= 16'sb0000000000011100;

in_5_24_r <= 16'sb0000000000011101;
in_5_24_i <= 16'sb0000000000011101;

in_5_25_r <= 16'sb0000000000011110;
in_5_25_i <= 16'sb0000000000011110;

in_5_26_r <= 16'sb0000000000011111;
in_5_26_i <= 16'sb0000000000011111;

in_5_27_r <= 16'sb0000000000100000;
in_5_27_i <= 16'sb0000000000100000;

in_5_28_r <= 16'sb0000000000100001;
in_5_28_i <= 16'sb0000000000100001;

in_5_29_r <= 16'sb0000000000100010;
in_5_29_i <= 16'sb0000000000100010;

in_5_30_r <= 16'sb0000000000100011;
in_5_30_i <= 16'sb0000000000100011;

in_5_31_r <= 16'sb0000000000100100;
in_5_31_i <= 16'sb0000000000100100;

in_5_32_r <= 16'sb0000000000100101;
in_5_32_i <= 16'sb0000000000100101;

in_6_1_r <= 16'sb0000000000000111;
in_6_1_i <= 16'sb0000000000000111;

in_6_2_r <= 16'sb0000000000001000;
in_6_2_i <= 16'sb0000000000001000;

in_6_3_r <= 16'sb0000000000001001;
in_6_3_i <= 16'sb0000000000001001;

in_6_4_r <= 16'sb0000000000001010;
in_6_4_i <= 16'sb0000000000001010;

in_6_5_r <= 16'sb0000000000001011;
in_6_5_i <= 16'sb0000000000001011;

in_6_6_r <= 16'sb0000000000001100;
in_6_6_i <= 16'sb0000000000001100;

in_6_7_r <= 16'sb0000000000001101;
in_6_7_i <= 16'sb0000000000001101;

in_6_8_r <= 16'sb0000000000001110;
in_6_8_i <= 16'sb0000000000001110;

in_6_9_r <= 16'sb0000000000001111;
in_6_9_i <= 16'sb0000000000001111;

in_6_10_r <= 16'sb0000000000010000;
in_6_10_i <= 16'sb0000000000010000;

in_6_11_r <= 16'sb0000000000010001;
in_6_11_i <= 16'sb0000000000010001;

in_6_12_r <= 16'sb0000000000010010;
in_6_12_i <= 16'sb0000000000010010;

in_6_13_r <= 16'sb0000000000010011;
in_6_13_i <= 16'sb0000000000010011;

in_6_14_r <= 16'sb0000000000010100;
in_6_14_i <= 16'sb0000000000010100;

in_6_15_r <= 16'sb0000000000010101;
in_6_15_i <= 16'sb0000000000010101;

in_6_16_r <= 16'sb0000000000010110;
in_6_16_i <= 16'sb0000000000010110;

in_6_17_r <= 16'sb0000000000010111;
in_6_17_i <= 16'sb0000000000010111;

in_6_18_r <= 16'sb0000000000011000;
in_6_18_i <= 16'sb0000000000011000;

in_6_19_r <= 16'sb0000000000011001;
in_6_19_i <= 16'sb0000000000011001;

in_6_20_r <= 16'sb0000000000011010;
in_6_20_i <= 16'sb0000000000011010;

in_6_21_r <= 16'sb0000000000011011;
in_6_21_i <= 16'sb0000000000011011;

in_6_22_r <= 16'sb0000000000011100;
in_6_22_i <= 16'sb0000000000011100;

in_6_23_r <= 16'sb0000000000011101;
in_6_23_i <= 16'sb0000000000011101;

in_6_24_r <= 16'sb0000000000011110;
in_6_24_i <= 16'sb0000000000011110;

in_6_25_r <= 16'sb0000000000011111;
in_6_25_i <= 16'sb0000000000011111;

in_6_26_r <= 16'sb0000000000100000;
in_6_26_i <= 16'sb0000000000100000;

in_6_27_r <= 16'sb0000000000100001;
in_6_27_i <= 16'sb0000000000100001;

in_6_28_r <= 16'sb0000000000100010;
in_6_28_i <= 16'sb0000000000100010;

in_6_29_r <= 16'sb0000000000100011;
in_6_29_i <= 16'sb0000000000100011;

in_6_30_r <= 16'sb0000000000100100;
in_6_30_i <= 16'sb0000000000100100;

in_6_31_r <= 16'sb0000000000100101;
in_6_31_i <= 16'sb0000000000100101;

in_6_32_r <= 16'sb0000000000100110;
in_6_32_i <= 16'sb0000000000100110;

in_7_1_r <= 16'sb0000000000001000;
in_7_1_i <= 16'sb0000000000001000;

in_7_2_r <= 16'sb0000000000001001;
in_7_2_i <= 16'sb0000000000001001;

in_7_3_r <= 16'sb0000000000001010;
in_7_3_i <= 16'sb0000000000001010;

in_7_4_r <= 16'sb0000000000001011;
in_7_4_i <= 16'sb0000000000001011;

in_7_5_r <= 16'sb0000000000001100;
in_7_5_i <= 16'sb0000000000001100;

in_7_6_r <= 16'sb0000000000001101;
in_7_6_i <= 16'sb0000000000001101;

in_7_7_r <= 16'sb0000000000001110;
in_7_7_i <= 16'sb0000000000001110;

in_7_8_r <= 16'sb0000000000001111;
in_7_8_i <= 16'sb0000000000001111;

in_7_9_r <= 16'sb0000000000010000;
in_7_9_i <= 16'sb0000000000010000;

in_7_10_r <= 16'sb0000000000010001;
in_7_10_i <= 16'sb0000000000010001;

in_7_11_r <= 16'sb0000000000010010;
in_7_11_i <= 16'sb0000000000010010;

in_7_12_r <= 16'sb0000000000010011;
in_7_12_i <= 16'sb0000000000010011;

in_7_13_r <= 16'sb0000000000010100;
in_7_13_i <= 16'sb0000000000010100;

in_7_14_r <= 16'sb0000000000010101;
in_7_14_i <= 16'sb0000000000010101;

in_7_15_r <= 16'sb0000000000010110;
in_7_15_i <= 16'sb0000000000010110;

in_7_16_r <= 16'sb0000000000010111;
in_7_16_i <= 16'sb0000000000010111;

in_7_17_r <= 16'sb0000000000011000;
in_7_17_i <= 16'sb0000000000011000;

in_7_18_r <= 16'sb0000000000011001;
in_7_18_i <= 16'sb0000000000011001;

in_7_19_r <= 16'sb0000000000011010;
in_7_19_i <= 16'sb0000000000011010;

in_7_20_r <= 16'sb0000000000011011;
in_7_20_i <= 16'sb0000000000011011;

in_7_21_r <= 16'sb0000000000011100;
in_7_21_i <= 16'sb0000000000011100;

in_7_22_r <= 16'sb0000000000011101;
in_7_22_i <= 16'sb0000000000011101;

in_7_23_r <= 16'sb0000000000011110;
in_7_23_i <= 16'sb0000000000011110;

in_7_24_r <= 16'sb0000000000011111;
in_7_24_i <= 16'sb0000000000011111;

in_7_25_r <= 16'sb0000000000100000;
in_7_25_i <= 16'sb0000000000100000;

in_7_26_r <= 16'sb0000000000100001;
in_7_26_i <= 16'sb0000000000100001;

in_7_27_r <= 16'sb0000000000100010;
in_7_27_i <= 16'sb0000000000100010;

in_7_28_r <= 16'sb0000000000100011;
in_7_28_i <= 16'sb0000000000100011;

in_7_29_r <= 16'sb0000000000100100;
in_7_29_i <= 16'sb0000000000100100;

in_7_30_r <= 16'sb0000000000100101;
in_7_30_i <= 16'sb0000000000100101;

in_7_31_r <= 16'sb0000000000100110;
in_7_31_i <= 16'sb0000000000100110;

in_7_32_r <= 16'sb0000000000100111;
in_7_32_i <= 16'sb0000000000100111;

in_8_1_r <= 16'sb0000000000001001;
in_8_1_i <= 16'sb0000000000001001;

in_8_2_r <= 16'sb0000000000001010;
in_8_2_i <= 16'sb0000000000001010;

in_8_3_r <= 16'sb0000000000001011;
in_8_3_i <= 16'sb0000000000001011;

in_8_4_r <= 16'sb0000000000001100;
in_8_4_i <= 16'sb0000000000001100;

in_8_5_r <= 16'sb0000000000001101;
in_8_5_i <= 16'sb0000000000001101;

in_8_6_r <= 16'sb0000000000001110;
in_8_6_i <= 16'sb0000000000001110;

in_8_7_r <= 16'sb0000000000001111;
in_8_7_i <= 16'sb0000000000001111;

in_8_8_r <= 16'sb0000000000010000;
in_8_8_i <= 16'sb0000000000010000;

in_8_9_r <= 16'sb0000000000010001;
in_8_9_i <= 16'sb0000000000010001;

in_8_10_r <= 16'sb0000000000010010;
in_8_10_i <= 16'sb0000000000010010;

in_8_11_r <= 16'sb0000000000010011;
in_8_11_i <= 16'sb0000000000010011;

in_8_12_r <= 16'sb0000000000010100;
in_8_12_i <= 16'sb0000000000010100;

in_8_13_r <= 16'sb0000000000010101;
in_8_13_i <= 16'sb0000000000010101;

in_8_14_r <= 16'sb0000000000010110;
in_8_14_i <= 16'sb0000000000010110;

in_8_15_r <= 16'sb0000000000010111;
in_8_15_i <= 16'sb0000000000010111;

in_8_16_r <= 16'sb0000000000011000;
in_8_16_i <= 16'sb0000000000011000;

in_8_17_r <= 16'sb0000000000011001;
in_8_17_i <= 16'sb0000000000011001;

in_8_18_r <= 16'sb0000000000011010;
in_8_18_i <= 16'sb0000000000011010;

in_8_19_r <= 16'sb0000000000011011;
in_8_19_i <= 16'sb0000000000011011;

in_8_20_r <= 16'sb0000000000011100;
in_8_20_i <= 16'sb0000000000011100;

in_8_21_r <= 16'sb0000000000011101;
in_8_21_i <= 16'sb0000000000011101;

in_8_22_r <= 16'sb0000000000011110;
in_8_22_i <= 16'sb0000000000011110;

in_8_23_r <= 16'sb0000000000011111;
in_8_23_i <= 16'sb0000000000011111;

in_8_24_r <= 16'sb0000000000100000;
in_8_24_i <= 16'sb0000000000100000;

in_8_25_r <= 16'sb0000000000100001;
in_8_25_i <= 16'sb0000000000100001;

in_8_26_r <= 16'sb0000000000100010;
in_8_26_i <= 16'sb0000000000100010;

in_8_27_r <= 16'sb0000000000100011;
in_8_27_i <= 16'sb0000000000100011;

in_8_28_r <= 16'sb0000000000100100;
in_8_28_i <= 16'sb0000000000100100;

in_8_29_r <= 16'sb0000000000100101;
in_8_29_i <= 16'sb0000000000100101;

in_8_30_r <= 16'sb0000000000100110;
in_8_30_i <= 16'sb0000000000100110;

in_8_31_r <= 16'sb0000000000100111;
in_8_31_i <= 16'sb0000000000100111;

in_8_32_r <= 16'sb0000000000101000;
in_8_32_i <= 16'sb0000000000101000;

in_9_1_r <= 16'sb0000000000001010;
in_9_1_i <= 16'sb0000000000001010;

in_9_2_r <= 16'sb0000000000001011;
in_9_2_i <= 16'sb0000000000001011;

in_9_3_r <= 16'sb0000000000001100;
in_9_3_i <= 16'sb0000000000001100;

in_9_4_r <= 16'sb0000000000001101;
in_9_4_i <= 16'sb0000000000001101;

in_9_5_r <= 16'sb0000000000001110;
in_9_5_i <= 16'sb0000000000001110;

in_9_6_r <= 16'sb0000000000001111;
in_9_6_i <= 16'sb0000000000001111;

in_9_7_r <= 16'sb0000000000010000;
in_9_7_i <= 16'sb0000000000010000;

in_9_8_r <= 16'sb0000000000010001;
in_9_8_i <= 16'sb0000000000010001;

in_9_9_r <= 16'sb0000000000010010;
in_9_9_i <= 16'sb0000000000010010;

in_9_10_r <= 16'sb0000000000010011;
in_9_10_i <= 16'sb0000000000010011;

in_9_11_r <= 16'sb0000000000010100;
in_9_11_i <= 16'sb0000000000010100;

in_9_12_r <= 16'sb0000000000010101;
in_9_12_i <= 16'sb0000000000010101;

in_9_13_r <= 16'sb0000000000010110;
in_9_13_i <= 16'sb0000000000010110;

in_9_14_r <= 16'sb0000000000010111;
in_9_14_i <= 16'sb0000000000010111;

in_9_15_r <= 16'sb0000000000011000;
in_9_15_i <= 16'sb0000000000011000;

in_9_16_r <= 16'sb0000000000011001;
in_9_16_i <= 16'sb0000000000011001;

in_9_17_r <= 16'sb0000000000011010;
in_9_17_i <= 16'sb0000000000011010;

in_9_18_r <= 16'sb0000000000011011;
in_9_18_i <= 16'sb0000000000011011;

in_9_19_r <= 16'sb0000000000011100;
in_9_19_i <= 16'sb0000000000011100;

in_9_20_r <= 16'sb0000000000011101;
in_9_20_i <= 16'sb0000000000011101;

in_9_21_r <= 16'sb0000000000011110;
in_9_21_i <= 16'sb0000000000011110;

in_9_22_r <= 16'sb0000000000011111;
in_9_22_i <= 16'sb0000000000011111;

in_9_23_r <= 16'sb0000000000100000;
in_9_23_i <= 16'sb0000000000100000;

in_9_24_r <= 16'sb0000000000100001;
in_9_24_i <= 16'sb0000000000100001;

in_9_25_r <= 16'sb0000000000100010;
in_9_25_i <= 16'sb0000000000100010;

in_9_26_r <= 16'sb0000000000100011;
in_9_26_i <= 16'sb0000000000100011;

in_9_27_r <= 16'sb0000000000100100;
in_9_27_i <= 16'sb0000000000100100;

in_9_28_r <= 16'sb0000000000100101;
in_9_28_i <= 16'sb0000000000100101;

in_9_29_r <= 16'sb0000000000100110;
in_9_29_i <= 16'sb0000000000100110;

in_9_30_r <= 16'sb0000000000100111;
in_9_30_i <= 16'sb0000000000100111;

in_9_31_r <= 16'sb0000000000101000;
in_9_31_i <= 16'sb0000000000101000;

in_9_32_r <= 16'sb0000000000101001;
in_9_32_i <= 16'sb0000000000101001;

in_10_1_r <= 16'sb0000000000001011;
in_10_1_i <= 16'sb0000000000001011;

in_10_2_r <= 16'sb0000000000001100;
in_10_2_i <= 16'sb0000000000001100;

in_10_3_r <= 16'sb0000000000001101;
in_10_3_i <= 16'sb0000000000001101;

in_10_4_r <= 16'sb0000000000001110;
in_10_4_i <= 16'sb0000000000001110;

in_10_5_r <= 16'sb0000000000001111;
in_10_5_i <= 16'sb0000000000001111;

in_10_6_r <= 16'sb0000000000010000;
in_10_6_i <= 16'sb0000000000010000;

in_10_7_r <= 16'sb0000000000010001;
in_10_7_i <= 16'sb0000000000010001;

in_10_8_r <= 16'sb0000000000010010;
in_10_8_i <= 16'sb0000000000010010;

in_10_9_r <= 16'sb0000000000010011;
in_10_9_i <= 16'sb0000000000010011;

in_10_10_r <= 16'sb0000000000010100;
in_10_10_i <= 16'sb0000000000010100;

in_10_11_r <= 16'sb0000000000010101;
in_10_11_i <= 16'sb0000000000010101;

in_10_12_r <= 16'sb0000000000010110;
in_10_12_i <= 16'sb0000000000010110;

in_10_13_r <= 16'sb0000000000010111;
in_10_13_i <= 16'sb0000000000010111;

in_10_14_r <= 16'sb0000000000011000;
in_10_14_i <= 16'sb0000000000011000;

in_10_15_r <= 16'sb0000000000011001;
in_10_15_i <= 16'sb0000000000011001;

in_10_16_r <= 16'sb0000000000011010;
in_10_16_i <= 16'sb0000000000011010;

in_10_17_r <= 16'sb0000000000011011;
in_10_17_i <= 16'sb0000000000011011;

in_10_18_r <= 16'sb0000000000011100;
in_10_18_i <= 16'sb0000000000011100;

in_10_19_r <= 16'sb0000000000011101;
in_10_19_i <= 16'sb0000000000011101;

in_10_20_r <= 16'sb0000000000011110;
in_10_20_i <= 16'sb0000000000011110;

in_10_21_r <= 16'sb0000000000011111;
in_10_21_i <= 16'sb0000000000011111;

in_10_22_r <= 16'sb0000000000100000;
in_10_22_i <= 16'sb0000000000100000;

in_10_23_r <= 16'sb0000000000100001;
in_10_23_i <= 16'sb0000000000100001;

in_10_24_r <= 16'sb0000000000100010;
in_10_24_i <= 16'sb0000000000100010;

in_10_25_r <= 16'sb0000000000100011;
in_10_25_i <= 16'sb0000000000100011;

in_10_26_r <= 16'sb0000000000100100;
in_10_26_i <= 16'sb0000000000100100;

in_10_27_r <= 16'sb0000000000100101;
in_10_27_i <= 16'sb0000000000100101;

in_10_28_r <= 16'sb0000000000100110;
in_10_28_i <= 16'sb0000000000100110;

in_10_29_r <= 16'sb0000000000100111;
in_10_29_i <= 16'sb0000000000100111;

in_10_30_r <= 16'sb0000000000101000;
in_10_30_i <= 16'sb0000000000101000;

in_10_31_r <= 16'sb0000000000101001;
in_10_31_i <= 16'sb0000000000101001;

in_10_32_r <= 16'sb0000000000101010;
in_10_32_i <= 16'sb0000000000101010;

in_11_1_r <= 16'sb0000000000001100;
in_11_1_i <= 16'sb0000000000001100;

in_11_2_r <= 16'sb0000000000001101;
in_11_2_i <= 16'sb0000000000001101;

in_11_3_r <= 16'sb0000000000001110;
in_11_3_i <= 16'sb0000000000001110;

in_11_4_r <= 16'sb0000000000001111;
in_11_4_i <= 16'sb0000000000001111;

in_11_5_r <= 16'sb0000000000010000;
in_11_5_i <= 16'sb0000000000010000;

in_11_6_r <= 16'sb0000000000010001;
in_11_6_i <= 16'sb0000000000010001;

in_11_7_r <= 16'sb0000000000010010;
in_11_7_i <= 16'sb0000000000010010;

in_11_8_r <= 16'sb0000000000010011;
in_11_8_i <= 16'sb0000000000010011;

in_11_9_r <= 16'sb0000000000010100;
in_11_9_i <= 16'sb0000000000010100;

in_11_10_r <= 16'sb0000000000010101;
in_11_10_i <= 16'sb0000000000010101;

in_11_11_r <= 16'sb0000000000010110;
in_11_11_i <= 16'sb0000000000010110;

in_11_12_r <= 16'sb0000000000010111;
in_11_12_i <= 16'sb0000000000010111;

in_11_13_r <= 16'sb0000000000011000;
in_11_13_i <= 16'sb0000000000011000;

in_11_14_r <= 16'sb0000000000011001;
in_11_14_i <= 16'sb0000000000011001;

in_11_15_r <= 16'sb0000000000011010;
in_11_15_i <= 16'sb0000000000011010;

in_11_16_r <= 16'sb0000000000011011;
in_11_16_i <= 16'sb0000000000011011;

in_11_17_r <= 16'sb0000000000011100;
in_11_17_i <= 16'sb0000000000011100;

in_11_18_r <= 16'sb0000000000011101;
in_11_18_i <= 16'sb0000000000011101;

in_11_19_r <= 16'sb0000000000011110;
in_11_19_i <= 16'sb0000000000011110;

in_11_20_r <= 16'sb0000000000011111;
in_11_20_i <= 16'sb0000000000011111;

in_11_21_r <= 16'sb0000000000100000;
in_11_21_i <= 16'sb0000000000100000;

in_11_22_r <= 16'sb0000000000100001;
in_11_22_i <= 16'sb0000000000100001;

in_11_23_r <= 16'sb0000000000100010;
in_11_23_i <= 16'sb0000000000100010;

in_11_24_r <= 16'sb0000000000100011;
in_11_24_i <= 16'sb0000000000100011;

in_11_25_r <= 16'sb0000000000100100;
in_11_25_i <= 16'sb0000000000100100;

in_11_26_r <= 16'sb0000000000100101;
in_11_26_i <= 16'sb0000000000100101;

in_11_27_r <= 16'sb0000000000100110;
in_11_27_i <= 16'sb0000000000100110;

in_11_28_r <= 16'sb0000000000100111;
in_11_28_i <= 16'sb0000000000100111;

in_11_29_r <= 16'sb0000000000101000;
in_11_29_i <= 16'sb0000000000101000;

in_11_30_r <= 16'sb0000000000101001;
in_11_30_i <= 16'sb0000000000101001;

in_11_31_r <= 16'sb0000000000101010;
in_11_31_i <= 16'sb0000000000101010;

in_11_32_r <= 16'sb0000000000101011;
in_11_32_i <= 16'sb0000000000101011;

in_12_1_r <= 16'sb0000000000001101;
in_12_1_i <= 16'sb0000000000001101;

in_12_2_r <= 16'sb0000000000001110;
in_12_2_i <= 16'sb0000000000001110;

in_12_3_r <= 16'sb0000000000001111;
in_12_3_i <= 16'sb0000000000001111;

in_12_4_r <= 16'sb0000000000010000;
in_12_4_i <= 16'sb0000000000010000;

in_12_5_r <= 16'sb0000000000010001;
in_12_5_i <= 16'sb0000000000010001;

in_12_6_r <= 16'sb0000000000010010;
in_12_6_i <= 16'sb0000000000010010;

in_12_7_r <= 16'sb0000000000010011;
in_12_7_i <= 16'sb0000000000010011;

in_12_8_r <= 16'sb0000000000010100;
in_12_8_i <= 16'sb0000000000010100;

in_12_9_r <= 16'sb0000000000010101;
in_12_9_i <= 16'sb0000000000010101;

in_12_10_r <= 16'sb0000000000010110;
in_12_10_i <= 16'sb0000000000010110;

in_12_11_r <= 16'sb0000000000010111;
in_12_11_i <= 16'sb0000000000010111;

in_12_12_r <= 16'sb0000000000011000;
in_12_12_i <= 16'sb0000000000011000;

in_12_13_r <= 16'sb0000000000011001;
in_12_13_i <= 16'sb0000000000011001;

in_12_14_r <= 16'sb0000000000011010;
in_12_14_i <= 16'sb0000000000011010;

in_12_15_r <= 16'sb0000000000011011;
in_12_15_i <= 16'sb0000000000011011;

in_12_16_r <= 16'sb0000000000011100;
in_12_16_i <= 16'sb0000000000011100;

in_12_17_r <= 16'sb0000000000011101;
in_12_17_i <= 16'sb0000000000011101;

in_12_18_r <= 16'sb0000000000011110;
in_12_18_i <= 16'sb0000000000011110;

in_12_19_r <= 16'sb0000000000011111;
in_12_19_i <= 16'sb0000000000011111;

in_12_20_r <= 16'sb0000000000100000;
in_12_20_i <= 16'sb0000000000100000;

in_12_21_r <= 16'sb0000000000100001;
in_12_21_i <= 16'sb0000000000100001;

in_12_22_r <= 16'sb0000000000100010;
in_12_22_i <= 16'sb0000000000100010;

in_12_23_r <= 16'sb0000000000100011;
in_12_23_i <= 16'sb0000000000100011;

in_12_24_r <= 16'sb0000000000100100;
in_12_24_i <= 16'sb0000000000100100;

in_12_25_r <= 16'sb0000000000100101;
in_12_25_i <= 16'sb0000000000100101;

in_12_26_r <= 16'sb0000000000100110;
in_12_26_i <= 16'sb0000000000100110;

in_12_27_r <= 16'sb0000000000100111;
in_12_27_i <= 16'sb0000000000100111;

in_12_28_r <= 16'sb0000000000101000;
in_12_28_i <= 16'sb0000000000101000;

in_12_29_r <= 16'sb0000000000101001;
in_12_29_i <= 16'sb0000000000101001;

in_12_30_r <= 16'sb0000000000101010;
in_12_30_i <= 16'sb0000000000101010;

in_12_31_r <= 16'sb0000000000101011;
in_12_31_i <= 16'sb0000000000101011;

in_12_32_r <= 16'sb0000000000101100;
in_12_32_i <= 16'sb0000000000101100;

in_13_1_r <= 16'sb0000000000001110;
in_13_1_i <= 16'sb0000000000001110;

in_13_2_r <= 16'sb0000000000001111;
in_13_2_i <= 16'sb0000000000001111;

in_13_3_r <= 16'sb0000000000010000;
in_13_3_i <= 16'sb0000000000010000;

in_13_4_r <= 16'sb0000000000010001;
in_13_4_i <= 16'sb0000000000010001;

in_13_5_r <= 16'sb0000000000010010;
in_13_5_i <= 16'sb0000000000010010;

in_13_6_r <= 16'sb0000000000010011;
in_13_6_i <= 16'sb0000000000010011;

in_13_7_r <= 16'sb0000000000010100;
in_13_7_i <= 16'sb0000000000010100;

in_13_8_r <= 16'sb0000000000010101;
in_13_8_i <= 16'sb0000000000010101;

in_13_9_r <= 16'sb0000000000010110;
in_13_9_i <= 16'sb0000000000010110;

in_13_10_r <= 16'sb0000000000010111;
in_13_10_i <= 16'sb0000000000010111;

in_13_11_r <= 16'sb0000000000011000;
in_13_11_i <= 16'sb0000000000011000;

in_13_12_r <= 16'sb0000000000011001;
in_13_12_i <= 16'sb0000000000011001;

in_13_13_r <= 16'sb0000000000011010;
in_13_13_i <= 16'sb0000000000011010;

in_13_14_r <= 16'sb0000000000011011;
in_13_14_i <= 16'sb0000000000011011;

in_13_15_r <= 16'sb0000000000011100;
in_13_15_i <= 16'sb0000000000011100;

in_13_16_r <= 16'sb0000000000011101;
in_13_16_i <= 16'sb0000000000011101;

in_13_17_r <= 16'sb0000000000011110;
in_13_17_i <= 16'sb0000000000011110;

in_13_18_r <= 16'sb0000000000011111;
in_13_18_i <= 16'sb0000000000011111;

in_13_19_r <= 16'sb0000000000100000;
in_13_19_i <= 16'sb0000000000100000;

in_13_20_r <= 16'sb0000000000100001;
in_13_20_i <= 16'sb0000000000100001;

in_13_21_r <= 16'sb0000000000100010;
in_13_21_i <= 16'sb0000000000100010;

in_13_22_r <= 16'sb0000000000100011;
in_13_22_i <= 16'sb0000000000100011;

in_13_23_r <= 16'sb0000000000100100;
in_13_23_i <= 16'sb0000000000100100;

in_13_24_r <= 16'sb0000000000100101;
in_13_24_i <= 16'sb0000000000100101;

in_13_25_r <= 16'sb0000000000100110;
in_13_25_i <= 16'sb0000000000100110;

in_13_26_r <= 16'sb0000000000100111;
in_13_26_i <= 16'sb0000000000100111;

in_13_27_r <= 16'sb0000000000101000;
in_13_27_i <= 16'sb0000000000101000;

in_13_28_r <= 16'sb0000000000101001;
in_13_28_i <= 16'sb0000000000101001;

in_13_29_r <= 16'sb0000000000101010;
in_13_29_i <= 16'sb0000000000101010;

in_13_30_r <= 16'sb0000000000101011;
in_13_30_i <= 16'sb0000000000101011;

in_13_31_r <= 16'sb0000000000101100;
in_13_31_i <= 16'sb0000000000101100;

in_13_32_r <= 16'sb0000000000101101;
in_13_32_i <= 16'sb0000000000101101;

in_14_1_r <= 16'sb0000000000001111;
in_14_1_i <= 16'sb0000000000001111;

in_14_2_r <= 16'sb0000000000010000;
in_14_2_i <= 16'sb0000000000010000;

in_14_3_r <= 16'sb0000000000010001;
in_14_3_i <= 16'sb0000000000010001;

in_14_4_r <= 16'sb0000000000010010;
in_14_4_i <= 16'sb0000000000010010;

in_14_5_r <= 16'sb0000000000010011;
in_14_5_i <= 16'sb0000000000010011;

in_14_6_r <= 16'sb0000000000010100;
in_14_6_i <= 16'sb0000000000010100;

in_14_7_r <= 16'sb0000000000010101;
in_14_7_i <= 16'sb0000000000010101;

in_14_8_r <= 16'sb0000000000010110;
in_14_8_i <= 16'sb0000000000010110;

in_14_9_r <= 16'sb0000000000010111;
in_14_9_i <= 16'sb0000000000010111;

in_14_10_r <= 16'sb0000000000011000;
in_14_10_i <= 16'sb0000000000011000;

in_14_11_r <= 16'sb0000000000011001;
in_14_11_i <= 16'sb0000000000011001;

in_14_12_r <= 16'sb0000000000011010;
in_14_12_i <= 16'sb0000000000011010;

in_14_13_r <= 16'sb0000000000011011;
in_14_13_i <= 16'sb0000000000011011;

in_14_14_r <= 16'sb0000000000011100;
in_14_14_i <= 16'sb0000000000011100;

in_14_15_r <= 16'sb0000000000011101;
in_14_15_i <= 16'sb0000000000011101;

in_14_16_r <= 16'sb0000000000011110;
in_14_16_i <= 16'sb0000000000011110;

in_14_17_r <= 16'sb0000000000011111;
in_14_17_i <= 16'sb0000000000011111;

in_14_18_r <= 16'sb0000000000100000;
in_14_18_i <= 16'sb0000000000100000;

in_14_19_r <= 16'sb0000000000100001;
in_14_19_i <= 16'sb0000000000100001;

in_14_20_r <= 16'sb0000000000100010;
in_14_20_i <= 16'sb0000000000100010;

in_14_21_r <= 16'sb0000000000100011;
in_14_21_i <= 16'sb0000000000100011;

in_14_22_r <= 16'sb0000000000100100;
in_14_22_i <= 16'sb0000000000100100;

in_14_23_r <= 16'sb0000000000100101;
in_14_23_i <= 16'sb0000000000100101;

in_14_24_r <= 16'sb0000000000100110;
in_14_24_i <= 16'sb0000000000100110;

in_14_25_r <= 16'sb0000000000100111;
in_14_25_i <= 16'sb0000000000100111;

in_14_26_r <= 16'sb0000000000101000;
in_14_26_i <= 16'sb0000000000101000;

in_14_27_r <= 16'sb0000000000101001;
in_14_27_i <= 16'sb0000000000101001;

in_14_28_r <= 16'sb0000000000101010;
in_14_28_i <= 16'sb0000000000101010;

in_14_29_r <= 16'sb0000000000101011;
in_14_29_i <= 16'sb0000000000101011;

in_14_30_r <= 16'sb0000000000101100;
in_14_30_i <= 16'sb0000000000101100;

in_14_31_r <= 16'sb0000000000101101;
in_14_31_i <= 16'sb0000000000101101;

in_14_32_r <= 16'sb0000000000101110;
in_14_32_i <= 16'sb0000000000101110;

in_15_1_r <= 16'sb0000000000010000;
in_15_1_i <= 16'sb0000000000010000;

in_15_2_r <= 16'sb0000000000010001;
in_15_2_i <= 16'sb0000000000010001;

in_15_3_r <= 16'sb0000000000010010;
in_15_3_i <= 16'sb0000000000010010;

in_15_4_r <= 16'sb0000000000010011;
in_15_4_i <= 16'sb0000000000010011;

in_15_5_r <= 16'sb0000000000010100;
in_15_5_i <= 16'sb0000000000010100;

in_15_6_r <= 16'sb0000000000010101;
in_15_6_i <= 16'sb0000000000010101;

in_15_7_r <= 16'sb0000000000010110;
in_15_7_i <= 16'sb0000000000010110;

in_15_8_r <= 16'sb0000000000010111;
in_15_8_i <= 16'sb0000000000010111;

in_15_9_r <= 16'sb0000000000011000;
in_15_9_i <= 16'sb0000000000011000;

in_15_10_r <= 16'sb0000000000011001;
in_15_10_i <= 16'sb0000000000011001;

in_15_11_r <= 16'sb0000000000011010;
in_15_11_i <= 16'sb0000000000011010;

in_15_12_r <= 16'sb0000000000011011;
in_15_12_i <= 16'sb0000000000011011;

in_15_13_r <= 16'sb0000000000011100;
in_15_13_i <= 16'sb0000000000011100;

in_15_14_r <= 16'sb0000000000011101;
in_15_14_i <= 16'sb0000000000011101;

in_15_15_r <= 16'sb0000000000011110;
in_15_15_i <= 16'sb0000000000011110;

in_15_16_r <= 16'sb0000000000011111;
in_15_16_i <= 16'sb0000000000011111;

in_15_17_r <= 16'sb0000000000100000;
in_15_17_i <= 16'sb0000000000100000;

in_15_18_r <= 16'sb0000000000100001;
in_15_18_i <= 16'sb0000000000100001;

in_15_19_r <= 16'sb0000000000100010;
in_15_19_i <= 16'sb0000000000100010;

in_15_20_r <= 16'sb0000000000100011;
in_15_20_i <= 16'sb0000000000100011;

in_15_21_r <= 16'sb0000000000100100;
in_15_21_i <= 16'sb0000000000100100;

in_15_22_r <= 16'sb0000000000100101;
in_15_22_i <= 16'sb0000000000100101;

in_15_23_r <= 16'sb0000000000100110;
in_15_23_i <= 16'sb0000000000100110;

in_15_24_r <= 16'sb0000000000100111;
in_15_24_i <= 16'sb0000000000100111;

in_15_25_r <= 16'sb0000000000101000;
in_15_25_i <= 16'sb0000000000101000;

in_15_26_r <= 16'sb0000000000101001;
in_15_26_i <= 16'sb0000000000101001;

in_15_27_r <= 16'sb0000000000101010;
in_15_27_i <= 16'sb0000000000101010;

in_15_28_r <= 16'sb0000000000101011;
in_15_28_i <= 16'sb0000000000101011;

in_15_29_r <= 16'sb0000000000101100;
in_15_29_i <= 16'sb0000000000101100;

in_15_30_r <= 16'sb0000000000101101;
in_15_30_i <= 16'sb0000000000101101;

in_15_31_r <= 16'sb0000000000101110;
in_15_31_i <= 16'sb0000000000101110;

in_15_32_r <= 16'sb0000000000101111;
in_15_32_i <= 16'sb0000000000101111;

in_16_1_r <= 16'sb0000000000010001;
in_16_1_i <= 16'sb0000000000010001;

in_16_2_r <= 16'sb0000000000010010;
in_16_2_i <= 16'sb0000000000010010;

in_16_3_r <= 16'sb0000000000010011;
in_16_3_i <= 16'sb0000000000010011;

in_16_4_r <= 16'sb0000000000010100;
in_16_4_i <= 16'sb0000000000010100;

in_16_5_r <= 16'sb0000000000010101;
in_16_5_i <= 16'sb0000000000010101;

in_16_6_r <= 16'sb0000000000010110;
in_16_6_i <= 16'sb0000000000010110;

in_16_7_r <= 16'sb0000000000010111;
in_16_7_i <= 16'sb0000000000010111;

in_16_8_r <= 16'sb0000000000011000;
in_16_8_i <= 16'sb0000000000011000;

in_16_9_r <= 16'sb0000000000011001;
in_16_9_i <= 16'sb0000000000011001;

in_16_10_r <= 16'sb0000000000011010;
in_16_10_i <= 16'sb0000000000011010;

in_16_11_r <= 16'sb0000000000011011;
in_16_11_i <= 16'sb0000000000011011;

in_16_12_r <= 16'sb0000000000011100;
in_16_12_i <= 16'sb0000000000011100;

in_16_13_r <= 16'sb0000000000011101;
in_16_13_i <= 16'sb0000000000011101;

in_16_14_r <= 16'sb0000000000011110;
in_16_14_i <= 16'sb0000000000011110;

in_16_15_r <= 16'sb0000000000011111;
in_16_15_i <= 16'sb0000000000011111;

in_16_16_r <= 16'sb0000000000100000;
in_16_16_i <= 16'sb0000000000100000;

in_16_17_r <= 16'sb0000000000100001;
in_16_17_i <= 16'sb0000000000100001;

in_16_18_r <= 16'sb0000000000100010;
in_16_18_i <= 16'sb0000000000100010;

in_16_19_r <= 16'sb0000000000100011;
in_16_19_i <= 16'sb0000000000100011;

in_16_20_r <= 16'sb0000000000100100;
in_16_20_i <= 16'sb0000000000100100;

in_16_21_r <= 16'sb0000000000100101;
in_16_21_i <= 16'sb0000000000100101;

in_16_22_r <= 16'sb0000000000100110;
in_16_22_i <= 16'sb0000000000100110;

in_16_23_r <= 16'sb0000000000100111;
in_16_23_i <= 16'sb0000000000100111;

in_16_24_r <= 16'sb0000000000101000;
in_16_24_i <= 16'sb0000000000101000;

in_16_25_r <= 16'sb0000000000101001;
in_16_25_i <= 16'sb0000000000101001;

in_16_26_r <= 16'sb0000000000101010;
in_16_26_i <= 16'sb0000000000101010;

in_16_27_r <= 16'sb0000000000101011;
in_16_27_i <= 16'sb0000000000101011;

in_16_28_r <= 16'sb0000000000101100;
in_16_28_i <= 16'sb0000000000101100;

in_16_29_r <= 16'sb0000000000101101;
in_16_29_i <= 16'sb0000000000101101;

in_16_30_r <= 16'sb0000000000101110;
in_16_30_i <= 16'sb0000000000101110;

in_16_31_r <= 16'sb0000000000101111;
in_16_31_i <= 16'sb0000000000101111;

in_16_32_r <= 16'sb0000000000110000;
in_16_32_i <= 16'sb0000000000110000;

in_17_1_r <= 16'sb0000000000010010;
in_17_1_i <= 16'sb0000000000010010;

in_17_2_r <= 16'sb0000000000010011;
in_17_2_i <= 16'sb0000000000010011;

in_17_3_r <= 16'sb0000000000010100;
in_17_3_i <= 16'sb0000000000010100;

in_17_4_r <= 16'sb0000000000010101;
in_17_4_i <= 16'sb0000000000010101;

in_17_5_r <= 16'sb0000000000010110;
in_17_5_i <= 16'sb0000000000010110;

in_17_6_r <= 16'sb0000000000010111;
in_17_6_i <= 16'sb0000000000010111;

in_17_7_r <= 16'sb0000000000011000;
in_17_7_i <= 16'sb0000000000011000;

in_17_8_r <= 16'sb0000000000011001;
in_17_8_i <= 16'sb0000000000011001;

in_17_9_r <= 16'sb0000000000011010;
in_17_9_i <= 16'sb0000000000011010;

in_17_10_r <= 16'sb0000000000011011;
in_17_10_i <= 16'sb0000000000011011;

in_17_11_r <= 16'sb0000000000011100;
in_17_11_i <= 16'sb0000000000011100;

in_17_12_r <= 16'sb0000000000011101;
in_17_12_i <= 16'sb0000000000011101;

in_17_13_r <= 16'sb0000000000011110;
in_17_13_i <= 16'sb0000000000011110;

in_17_14_r <= 16'sb0000000000011111;
in_17_14_i <= 16'sb0000000000011111;

in_17_15_r <= 16'sb0000000000100000;
in_17_15_i <= 16'sb0000000000100000;

in_17_16_r <= 16'sb0000000000100001;
in_17_16_i <= 16'sb0000000000100001;

in_17_17_r <= 16'sb0000000000100010;
in_17_17_i <= 16'sb0000000000100010;

in_17_18_r <= 16'sb0000000000100011;
in_17_18_i <= 16'sb0000000000100011;

in_17_19_r <= 16'sb0000000000100100;
in_17_19_i <= 16'sb0000000000100100;

in_17_20_r <= 16'sb0000000000100101;
in_17_20_i <= 16'sb0000000000100101;

in_17_21_r <= 16'sb0000000000100110;
in_17_21_i <= 16'sb0000000000100110;

in_17_22_r <= 16'sb0000000000100111;
in_17_22_i <= 16'sb0000000000100111;

in_17_23_r <= 16'sb0000000000101000;
in_17_23_i <= 16'sb0000000000101000;

in_17_24_r <= 16'sb0000000000101001;
in_17_24_i <= 16'sb0000000000101001;

in_17_25_r <= 16'sb0000000000101010;
in_17_25_i <= 16'sb0000000000101010;

in_17_26_r <= 16'sb0000000000101011;
in_17_26_i <= 16'sb0000000000101011;

in_17_27_r <= 16'sb0000000000101100;
in_17_27_i <= 16'sb0000000000101100;

in_17_28_r <= 16'sb0000000000101101;
in_17_28_i <= 16'sb0000000000101101;

in_17_29_r <= 16'sb0000000000101110;
in_17_29_i <= 16'sb0000000000101110;

in_17_30_r <= 16'sb0000000000101111;
in_17_30_i <= 16'sb0000000000101111;

in_17_31_r <= 16'sb0000000000110000;
in_17_31_i <= 16'sb0000000000110000;

in_17_32_r <= 16'sb0000000000110001;
in_17_32_i <= 16'sb0000000000110001;

in_18_1_r <= 16'sb0000000000010011;
in_18_1_i <= 16'sb0000000000010011;

in_18_2_r <= 16'sb0000000000010100;
in_18_2_i <= 16'sb0000000000010100;

in_18_3_r <= 16'sb0000000000010101;
in_18_3_i <= 16'sb0000000000010101;

in_18_4_r <= 16'sb0000000000010110;
in_18_4_i <= 16'sb0000000000010110;

in_18_5_r <= 16'sb0000000000010111;
in_18_5_i <= 16'sb0000000000010111;

in_18_6_r <= 16'sb0000000000011000;
in_18_6_i <= 16'sb0000000000011000;

in_18_7_r <= 16'sb0000000000011001;
in_18_7_i <= 16'sb0000000000011001;

in_18_8_r <= 16'sb0000000000011010;
in_18_8_i <= 16'sb0000000000011010;

in_18_9_r <= 16'sb0000000000011011;
in_18_9_i <= 16'sb0000000000011011;

in_18_10_r <= 16'sb0000000000011100;
in_18_10_i <= 16'sb0000000000011100;

in_18_11_r <= 16'sb0000000000011101;
in_18_11_i <= 16'sb0000000000011101;

in_18_12_r <= 16'sb0000000000011110;
in_18_12_i <= 16'sb0000000000011110;

in_18_13_r <= 16'sb0000000000011111;
in_18_13_i <= 16'sb0000000000011111;

in_18_14_r <= 16'sb0000000000100000;
in_18_14_i <= 16'sb0000000000100000;

in_18_15_r <= 16'sb0000000000100001;
in_18_15_i <= 16'sb0000000000100001;

in_18_16_r <= 16'sb0000000000100010;
in_18_16_i <= 16'sb0000000000100010;

in_18_17_r <= 16'sb0000000000100011;
in_18_17_i <= 16'sb0000000000100011;

in_18_18_r <= 16'sb0000000000100100;
in_18_18_i <= 16'sb0000000000100100;

in_18_19_r <= 16'sb0000000000100101;
in_18_19_i <= 16'sb0000000000100101;

in_18_20_r <= 16'sb0000000000100110;
in_18_20_i <= 16'sb0000000000100110;

in_18_21_r <= 16'sb0000000000100111;
in_18_21_i <= 16'sb0000000000100111;

in_18_22_r <= 16'sb0000000000101000;
in_18_22_i <= 16'sb0000000000101000;

in_18_23_r <= 16'sb0000000000101001;
in_18_23_i <= 16'sb0000000000101001;

in_18_24_r <= 16'sb0000000000101010;
in_18_24_i <= 16'sb0000000000101010;

in_18_25_r <= 16'sb0000000000101011;
in_18_25_i <= 16'sb0000000000101011;

in_18_26_r <= 16'sb0000000000101100;
in_18_26_i <= 16'sb0000000000101100;

in_18_27_r <= 16'sb0000000000101101;
in_18_27_i <= 16'sb0000000000101101;

in_18_28_r <= 16'sb0000000000101110;
in_18_28_i <= 16'sb0000000000101110;

in_18_29_r <= 16'sb0000000000101111;
in_18_29_i <= 16'sb0000000000101111;

in_18_30_r <= 16'sb0000000000110000;
in_18_30_i <= 16'sb0000000000110000;

in_18_31_r <= 16'sb0000000000110001;
in_18_31_i <= 16'sb0000000000110001;

in_18_32_r <= 16'sb0000000000110010;
in_18_32_i <= 16'sb0000000000110010;

in_19_1_r <= 16'sb0000000000010100;
in_19_1_i <= 16'sb0000000000010100;

in_19_2_r <= 16'sb0000000000010101;
in_19_2_i <= 16'sb0000000000010101;

in_19_3_r <= 16'sb0000000000010110;
in_19_3_i <= 16'sb0000000000010110;

in_19_4_r <= 16'sb0000000000010111;
in_19_4_i <= 16'sb0000000000010111;

in_19_5_r <= 16'sb0000000000011000;
in_19_5_i <= 16'sb0000000000011000;

in_19_6_r <= 16'sb0000000000011001;
in_19_6_i <= 16'sb0000000000011001;

in_19_7_r <= 16'sb0000000000011010;
in_19_7_i <= 16'sb0000000000011010;

in_19_8_r <= 16'sb0000000000011011;
in_19_8_i <= 16'sb0000000000011011;

in_19_9_r <= 16'sb0000000000011100;
in_19_9_i <= 16'sb0000000000011100;

in_19_10_r <= 16'sb0000000000011101;
in_19_10_i <= 16'sb0000000000011101;

in_19_11_r <= 16'sb0000000000011110;
in_19_11_i <= 16'sb0000000000011110;

in_19_12_r <= 16'sb0000000000011111;
in_19_12_i <= 16'sb0000000000011111;

in_19_13_r <= 16'sb0000000000100000;
in_19_13_i <= 16'sb0000000000100000;

in_19_14_r <= 16'sb0000000000100001;
in_19_14_i <= 16'sb0000000000100001;

in_19_15_r <= 16'sb0000000000100010;
in_19_15_i <= 16'sb0000000000100010;

in_19_16_r <= 16'sb0000000000100011;
in_19_16_i <= 16'sb0000000000100011;

in_19_17_r <= 16'sb0000000000100100;
in_19_17_i <= 16'sb0000000000100100;

in_19_18_r <= 16'sb0000000000100101;
in_19_18_i <= 16'sb0000000000100101;

in_19_19_r <= 16'sb0000000000100110;
in_19_19_i <= 16'sb0000000000100110;

in_19_20_r <= 16'sb0000000000100111;
in_19_20_i <= 16'sb0000000000100111;

in_19_21_r <= 16'sb0000000000101000;
in_19_21_i <= 16'sb0000000000101000;

in_19_22_r <= 16'sb0000000000101001;
in_19_22_i <= 16'sb0000000000101001;

in_19_23_r <= 16'sb0000000000101010;
in_19_23_i <= 16'sb0000000000101010;

in_19_24_r <= 16'sb0000000000101011;
in_19_24_i <= 16'sb0000000000101011;

in_19_25_r <= 16'sb0000000000101100;
in_19_25_i <= 16'sb0000000000101100;

in_19_26_r <= 16'sb0000000000101101;
in_19_26_i <= 16'sb0000000000101101;

in_19_27_r <= 16'sb0000000000101110;
in_19_27_i <= 16'sb0000000000101110;

in_19_28_r <= 16'sb0000000000101111;
in_19_28_i <= 16'sb0000000000101111;

in_19_29_r <= 16'sb0000000000110000;
in_19_29_i <= 16'sb0000000000110000;

in_19_30_r <= 16'sb0000000000110001;
in_19_30_i <= 16'sb0000000000110001;

in_19_31_r <= 16'sb0000000000110010;
in_19_31_i <= 16'sb0000000000110010;

in_19_32_r <= 16'sb0000000000110011;
in_19_32_i <= 16'sb0000000000110011;

in_20_1_r <= 16'sb0000000000010101;
in_20_1_i <= 16'sb0000000000010101;

in_20_2_r <= 16'sb0000000000010110;
in_20_2_i <= 16'sb0000000000010110;

in_20_3_r <= 16'sb0000000000010111;
in_20_3_i <= 16'sb0000000000010111;

in_20_4_r <= 16'sb0000000000011000;
in_20_4_i <= 16'sb0000000000011000;

in_20_5_r <= 16'sb0000000000011001;
in_20_5_i <= 16'sb0000000000011001;

in_20_6_r <= 16'sb0000000000011010;
in_20_6_i <= 16'sb0000000000011010;

in_20_7_r <= 16'sb0000000000011011;
in_20_7_i <= 16'sb0000000000011011;

in_20_8_r <= 16'sb0000000000011100;
in_20_8_i <= 16'sb0000000000011100;

in_20_9_r <= 16'sb0000000000011101;
in_20_9_i <= 16'sb0000000000011101;

in_20_10_r <= 16'sb0000000000011110;
in_20_10_i <= 16'sb0000000000011110;

in_20_11_r <= 16'sb0000000000011111;
in_20_11_i <= 16'sb0000000000011111;

in_20_12_r <= 16'sb0000000000100000;
in_20_12_i <= 16'sb0000000000100000;

in_20_13_r <= 16'sb0000000000100001;
in_20_13_i <= 16'sb0000000000100001;

in_20_14_r <= 16'sb0000000000100010;
in_20_14_i <= 16'sb0000000000100010;

in_20_15_r <= 16'sb0000000000100011;
in_20_15_i <= 16'sb0000000000100011;

in_20_16_r <= 16'sb0000000000100100;
in_20_16_i <= 16'sb0000000000100100;

in_20_17_r <= 16'sb0000000000100101;
in_20_17_i <= 16'sb0000000000100101;

in_20_18_r <= 16'sb0000000000100110;
in_20_18_i <= 16'sb0000000000100110;

in_20_19_r <= 16'sb0000000000100111;
in_20_19_i <= 16'sb0000000000100111;

in_20_20_r <= 16'sb0000000000101000;
in_20_20_i <= 16'sb0000000000101000;

in_20_21_r <= 16'sb0000000000101001;
in_20_21_i <= 16'sb0000000000101001;

in_20_22_r <= 16'sb0000000000101010;
in_20_22_i <= 16'sb0000000000101010;

in_20_23_r <= 16'sb0000000000101011;
in_20_23_i <= 16'sb0000000000101011;

in_20_24_r <= 16'sb0000000000101100;
in_20_24_i <= 16'sb0000000000101100;

in_20_25_r <= 16'sb0000000000101101;
in_20_25_i <= 16'sb0000000000101101;

in_20_26_r <= 16'sb0000000000101110;
in_20_26_i <= 16'sb0000000000101110;

in_20_27_r <= 16'sb0000000000101111;
in_20_27_i <= 16'sb0000000000101111;

in_20_28_r <= 16'sb0000000000110000;
in_20_28_i <= 16'sb0000000000110000;

in_20_29_r <= 16'sb0000000000110001;
in_20_29_i <= 16'sb0000000000110001;

in_20_30_r <= 16'sb0000000000110010;
in_20_30_i <= 16'sb0000000000110010;

in_20_31_r <= 16'sb0000000000110011;
in_20_31_i <= 16'sb0000000000110011;

in_20_32_r <= 16'sb0000000000110100;
in_20_32_i <= 16'sb0000000000110100;

in_21_1_r <= 16'sb0000000000010110;
in_21_1_i <= 16'sb0000000000010110;

in_21_2_r <= 16'sb0000000000010111;
in_21_2_i <= 16'sb0000000000010111;

in_21_3_r <= 16'sb0000000000011000;
in_21_3_i <= 16'sb0000000000011000;

in_21_4_r <= 16'sb0000000000011001;
in_21_4_i <= 16'sb0000000000011001;

in_21_5_r <= 16'sb0000000000011010;
in_21_5_i <= 16'sb0000000000011010;

in_21_6_r <= 16'sb0000000000011011;
in_21_6_i <= 16'sb0000000000011011;

in_21_7_r <= 16'sb0000000000011100;
in_21_7_i <= 16'sb0000000000011100;

in_21_8_r <= 16'sb0000000000011101;
in_21_8_i <= 16'sb0000000000011101;

in_21_9_r <= 16'sb0000000000011110;
in_21_9_i <= 16'sb0000000000011110;

in_21_10_r <= 16'sb0000000000011111;
in_21_10_i <= 16'sb0000000000011111;

in_21_11_r <= 16'sb0000000000100000;
in_21_11_i <= 16'sb0000000000100000;

in_21_12_r <= 16'sb0000000000100001;
in_21_12_i <= 16'sb0000000000100001;

in_21_13_r <= 16'sb0000000000100010;
in_21_13_i <= 16'sb0000000000100010;

in_21_14_r <= 16'sb0000000000100011;
in_21_14_i <= 16'sb0000000000100011;

in_21_15_r <= 16'sb0000000000100100;
in_21_15_i <= 16'sb0000000000100100;

in_21_16_r <= 16'sb0000000000100101;
in_21_16_i <= 16'sb0000000000100101;

in_21_17_r <= 16'sb0000000000100110;
in_21_17_i <= 16'sb0000000000100110;

in_21_18_r <= 16'sb0000000000100111;
in_21_18_i <= 16'sb0000000000100111;

in_21_19_r <= 16'sb0000000000101000;
in_21_19_i <= 16'sb0000000000101000;

in_21_20_r <= 16'sb0000000000101001;
in_21_20_i <= 16'sb0000000000101001;

in_21_21_r <= 16'sb0000000000101010;
in_21_21_i <= 16'sb0000000000101010;

in_21_22_r <= 16'sb0000000000101011;
in_21_22_i <= 16'sb0000000000101011;

in_21_23_r <= 16'sb0000000000101100;
in_21_23_i <= 16'sb0000000000101100;

in_21_24_r <= 16'sb0000000000101101;
in_21_24_i <= 16'sb0000000000101101;

in_21_25_r <= 16'sb0000000000101110;
in_21_25_i <= 16'sb0000000000101110;

in_21_26_r <= 16'sb0000000000101111;
in_21_26_i <= 16'sb0000000000101111;

in_21_27_r <= 16'sb0000000000110000;
in_21_27_i <= 16'sb0000000000110000;

in_21_28_r <= 16'sb0000000000110001;
in_21_28_i <= 16'sb0000000000110001;

in_21_29_r <= 16'sb0000000000110010;
in_21_29_i <= 16'sb0000000000110010;

in_21_30_r <= 16'sb0000000000110011;
in_21_30_i <= 16'sb0000000000110011;

in_21_31_r <= 16'sb0000000000110100;
in_21_31_i <= 16'sb0000000000110100;

in_21_32_r <= 16'sb0000000000110101;
in_21_32_i <= 16'sb0000000000110101;

in_22_1_r <= 16'sb0000000000010111;
in_22_1_i <= 16'sb0000000000010111;

in_22_2_r <= 16'sb0000000000011000;
in_22_2_i <= 16'sb0000000000011000;

in_22_3_r <= 16'sb0000000000011001;
in_22_3_i <= 16'sb0000000000011001;

in_22_4_r <= 16'sb0000000000011010;
in_22_4_i <= 16'sb0000000000011010;

in_22_5_r <= 16'sb0000000000011011;
in_22_5_i <= 16'sb0000000000011011;

in_22_6_r <= 16'sb0000000000011100;
in_22_6_i <= 16'sb0000000000011100;

in_22_7_r <= 16'sb0000000000011101;
in_22_7_i <= 16'sb0000000000011101;

in_22_8_r <= 16'sb0000000000011110;
in_22_8_i <= 16'sb0000000000011110;

in_22_9_r <= 16'sb0000000000011111;
in_22_9_i <= 16'sb0000000000011111;

in_22_10_r <= 16'sb0000000000100000;
in_22_10_i <= 16'sb0000000000100000;

in_22_11_r <= 16'sb0000000000100001;
in_22_11_i <= 16'sb0000000000100001;

in_22_12_r <= 16'sb0000000000100010;
in_22_12_i <= 16'sb0000000000100010;

in_22_13_r <= 16'sb0000000000100011;
in_22_13_i <= 16'sb0000000000100011;

in_22_14_r <= 16'sb0000000000100100;
in_22_14_i <= 16'sb0000000000100100;

in_22_15_r <= 16'sb0000000000100101;
in_22_15_i <= 16'sb0000000000100101;

in_22_16_r <= 16'sb0000000000100110;
in_22_16_i <= 16'sb0000000000100110;

in_22_17_r <= 16'sb0000000000100111;
in_22_17_i <= 16'sb0000000000100111;

in_22_18_r <= 16'sb0000000000101000;
in_22_18_i <= 16'sb0000000000101000;

in_22_19_r <= 16'sb0000000000101001;
in_22_19_i <= 16'sb0000000000101001;

in_22_20_r <= 16'sb0000000000101010;
in_22_20_i <= 16'sb0000000000101010;

in_22_21_r <= 16'sb0000000000101011;
in_22_21_i <= 16'sb0000000000101011;

in_22_22_r <= 16'sb0000000000101100;
in_22_22_i <= 16'sb0000000000101100;

in_22_23_r <= 16'sb0000000000101101;
in_22_23_i <= 16'sb0000000000101101;

in_22_24_r <= 16'sb0000000000101110;
in_22_24_i <= 16'sb0000000000101110;

in_22_25_r <= 16'sb0000000000101111;
in_22_25_i <= 16'sb0000000000101111;

in_22_26_r <= 16'sb0000000000110000;
in_22_26_i <= 16'sb0000000000110000;

in_22_27_r <= 16'sb0000000000110001;
in_22_27_i <= 16'sb0000000000110001;

in_22_28_r <= 16'sb0000000000110010;
in_22_28_i <= 16'sb0000000000110010;

in_22_29_r <= 16'sb0000000000110011;
in_22_29_i <= 16'sb0000000000110011;

in_22_30_r <= 16'sb0000000000110100;
in_22_30_i <= 16'sb0000000000110100;

in_22_31_r <= 16'sb0000000000110101;
in_22_31_i <= 16'sb0000000000110101;

in_22_32_r <= 16'sb0000000000110110;
in_22_32_i <= 16'sb0000000000110110;

in_23_1_r <= 16'sb0000000000011000;
in_23_1_i <= 16'sb0000000000011000;

in_23_2_r <= 16'sb0000000000011001;
in_23_2_i <= 16'sb0000000000011001;

in_23_3_r <= 16'sb0000000000011010;
in_23_3_i <= 16'sb0000000000011010;

in_23_4_r <= 16'sb0000000000011011;
in_23_4_i <= 16'sb0000000000011011;

in_23_5_r <= 16'sb0000000000011100;
in_23_5_i <= 16'sb0000000000011100;

in_23_6_r <= 16'sb0000000000011101;
in_23_6_i <= 16'sb0000000000011101;

in_23_7_r <= 16'sb0000000000011110;
in_23_7_i <= 16'sb0000000000011110;

in_23_8_r <= 16'sb0000000000011111;
in_23_8_i <= 16'sb0000000000011111;

in_23_9_r <= 16'sb0000000000100000;
in_23_9_i <= 16'sb0000000000100000;

in_23_10_r <= 16'sb0000000000100001;
in_23_10_i <= 16'sb0000000000100001;

in_23_11_r <= 16'sb0000000000100010;
in_23_11_i <= 16'sb0000000000100010;

in_23_12_r <= 16'sb0000000000100011;
in_23_12_i <= 16'sb0000000000100011;

in_23_13_r <= 16'sb0000000000100100;
in_23_13_i <= 16'sb0000000000100100;

in_23_14_r <= 16'sb0000000000100101;
in_23_14_i <= 16'sb0000000000100101;

in_23_15_r <= 16'sb0000000000100110;
in_23_15_i <= 16'sb0000000000100110;

in_23_16_r <= 16'sb0000000000100111;
in_23_16_i <= 16'sb0000000000100111;

in_23_17_r <= 16'sb0000000000101000;
in_23_17_i <= 16'sb0000000000101000;

in_23_18_r <= 16'sb0000000000101001;
in_23_18_i <= 16'sb0000000000101001;

in_23_19_r <= 16'sb0000000000101010;
in_23_19_i <= 16'sb0000000000101010;

in_23_20_r <= 16'sb0000000000101011;
in_23_20_i <= 16'sb0000000000101011;

in_23_21_r <= 16'sb0000000000101100;
in_23_21_i <= 16'sb0000000000101100;

in_23_22_r <= 16'sb0000000000101101;
in_23_22_i <= 16'sb0000000000101101;

in_23_23_r <= 16'sb0000000000101110;
in_23_23_i <= 16'sb0000000000101110;

in_23_24_r <= 16'sb0000000000101111;
in_23_24_i <= 16'sb0000000000101111;

in_23_25_r <= 16'sb0000000000110000;
in_23_25_i <= 16'sb0000000000110000;

in_23_26_r <= 16'sb0000000000110001;
in_23_26_i <= 16'sb0000000000110001;

in_23_27_r <= 16'sb0000000000110010;
in_23_27_i <= 16'sb0000000000110010;

in_23_28_r <= 16'sb0000000000110011;
in_23_28_i <= 16'sb0000000000110011;

in_23_29_r <= 16'sb0000000000110100;
in_23_29_i <= 16'sb0000000000110100;

in_23_30_r <= 16'sb0000000000110101;
in_23_30_i <= 16'sb0000000000110101;

in_23_31_r <= 16'sb0000000000110110;
in_23_31_i <= 16'sb0000000000110110;

in_23_32_r <= 16'sb0000000000110111;
in_23_32_i <= 16'sb0000000000110111;

in_24_1_r <= 16'sb0000000000011001;
in_24_1_i <= 16'sb0000000000011001;

in_24_2_r <= 16'sb0000000000011010;
in_24_2_i <= 16'sb0000000000011010;

in_24_3_r <= 16'sb0000000000011011;
in_24_3_i <= 16'sb0000000000011011;

in_24_4_r <= 16'sb0000000000011100;
in_24_4_i <= 16'sb0000000000011100;

in_24_5_r <= 16'sb0000000000011101;
in_24_5_i <= 16'sb0000000000011101;

in_24_6_r <= 16'sb0000000000011110;
in_24_6_i <= 16'sb0000000000011110;

in_24_7_r <= 16'sb0000000000011111;
in_24_7_i <= 16'sb0000000000011111;

in_24_8_r <= 16'sb0000000000100000;
in_24_8_i <= 16'sb0000000000100000;

in_24_9_r <= 16'sb0000000000100001;
in_24_9_i <= 16'sb0000000000100001;

in_24_10_r <= 16'sb0000000000100010;
in_24_10_i <= 16'sb0000000000100010;

in_24_11_r <= 16'sb0000000000100011;
in_24_11_i <= 16'sb0000000000100011;

in_24_12_r <= 16'sb0000000000100100;
in_24_12_i <= 16'sb0000000000100100;

in_24_13_r <= 16'sb0000000000100101;
in_24_13_i <= 16'sb0000000000100101;

in_24_14_r <= 16'sb0000000000100110;
in_24_14_i <= 16'sb0000000000100110;

in_24_15_r <= 16'sb0000000000100111;
in_24_15_i <= 16'sb0000000000100111;

in_24_16_r <= 16'sb0000000000101000;
in_24_16_i <= 16'sb0000000000101000;

in_24_17_r <= 16'sb0000000000101001;
in_24_17_i <= 16'sb0000000000101001;

in_24_18_r <= 16'sb0000000000101010;
in_24_18_i <= 16'sb0000000000101010;

in_24_19_r <= 16'sb0000000000101011;
in_24_19_i <= 16'sb0000000000101011;

in_24_20_r <= 16'sb0000000000101100;
in_24_20_i <= 16'sb0000000000101100;

in_24_21_r <= 16'sb0000000000101101;
in_24_21_i <= 16'sb0000000000101101;

in_24_22_r <= 16'sb0000000000101110;
in_24_22_i <= 16'sb0000000000101110;

in_24_23_r <= 16'sb0000000000101111;
in_24_23_i <= 16'sb0000000000101111;

in_24_24_r <= 16'sb0000000000110000;
in_24_24_i <= 16'sb0000000000110000;

in_24_25_r <= 16'sb0000000000110001;
in_24_25_i <= 16'sb0000000000110001;

in_24_26_r <= 16'sb0000000000110010;
in_24_26_i <= 16'sb0000000000110010;

in_24_27_r <= 16'sb0000000000110011;
in_24_27_i <= 16'sb0000000000110011;

in_24_28_r <= 16'sb0000000000110100;
in_24_28_i <= 16'sb0000000000110100;

in_24_29_r <= 16'sb0000000000110101;
in_24_29_i <= 16'sb0000000000110101;

in_24_30_r <= 16'sb0000000000110110;
in_24_30_i <= 16'sb0000000000110110;

in_24_31_r <= 16'sb0000000000110111;
in_24_31_i <= 16'sb0000000000110111;

in_24_32_r <= 16'sb0000000000111000;
in_24_32_i <= 16'sb0000000000111000;

in_25_1_r <= 16'sb0000000000011010;
in_25_1_i <= 16'sb0000000000011010;

in_25_2_r <= 16'sb0000000000011011;
in_25_2_i <= 16'sb0000000000011011;

in_25_3_r <= 16'sb0000000000011100;
in_25_3_i <= 16'sb0000000000011100;

in_25_4_r <= 16'sb0000000000011101;
in_25_4_i <= 16'sb0000000000011101;

in_25_5_r <= 16'sb0000000000011110;
in_25_5_i <= 16'sb0000000000011110;

in_25_6_r <= 16'sb0000000000011111;
in_25_6_i <= 16'sb0000000000011111;

in_25_7_r <= 16'sb0000000000100000;
in_25_7_i <= 16'sb0000000000100000;

in_25_8_r <= 16'sb0000000000100001;
in_25_8_i <= 16'sb0000000000100001;

in_25_9_r <= 16'sb0000000000100010;
in_25_9_i <= 16'sb0000000000100010;

in_25_10_r <= 16'sb0000000000100011;
in_25_10_i <= 16'sb0000000000100011;

in_25_11_r <= 16'sb0000000000100100;
in_25_11_i <= 16'sb0000000000100100;

in_25_12_r <= 16'sb0000000000100101;
in_25_12_i <= 16'sb0000000000100101;

in_25_13_r <= 16'sb0000000000100110;
in_25_13_i <= 16'sb0000000000100110;

in_25_14_r <= 16'sb0000000000100111;
in_25_14_i <= 16'sb0000000000100111;

in_25_15_r <= 16'sb0000000000101000;
in_25_15_i <= 16'sb0000000000101000;

in_25_16_r <= 16'sb0000000000101001;
in_25_16_i <= 16'sb0000000000101001;

in_25_17_r <= 16'sb0000000000101010;
in_25_17_i <= 16'sb0000000000101010;

in_25_18_r <= 16'sb0000000000101011;
in_25_18_i <= 16'sb0000000000101011;

in_25_19_r <= 16'sb0000000000101100;
in_25_19_i <= 16'sb0000000000101100;

in_25_20_r <= 16'sb0000000000101101;
in_25_20_i <= 16'sb0000000000101101;

in_25_21_r <= 16'sb0000000000101110;
in_25_21_i <= 16'sb0000000000101110;

in_25_22_r <= 16'sb0000000000101111;
in_25_22_i <= 16'sb0000000000101111;

in_25_23_r <= 16'sb0000000000110000;
in_25_23_i <= 16'sb0000000000110000;

in_25_24_r <= 16'sb0000000000110001;
in_25_24_i <= 16'sb0000000000110001;

in_25_25_r <= 16'sb0000000000110010;
in_25_25_i <= 16'sb0000000000110010;

in_25_26_r <= 16'sb0000000000110011;
in_25_26_i <= 16'sb0000000000110011;

in_25_27_r <= 16'sb0000000000110100;
in_25_27_i <= 16'sb0000000000110100;

in_25_28_r <= 16'sb0000000000110101;
in_25_28_i <= 16'sb0000000000110101;

in_25_29_r <= 16'sb0000000000110110;
in_25_29_i <= 16'sb0000000000110110;

in_25_30_r <= 16'sb0000000000110111;
in_25_30_i <= 16'sb0000000000110111;

in_25_31_r <= 16'sb0000000000111000;
in_25_31_i <= 16'sb0000000000111000;

in_25_32_r <= 16'sb0000000000111001;
in_25_32_i <= 16'sb0000000000111001;

in_26_1_r <= 16'sb0000000000011011;
in_26_1_i <= 16'sb0000000000011011;

in_26_2_r <= 16'sb0000000000011100;
in_26_2_i <= 16'sb0000000000011100;

in_26_3_r <= 16'sb0000000000011101;
in_26_3_i <= 16'sb0000000000011101;

in_26_4_r <= 16'sb0000000000011110;
in_26_4_i <= 16'sb0000000000011110;

in_26_5_r <= 16'sb0000000000011111;
in_26_5_i <= 16'sb0000000000011111;

in_26_6_r <= 16'sb0000000000100000;
in_26_6_i <= 16'sb0000000000100000;

in_26_7_r <= 16'sb0000000000100001;
in_26_7_i <= 16'sb0000000000100001;

in_26_8_r <= 16'sb0000000000100010;
in_26_8_i <= 16'sb0000000000100010;

in_26_9_r <= 16'sb0000000000100011;
in_26_9_i <= 16'sb0000000000100011;

in_26_10_r <= 16'sb0000000000100100;
in_26_10_i <= 16'sb0000000000100100;

in_26_11_r <= 16'sb0000000000100101;
in_26_11_i <= 16'sb0000000000100101;

in_26_12_r <= 16'sb0000000000100110;
in_26_12_i <= 16'sb0000000000100110;

in_26_13_r <= 16'sb0000000000100111;
in_26_13_i <= 16'sb0000000000100111;

in_26_14_r <= 16'sb0000000000101000;
in_26_14_i <= 16'sb0000000000101000;

in_26_15_r <= 16'sb0000000000101001;
in_26_15_i <= 16'sb0000000000101001;

in_26_16_r <= 16'sb0000000000101010;
in_26_16_i <= 16'sb0000000000101010;

in_26_17_r <= 16'sb0000000000101011;
in_26_17_i <= 16'sb0000000000101011;

in_26_18_r <= 16'sb0000000000101100;
in_26_18_i <= 16'sb0000000000101100;

in_26_19_r <= 16'sb0000000000101101;
in_26_19_i <= 16'sb0000000000101101;

in_26_20_r <= 16'sb0000000000101110;
in_26_20_i <= 16'sb0000000000101110;

in_26_21_r <= 16'sb0000000000101111;
in_26_21_i <= 16'sb0000000000101111;

in_26_22_r <= 16'sb0000000000110000;
in_26_22_i <= 16'sb0000000000110000;

in_26_23_r <= 16'sb0000000000110001;
in_26_23_i <= 16'sb0000000000110001;

in_26_24_r <= 16'sb0000000000110010;
in_26_24_i <= 16'sb0000000000110010;

in_26_25_r <= 16'sb0000000000110011;
in_26_25_i <= 16'sb0000000000110011;

in_26_26_r <= 16'sb0000000000110100;
in_26_26_i <= 16'sb0000000000110100;

in_26_27_r <= 16'sb0000000000110101;
in_26_27_i <= 16'sb0000000000110101;

in_26_28_r <= 16'sb0000000000110110;
in_26_28_i <= 16'sb0000000000110110;

in_26_29_r <= 16'sb0000000000110111;
in_26_29_i <= 16'sb0000000000110111;

in_26_30_r <= 16'sb0000000000111000;
in_26_30_i <= 16'sb0000000000111000;

in_26_31_r <= 16'sb0000000000111001;
in_26_31_i <= 16'sb0000000000111001;

in_26_32_r <= 16'sb0000000000111010;
in_26_32_i <= 16'sb0000000000111010;

in_27_1_r <= 16'sb0000000000011100;
in_27_1_i <= 16'sb0000000000011100;

in_27_2_r <= 16'sb0000000000011101;
in_27_2_i <= 16'sb0000000000011101;

in_27_3_r <= 16'sb0000000000011110;
in_27_3_i <= 16'sb0000000000011110;

in_27_4_r <= 16'sb0000000000011111;
in_27_4_i <= 16'sb0000000000011111;

in_27_5_r <= 16'sb0000000000100000;
in_27_5_i <= 16'sb0000000000100000;

in_27_6_r <= 16'sb0000000000100001;
in_27_6_i <= 16'sb0000000000100001;

in_27_7_r <= 16'sb0000000000100010;
in_27_7_i <= 16'sb0000000000100010;

in_27_8_r <= 16'sb0000000000100011;
in_27_8_i <= 16'sb0000000000100011;

in_27_9_r <= 16'sb0000000000100100;
in_27_9_i <= 16'sb0000000000100100;

in_27_10_r <= 16'sb0000000000100101;
in_27_10_i <= 16'sb0000000000100101;

in_27_11_r <= 16'sb0000000000100110;
in_27_11_i <= 16'sb0000000000100110;

in_27_12_r <= 16'sb0000000000100111;
in_27_12_i <= 16'sb0000000000100111;

in_27_13_r <= 16'sb0000000000101000;
in_27_13_i <= 16'sb0000000000101000;

in_27_14_r <= 16'sb0000000000101001;
in_27_14_i <= 16'sb0000000000101001;

in_27_15_r <= 16'sb0000000000101010;
in_27_15_i <= 16'sb0000000000101010;

in_27_16_r <= 16'sb0000000000101011;
in_27_16_i <= 16'sb0000000000101011;

in_27_17_r <= 16'sb0000000000101100;
in_27_17_i <= 16'sb0000000000101100;

in_27_18_r <= 16'sb0000000000101101;
in_27_18_i <= 16'sb0000000000101101;

in_27_19_r <= 16'sb0000000000101110;
in_27_19_i <= 16'sb0000000000101110;

in_27_20_r <= 16'sb0000000000101111;
in_27_20_i <= 16'sb0000000000101111;

in_27_21_r <= 16'sb0000000000110000;
in_27_21_i <= 16'sb0000000000110000;

in_27_22_r <= 16'sb0000000000110001;
in_27_22_i <= 16'sb0000000000110001;

in_27_23_r <= 16'sb0000000000110010;
in_27_23_i <= 16'sb0000000000110010;

in_27_24_r <= 16'sb0000000000110011;
in_27_24_i <= 16'sb0000000000110011;

in_27_25_r <= 16'sb0000000000110100;
in_27_25_i <= 16'sb0000000000110100;

in_27_26_r <= 16'sb0000000000110101;
in_27_26_i <= 16'sb0000000000110101;

in_27_27_r <= 16'sb0000000000110110;
in_27_27_i <= 16'sb0000000000110110;

in_27_28_r <= 16'sb0000000000110111;
in_27_28_i <= 16'sb0000000000110111;

in_27_29_r <= 16'sb0000000000111000;
in_27_29_i <= 16'sb0000000000111000;

in_27_30_r <= 16'sb0000000000111001;
in_27_30_i <= 16'sb0000000000111001;

in_27_31_r <= 16'sb0000000000111010;
in_27_31_i <= 16'sb0000000000111010;

in_27_32_r <= 16'sb0000000000111011;
in_27_32_i <= 16'sb0000000000111011;

in_28_1_r <= 16'sb0000000000011101;
in_28_1_i <= 16'sb0000000000011101;

in_28_2_r <= 16'sb0000000000011110;
in_28_2_i <= 16'sb0000000000011110;

in_28_3_r <= 16'sb0000000000011111;
in_28_3_i <= 16'sb0000000000011111;

in_28_4_r <= 16'sb0000000000100000;
in_28_4_i <= 16'sb0000000000100000;

in_28_5_r <= 16'sb0000000000100001;
in_28_5_i <= 16'sb0000000000100001;

in_28_6_r <= 16'sb0000000000100010;
in_28_6_i <= 16'sb0000000000100010;

in_28_7_r <= 16'sb0000000000100011;
in_28_7_i <= 16'sb0000000000100011;

in_28_8_r <= 16'sb0000000000100100;
in_28_8_i <= 16'sb0000000000100100;

in_28_9_r <= 16'sb0000000000100101;
in_28_9_i <= 16'sb0000000000100101;

in_28_10_r <= 16'sb0000000000100110;
in_28_10_i <= 16'sb0000000000100110;

in_28_11_r <= 16'sb0000000000100111;
in_28_11_i <= 16'sb0000000000100111;

in_28_12_r <= 16'sb0000000000101000;
in_28_12_i <= 16'sb0000000000101000;

in_28_13_r <= 16'sb0000000000101001;
in_28_13_i <= 16'sb0000000000101001;

in_28_14_r <= 16'sb0000000000101010;
in_28_14_i <= 16'sb0000000000101010;

in_28_15_r <= 16'sb0000000000101011;
in_28_15_i <= 16'sb0000000000101011;

in_28_16_r <= 16'sb0000000000101100;
in_28_16_i <= 16'sb0000000000101100;

in_28_17_r <= 16'sb0000000000101101;
in_28_17_i <= 16'sb0000000000101101;

in_28_18_r <= 16'sb0000000000101110;
in_28_18_i <= 16'sb0000000000101110;

in_28_19_r <= 16'sb0000000000101111;
in_28_19_i <= 16'sb0000000000101111;

in_28_20_r <= 16'sb0000000000110000;
in_28_20_i <= 16'sb0000000000110000;

in_28_21_r <= 16'sb0000000000110001;
in_28_21_i <= 16'sb0000000000110001;

in_28_22_r <= 16'sb0000000000110010;
in_28_22_i <= 16'sb0000000000110010;

in_28_23_r <= 16'sb0000000000110011;
in_28_23_i <= 16'sb0000000000110011;

in_28_24_r <= 16'sb0000000000110100;
in_28_24_i <= 16'sb0000000000110100;

in_28_25_r <= 16'sb0000000000110101;
in_28_25_i <= 16'sb0000000000110101;

in_28_26_r <= 16'sb0000000000110110;
in_28_26_i <= 16'sb0000000000110110;

in_28_27_r <= 16'sb0000000000110111;
in_28_27_i <= 16'sb0000000000110111;

in_28_28_r <= 16'sb0000000000111000;
in_28_28_i <= 16'sb0000000000111000;

in_28_29_r <= 16'sb0000000000111001;
in_28_29_i <= 16'sb0000000000111001;

in_28_30_r <= 16'sb0000000000111010;
in_28_30_i <= 16'sb0000000000111010;

in_28_31_r <= 16'sb0000000000111011;
in_28_31_i <= 16'sb0000000000111011;

in_28_32_r <= 16'sb0000000000111100;
in_28_32_i <= 16'sb0000000000111100;

in_29_1_r <= 16'sb0000000000011110;
in_29_1_i <= 16'sb0000000000011110;

in_29_2_r <= 16'sb0000000000011111;
in_29_2_i <= 16'sb0000000000011111;

in_29_3_r <= 16'sb0000000000100000;
in_29_3_i <= 16'sb0000000000100000;

in_29_4_r <= 16'sb0000000000100001;
in_29_4_i <= 16'sb0000000000100001;

in_29_5_r <= 16'sb0000000000100010;
in_29_5_i <= 16'sb0000000000100010;

in_29_6_r <= 16'sb0000000000100011;
in_29_6_i <= 16'sb0000000000100011;

in_29_7_r <= 16'sb0000000000100100;
in_29_7_i <= 16'sb0000000000100100;

in_29_8_r <= 16'sb0000000000100101;
in_29_8_i <= 16'sb0000000000100101;

in_29_9_r <= 16'sb0000000000100110;
in_29_9_i <= 16'sb0000000000100110;

in_29_10_r <= 16'sb0000000000100111;
in_29_10_i <= 16'sb0000000000100111;

in_29_11_r <= 16'sb0000000000101000;
in_29_11_i <= 16'sb0000000000101000;

in_29_12_r <= 16'sb0000000000101001;
in_29_12_i <= 16'sb0000000000101001;

in_29_13_r <= 16'sb0000000000101010;
in_29_13_i <= 16'sb0000000000101010;

in_29_14_r <= 16'sb0000000000101011;
in_29_14_i <= 16'sb0000000000101011;

in_29_15_r <= 16'sb0000000000101100;
in_29_15_i <= 16'sb0000000000101100;

in_29_16_r <= 16'sb0000000000101101;
in_29_16_i <= 16'sb0000000000101101;

in_29_17_r <= 16'sb0000000000101110;
in_29_17_i <= 16'sb0000000000101110;

in_29_18_r <= 16'sb0000000000101111;
in_29_18_i <= 16'sb0000000000101111;

in_29_19_r <= 16'sb0000000000110000;
in_29_19_i <= 16'sb0000000000110000;

in_29_20_r <= 16'sb0000000000110001;
in_29_20_i <= 16'sb0000000000110001;

in_29_21_r <= 16'sb0000000000110010;
in_29_21_i <= 16'sb0000000000110010;

in_29_22_r <= 16'sb0000000000110011;
in_29_22_i <= 16'sb0000000000110011;

in_29_23_r <= 16'sb0000000000110100;
in_29_23_i <= 16'sb0000000000110100;

in_29_24_r <= 16'sb0000000000110101;
in_29_24_i <= 16'sb0000000000110101;

in_29_25_r <= 16'sb0000000000110110;
in_29_25_i <= 16'sb0000000000110110;

in_29_26_r <= 16'sb0000000000110111;
in_29_26_i <= 16'sb0000000000110111;

in_29_27_r <= 16'sb0000000000111000;
in_29_27_i <= 16'sb0000000000111000;

in_29_28_r <= 16'sb0000000000111001;
in_29_28_i <= 16'sb0000000000111001;

in_29_29_r <= 16'sb0000000000111010;
in_29_29_i <= 16'sb0000000000111010;

in_29_30_r <= 16'sb0000000000111011;
in_29_30_i <= 16'sb0000000000111011;

in_29_31_r <= 16'sb0000000000111100;
in_29_31_i <= 16'sb0000000000111100;

in_29_32_r <= 16'sb0000000000111101;
in_29_32_i <= 16'sb0000000000111101;

in_30_1_r <= 16'sb0000000000011111;
in_30_1_i <= 16'sb0000000000011111;

in_30_2_r <= 16'sb0000000000100000;
in_30_2_i <= 16'sb0000000000100000;

in_30_3_r <= 16'sb0000000000100001;
in_30_3_i <= 16'sb0000000000100001;

in_30_4_r <= 16'sb0000000000100010;
in_30_4_i <= 16'sb0000000000100010;

in_30_5_r <= 16'sb0000000000100011;
in_30_5_i <= 16'sb0000000000100011;

in_30_6_r <= 16'sb0000000000100100;
in_30_6_i <= 16'sb0000000000100100;

in_30_7_r <= 16'sb0000000000100101;
in_30_7_i <= 16'sb0000000000100101;

in_30_8_r <= 16'sb0000000000100110;
in_30_8_i <= 16'sb0000000000100110;

in_30_9_r <= 16'sb0000000000100111;
in_30_9_i <= 16'sb0000000000100111;

in_30_10_r <= 16'sb0000000000101000;
in_30_10_i <= 16'sb0000000000101000;

in_30_11_r <= 16'sb0000000000101001;
in_30_11_i <= 16'sb0000000000101001;

in_30_12_r <= 16'sb0000000000101010;
in_30_12_i <= 16'sb0000000000101010;

in_30_13_r <= 16'sb0000000000101011;
in_30_13_i <= 16'sb0000000000101011;

in_30_14_r <= 16'sb0000000000101100;
in_30_14_i <= 16'sb0000000000101100;

in_30_15_r <= 16'sb0000000000101101;
in_30_15_i <= 16'sb0000000000101101;

in_30_16_r <= 16'sb0000000000101110;
in_30_16_i <= 16'sb0000000000101110;

in_30_17_r <= 16'sb0000000000101111;
in_30_17_i <= 16'sb0000000000101111;

in_30_18_r <= 16'sb0000000000110000;
in_30_18_i <= 16'sb0000000000110000;

in_30_19_r <= 16'sb0000000000110001;
in_30_19_i <= 16'sb0000000000110001;

in_30_20_r <= 16'sb0000000000110010;
in_30_20_i <= 16'sb0000000000110010;

in_30_21_r <= 16'sb0000000000110011;
in_30_21_i <= 16'sb0000000000110011;

in_30_22_r <= 16'sb0000000000110100;
in_30_22_i <= 16'sb0000000000110100;

in_30_23_r <= 16'sb0000000000110101;
in_30_23_i <= 16'sb0000000000110101;

in_30_24_r <= 16'sb0000000000110110;
in_30_24_i <= 16'sb0000000000110110;

in_30_25_r <= 16'sb0000000000110111;
in_30_25_i <= 16'sb0000000000110111;

in_30_26_r <= 16'sb0000000000111000;
in_30_26_i <= 16'sb0000000000111000;

in_30_27_r <= 16'sb0000000000111001;
in_30_27_i <= 16'sb0000000000111001;

in_30_28_r <= 16'sb0000000000111010;
in_30_28_i <= 16'sb0000000000111010;

in_30_29_r <= 16'sb0000000000111011;
in_30_29_i <= 16'sb0000000000111011;

in_30_30_r <= 16'sb0000000000111100;
in_30_30_i <= 16'sb0000000000111100;

in_30_31_r <= 16'sb0000000000111101;
in_30_31_i <= 16'sb0000000000111101;

in_30_32_r <= 16'sb0000000000111110;
in_30_32_i <= 16'sb0000000000111110;

in_31_1_r <= 16'sb0000000000100000;
in_31_1_i <= 16'sb0000000000100000;

in_31_2_r <= 16'sb0000000000100001;
in_31_2_i <= 16'sb0000000000100001;

in_31_3_r <= 16'sb0000000000100010;
in_31_3_i <= 16'sb0000000000100010;

in_31_4_r <= 16'sb0000000000100011;
in_31_4_i <= 16'sb0000000000100011;

in_31_5_r <= 16'sb0000000000100100;
in_31_5_i <= 16'sb0000000000100100;

in_31_6_r <= 16'sb0000000000100101;
in_31_6_i <= 16'sb0000000000100101;

in_31_7_r <= 16'sb0000000000100110;
in_31_7_i <= 16'sb0000000000100110;

in_31_8_r <= 16'sb0000000000100111;
in_31_8_i <= 16'sb0000000000100111;

in_31_9_r <= 16'sb0000000000101000;
in_31_9_i <= 16'sb0000000000101000;

in_31_10_r <= 16'sb0000000000101001;
in_31_10_i <= 16'sb0000000000101001;

in_31_11_r <= 16'sb0000000000101010;
in_31_11_i <= 16'sb0000000000101010;

in_31_12_r <= 16'sb0000000000101011;
in_31_12_i <= 16'sb0000000000101011;

in_31_13_r <= 16'sb0000000000101100;
in_31_13_i <= 16'sb0000000000101100;

in_31_14_r <= 16'sb0000000000101101;
in_31_14_i <= 16'sb0000000000101101;

in_31_15_r <= 16'sb0000000000101110;
in_31_15_i <= 16'sb0000000000101110;

in_31_16_r <= 16'sb0000000000101111;
in_31_16_i <= 16'sb0000000000101111;

in_31_17_r <= 16'sb0000000000110000;
in_31_17_i <= 16'sb0000000000110000;

in_31_18_r <= 16'sb0000000000110001;
in_31_18_i <= 16'sb0000000000110001;

in_31_19_r <= 16'sb0000000000110010;
in_31_19_i <= 16'sb0000000000110010;

in_31_20_r <= 16'sb0000000000110011;
in_31_20_i <= 16'sb0000000000110011;

in_31_21_r <= 16'sb0000000000110100;
in_31_21_i <= 16'sb0000000000110100;

in_31_22_r <= 16'sb0000000000110101;
in_31_22_i <= 16'sb0000000000110101;

in_31_23_r <= 16'sb0000000000110110;
in_31_23_i <= 16'sb0000000000110110;

in_31_24_r <= 16'sb0000000000110111;
in_31_24_i <= 16'sb0000000000110111;

in_31_25_r <= 16'sb0000000000111000;
in_31_25_i <= 16'sb0000000000111000;

in_31_26_r <= 16'sb0000000000111001;
in_31_26_i <= 16'sb0000000000111001;

in_31_27_r <= 16'sb0000000000111010;
in_31_27_i <= 16'sb0000000000111010;

in_31_28_r <= 16'sb0000000000111011;
in_31_28_i <= 16'sb0000000000111011;

in_31_29_r <= 16'sb0000000000111100;
in_31_29_i <= 16'sb0000000000111100;

in_31_30_r <= 16'sb0000000000111101;
in_31_30_i <= 16'sb0000000000111101;

in_31_31_r <= 16'sb0000000000111110;
in_31_31_i <= 16'sb0000000000111110;

in_31_32_r <= 16'sb0000000000111111;
in_31_32_i <= 16'sb0000000000111111;

in_32_1_r <= 16'sb0000000000100001;
in_32_1_i <= 16'sb0000000000100001;

in_32_2_r <= 16'sb0000000000100010;
in_32_2_i <= 16'sb0000000000100010;

in_32_3_r <= 16'sb0000000000100011;
in_32_3_i <= 16'sb0000000000100011;

in_32_4_r <= 16'sb0000000000100100;
in_32_4_i <= 16'sb0000000000100100;

in_32_5_r <= 16'sb0000000000100101;
in_32_5_i <= 16'sb0000000000100101;

in_32_6_r <= 16'sb0000000000100110;
in_32_6_i <= 16'sb0000000000100110;

in_32_7_r <= 16'sb0000000000100111;
in_32_7_i <= 16'sb0000000000100111;

in_32_8_r <= 16'sb0000000000101000;
in_32_8_i <= 16'sb0000000000101000;

in_32_9_r <= 16'sb0000000000101001;
in_32_9_i <= 16'sb0000000000101001;

in_32_10_r <= 16'sb0000000000101010;
in_32_10_i <= 16'sb0000000000101010;

in_32_11_r <= 16'sb0000000000101011;
in_32_11_i <= 16'sb0000000000101011;

in_32_12_r <= 16'sb0000000000101100;
in_32_12_i <= 16'sb0000000000101100;

in_32_13_r <= 16'sb0000000000101101;
in_32_13_i <= 16'sb0000000000101101;

in_32_14_r <= 16'sb0000000000101110;
in_32_14_i <= 16'sb0000000000101110;

in_32_15_r <= 16'sb0000000000101111;
in_32_15_i <= 16'sb0000000000101111;

in_32_16_r <= 16'sb0000000000110000;
in_32_16_i <= 16'sb0000000000110000;

in_32_17_r <= 16'sb0000000000110001;
in_32_17_i <= 16'sb0000000000110001;

in_32_18_r <= 16'sb0000000000110010;
in_32_18_i <= 16'sb0000000000110010;

in_32_19_r <= 16'sb0000000000110011;
in_32_19_i <= 16'sb0000000000110011;

in_32_20_r <= 16'sb0000000000110100;
in_32_20_i <= 16'sb0000000000110100;

in_32_21_r <= 16'sb0000000000110101;
in_32_21_i <= 16'sb0000000000110101;

in_32_22_r <= 16'sb0000000000110110;
in_32_22_i <= 16'sb0000000000110110;

in_32_23_r <= 16'sb0000000000110111;
in_32_23_i <= 16'sb0000000000110111;

in_32_24_r <= 16'sb0000000000111000;
in_32_24_i <= 16'sb0000000000111000;

in_32_25_r <= 16'sb0000000000111001;
in_32_25_i <= 16'sb0000000000111001;

in_32_26_r <= 16'sb0000000000111010;
in_32_26_i <= 16'sb0000000000111010;

in_32_27_r <= 16'sb0000000000111011;
in_32_27_i <= 16'sb0000000000111011;

in_32_28_r <= 16'sb0000000000111100;
in_32_28_i <= 16'sb0000000000111100;

in_32_29_r <= 16'sb0000000000111101;
in_32_29_i <= 16'sb0000000000111101;

in_32_30_r <= 16'sb0000000000111110;
in_32_30_i <= 16'sb0000000000111110;

in_32_31_r <= 16'sb0000000000111111;
in_32_31_i <= 16'sb0000000000111111;

in_32_32_r <= 16'sb0000000001000000;
in_32_32_i <= 16'sb0000000001000000;


#500
$finish;

end


always #5 begin
            clk <= ~clk;
        end
        
        
endmodule
