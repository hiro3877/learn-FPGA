`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/05/31 16:18:23
// Design Name: 
// Module Name: top_sim
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module top_sim();

    reg d_in_;              //����񂯂�I������M��
    reg gtp_;               //�O�[�`���L�p�[���͂���M��
    reg pon;                //����񂯂�ۂ�I
    wire [`L_DataBus] led_;   //�\���p7segLED
    
    
    top top1 (d_in_,gtp_,pon,led_);
    
    
    initial begin
        d_in_ <= 1'b1;
        gtp_  <= 1'b1;
        pon   <= 1'b0;
        
    #20
        gtp_ <= 1'b0;
    
    #20
        gtp_ <= 1'b1;       //������
                
    /********************************/
        
    #20
        d_in_ <= 1'b0;      //�O�[
    
    #20
        d_in_ <= 1'b1; 

    #20
        d_in_ <= 1'b0;      //�`���L
    
    #20
        d_in_ <= 1'b1; 
        
    #20
        d_in_ <= 1'b0;      //�p�[
        
    #20
        d_in_ <= 1'b1; 

    #20
        d_in_ <= 1'b0;      //�O�[
        
    #20
        d_in_ <= 1'b1; 
        
    /*************************/
    
    #20
        gtp_ <= 1'b0;       //�O�[����
        
    #20
        gtp_ <= 1'b1;       //�O�[����
                    
        
    /*************************/
        
        
    #20
        d_in_ <= 1'b0;      //�O�[
        
    #20
        d_in_ <= 1'b1; 
    
    #20
        d_in_ <= 1'b0;      //�`���L
        
    #20
        d_in_ <= 1'b1; 
        
    /*************************/
    
    #20
        gtp_ <= 1'b0;       //�`���L����
    
    #20
        gtp_ <= 1'b1;       //�`���L����
                
        
    /**************************/
    
    #20
        d_in_ <= 1'b0;      //�O�[
    
    #20
        d_in_ <= 1'b1; 

    #20
        d_in_ <= 1'b0;      //�`���L
    
    #20
        d_in_ <= 1'b1; 
        
    #20
        d_in_ <= 1'b0;      //�p�[
        
    #20
        d_in_ <= 1'b1; 

    /*************************/
    
    #20
        gtp_ <= 1'b0;       //�p�[����
  
    #20
        gtp_ <= 1'b1;       //�p�[����
                    
    /*************************/
    
    #20
        pon <= 1'b1;        //����񂯂�ۂ�I
    
    /************************/
    
    #20
        $finish;
    end
    
        
    

endmodule
