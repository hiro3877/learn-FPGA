`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/08/20 20:43:41
// Design Name: 
// Module Name: top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
/////////////////////////////////////////////////////////////////////////////////

`include "./nettype.h"
`include "./std_define.h"

module top_io(
input wire clk,
input wire signed [`InBus]		in_r,
input wire signed [`InBus]		in_i,
output wire signed [`OutBus]		out_r,
output wire signed [`OutBus]		out_i

);

wire signed [`InBus]		in_1_1_r;
wire signed [`InBus]		in_1_1_i;
wire signed [`InBus]		in_1_2_r;
wire signed [`InBus]		in_1_2_i;
wire signed [`InBus]		in_1_3_r;
wire signed [`InBus]		in_1_3_i;
wire signed [`InBus]		in_1_4_r;
wire signed [`InBus]		in_1_4_i;
wire signed [`InBus]		in_1_5_r;
wire signed [`InBus]		in_1_5_i;
wire signed [`InBus]		in_1_6_r;
wire signed [`InBus]		in_1_6_i;
wire signed [`InBus]		in_1_7_r;
wire signed [`InBus]		in_1_7_i;
wire signed [`InBus]		in_1_8_r;
wire signed [`InBus]		in_1_8_i;
wire signed [`InBus]		in_1_9_r;
wire signed [`InBus]		in_1_9_i;
wire signed [`InBus]		in_1_10_r;
wire signed [`InBus]		in_1_10_i;
wire signed [`InBus]		in_1_11_r;
wire signed [`InBus]		in_1_11_i;
wire signed [`InBus]		in_1_12_r;
wire signed [`InBus]		in_1_12_i;
wire signed [`InBus]		in_1_13_r;
wire signed [`InBus]		in_1_13_i;
wire signed [`InBus]		in_1_14_r;
wire signed [`InBus]		in_1_14_i;
wire signed [`InBus]		in_1_15_r;
wire signed [`InBus]		in_1_15_i;
wire signed [`InBus]		in_1_16_r;
wire signed [`InBus]		in_1_16_i;
wire signed [`InBus]		in_2_1_r;
wire signed [`InBus]		in_2_1_i;
wire signed [`InBus]		in_2_2_r;
wire signed [`InBus]		in_2_2_i;
wire signed [`InBus]		in_2_3_r;
wire signed [`InBus]		in_2_3_i;
wire signed [`InBus]		in_2_4_r;
wire signed [`InBus]		in_2_4_i;
wire signed [`InBus]		in_2_5_r;
wire signed [`InBus]		in_2_5_i;
wire signed [`InBus]		in_2_6_r;
wire signed [`InBus]		in_2_6_i;
wire signed [`InBus]		in_2_7_r;
wire signed [`InBus]		in_2_7_i;
wire signed [`InBus]		in_2_8_r;
wire signed [`InBus]		in_2_8_i;
wire signed [`InBus]		in_2_9_r;
wire signed [`InBus]		in_2_9_i;
wire signed [`InBus]		in_2_10_r;
wire signed [`InBus]		in_2_10_i;
wire signed [`InBus]		in_2_11_r;
wire signed [`InBus]		in_2_11_i;
wire signed [`InBus]		in_2_12_r;
wire signed [`InBus]		in_2_12_i;
wire signed [`InBus]		in_2_13_r;
wire signed [`InBus]		in_2_13_i;
wire signed [`InBus]		in_2_14_r;
wire signed [`InBus]		in_2_14_i;
wire signed [`InBus]		in_2_15_r;
wire signed [`InBus]		in_2_15_i;
wire signed [`InBus]		in_2_16_r;
wire signed [`InBus]		in_2_16_i;
wire signed [`InBus]		in_3_1_r;
wire signed [`InBus]		in_3_1_i;
wire signed [`InBus]		in_3_2_r;
wire signed [`InBus]		in_3_2_i;
wire signed [`InBus]		in_3_3_r;
wire signed [`InBus]		in_3_3_i;
wire signed [`InBus]		in_3_4_r;
wire signed [`InBus]		in_3_4_i;
wire signed [`InBus]		in_3_5_r;
wire signed [`InBus]		in_3_5_i;
wire signed [`InBus]		in_3_6_r;
wire signed [`InBus]		in_3_6_i;
wire signed [`InBus]		in_3_7_r;
wire signed [`InBus]		in_3_7_i;
wire signed [`InBus]		in_3_8_r;
wire signed [`InBus]		in_3_8_i;
wire signed [`InBus]		in_3_9_r;
wire signed [`InBus]		in_3_9_i;
wire signed [`InBus]		in_3_10_r;
wire signed [`InBus]		in_3_10_i;
wire signed [`InBus]		in_3_11_r;
wire signed [`InBus]		in_3_11_i;
wire signed [`InBus]		in_3_12_r;
wire signed [`InBus]		in_3_12_i;
wire signed [`InBus]		in_3_13_r;
wire signed [`InBus]		in_3_13_i;
wire signed [`InBus]		in_3_14_r;
wire signed [`InBus]		in_3_14_i;
wire signed [`InBus]		in_3_15_r;
wire signed [`InBus]		in_3_15_i;
wire signed [`InBus]		in_3_16_r;
wire signed [`InBus]		in_3_16_i;
wire signed [`InBus]		in_4_1_r;
wire signed [`InBus]		in_4_1_i;
wire signed [`InBus]		in_4_2_r;
wire signed [`InBus]		in_4_2_i;
wire signed [`InBus]		in_4_3_r;
wire signed [`InBus]		in_4_3_i;
wire signed [`InBus]		in_4_4_r;
wire signed [`InBus]		in_4_4_i;
wire signed [`InBus]		in_4_5_r;
wire signed [`InBus]		in_4_5_i;
wire signed [`InBus]		in_4_6_r;
wire signed [`InBus]		in_4_6_i;
wire signed [`InBus]		in_4_7_r;
wire signed [`InBus]		in_4_7_i;
wire signed [`InBus]		in_4_8_r;
wire signed [`InBus]		in_4_8_i;
wire signed [`InBus]		in_4_9_r;
wire signed [`InBus]		in_4_9_i;
wire signed [`InBus]		in_4_10_r;
wire signed [`InBus]		in_4_10_i;
wire signed [`InBus]		in_4_11_r;
wire signed [`InBus]		in_4_11_i;
wire signed [`InBus]		in_4_12_r;
wire signed [`InBus]		in_4_12_i;
wire signed [`InBus]		in_4_13_r;
wire signed [`InBus]		in_4_13_i;
wire signed [`InBus]		in_4_14_r;
wire signed [`InBus]		in_4_14_i;
wire signed [`InBus]		in_4_15_r;
wire signed [`InBus]		in_4_15_i;
wire signed [`InBus]		in_4_16_r;
wire signed [`InBus]		in_4_16_i;
wire signed [`InBus]		in_5_1_r;
wire signed [`InBus]		in_5_1_i;
wire signed [`InBus]		in_5_2_r;
wire signed [`InBus]		in_5_2_i;
wire signed [`InBus]		in_5_3_r;
wire signed [`InBus]		in_5_3_i;
wire signed [`InBus]		in_5_4_r;
wire signed [`InBus]		in_5_4_i;
wire signed [`InBus]		in_5_5_r;
wire signed [`InBus]		in_5_5_i;
wire signed [`InBus]		in_5_6_r;
wire signed [`InBus]		in_5_6_i;
wire signed [`InBus]		in_5_7_r;
wire signed [`InBus]		in_5_7_i;
wire signed [`InBus]		in_5_8_r;
wire signed [`InBus]		in_5_8_i;
wire signed [`InBus]		in_5_9_r;
wire signed [`InBus]		in_5_9_i;
wire signed [`InBus]		in_5_10_r;
wire signed [`InBus]		in_5_10_i;
wire signed [`InBus]		in_5_11_r;
wire signed [`InBus]		in_5_11_i;
wire signed [`InBus]		in_5_12_r;
wire signed [`InBus]		in_5_12_i;
wire signed [`InBus]		in_5_13_r;
wire signed [`InBus]		in_5_13_i;
wire signed [`InBus]		in_5_14_r;
wire signed [`InBus]		in_5_14_i;
wire signed [`InBus]		in_5_15_r;
wire signed [`InBus]		in_5_15_i;
wire signed [`InBus]		in_5_16_r;
wire signed [`InBus]		in_5_16_i;
wire signed [`InBus]		in_6_1_r;
wire signed [`InBus]		in_6_1_i;
wire signed [`InBus]		in_6_2_r;
wire signed [`InBus]		in_6_2_i;
wire signed [`InBus]		in_6_3_r;
wire signed [`InBus]		in_6_3_i;
wire signed [`InBus]		in_6_4_r;
wire signed [`InBus]		in_6_4_i;
wire signed [`InBus]		in_6_5_r;
wire signed [`InBus]		in_6_5_i;
wire signed [`InBus]		in_6_6_r;
wire signed [`InBus]		in_6_6_i;
wire signed [`InBus]		in_6_7_r;
wire signed [`InBus]		in_6_7_i;
wire signed [`InBus]		in_6_8_r;
wire signed [`InBus]		in_6_8_i;
wire signed [`InBus]		in_6_9_r;
wire signed [`InBus]		in_6_9_i;
wire signed [`InBus]		in_6_10_r;
wire signed [`InBus]		in_6_10_i;
wire signed [`InBus]		in_6_11_r;
wire signed [`InBus]		in_6_11_i;
wire signed [`InBus]		in_6_12_r;
wire signed [`InBus]		in_6_12_i;
wire signed [`InBus]		in_6_13_r;
wire signed [`InBus]		in_6_13_i;
wire signed [`InBus]		in_6_14_r;
wire signed [`InBus]		in_6_14_i;
wire signed [`InBus]		in_6_15_r;
wire signed [`InBus]		in_6_15_i;
wire signed [`InBus]		in_6_16_r;
wire signed [`InBus]		in_6_16_i;
wire signed [`InBus]		in_7_1_r;
wire signed [`InBus]		in_7_1_i;
wire signed [`InBus]		in_7_2_r;
wire signed [`InBus]		in_7_2_i;
wire signed [`InBus]		in_7_3_r;
wire signed [`InBus]		in_7_3_i;
wire signed [`InBus]		in_7_4_r;
wire signed [`InBus]		in_7_4_i;
wire signed [`InBus]		in_7_5_r;
wire signed [`InBus]		in_7_5_i;
wire signed [`InBus]		in_7_6_r;
wire signed [`InBus]		in_7_6_i;
wire signed [`InBus]		in_7_7_r;
wire signed [`InBus]		in_7_7_i;
wire signed [`InBus]		in_7_8_r;
wire signed [`InBus]		in_7_8_i;
wire signed [`InBus]		in_7_9_r;
wire signed [`InBus]		in_7_9_i;
wire signed [`InBus]		in_7_10_r;
wire signed [`InBus]		in_7_10_i;
wire signed [`InBus]		in_7_11_r;
wire signed [`InBus]		in_7_11_i;
wire signed [`InBus]		in_7_12_r;
wire signed [`InBus]		in_7_12_i;
wire signed [`InBus]		in_7_13_r;
wire signed [`InBus]		in_7_13_i;
wire signed [`InBus]		in_7_14_r;
wire signed [`InBus]		in_7_14_i;
wire signed [`InBus]		in_7_15_r;
wire signed [`InBus]		in_7_15_i;
wire signed [`InBus]		in_7_16_r;
wire signed [`InBus]		in_7_16_i;
wire signed [`InBus]		in_8_1_r;
wire signed [`InBus]		in_8_1_i;
wire signed [`InBus]		in_8_2_r;
wire signed [`InBus]		in_8_2_i;
wire signed [`InBus]		in_8_3_r;
wire signed [`InBus]		in_8_3_i;
wire signed [`InBus]		in_8_4_r;
wire signed [`InBus]		in_8_4_i;
wire signed [`InBus]		in_8_5_r;
wire signed [`InBus]		in_8_5_i;
wire signed [`InBus]		in_8_6_r;
wire signed [`InBus]		in_8_6_i;
wire signed [`InBus]		in_8_7_r;
wire signed [`InBus]		in_8_7_i;
wire signed [`InBus]		in_8_8_r;
wire signed [`InBus]		in_8_8_i;
wire signed [`InBus]		in_8_9_r;
wire signed [`InBus]		in_8_9_i;
wire signed [`InBus]		in_8_10_r;
wire signed [`InBus]		in_8_10_i;
wire signed [`InBus]		in_8_11_r;
wire signed [`InBus]		in_8_11_i;
wire signed [`InBus]		in_8_12_r;
wire signed [`InBus]		in_8_12_i;
wire signed [`InBus]		in_8_13_r;
wire signed [`InBus]		in_8_13_i;
wire signed [`InBus]		in_8_14_r;
wire signed [`InBus]		in_8_14_i;
wire signed [`InBus]		in_8_15_r;
wire signed [`InBus]		in_8_15_i;
wire signed [`InBus]		in_8_16_r;
wire signed [`InBus]		in_8_16_i;
wire signed [`InBus]		in_9_1_r;
wire signed [`InBus]		in_9_1_i;
wire signed [`InBus]		in_9_2_r;
wire signed [`InBus]		in_9_2_i;
wire signed [`InBus]		in_9_3_r;
wire signed [`InBus]		in_9_3_i;
wire signed [`InBus]		in_9_4_r;
wire signed [`InBus]		in_9_4_i;
wire signed [`InBus]		in_9_5_r;
wire signed [`InBus]		in_9_5_i;
wire signed [`InBus]		in_9_6_r;
wire signed [`InBus]		in_9_6_i;
wire signed [`InBus]		in_9_7_r;
wire signed [`InBus]		in_9_7_i;
wire signed [`InBus]		in_9_8_r;
wire signed [`InBus]		in_9_8_i;
wire signed [`InBus]		in_9_9_r;
wire signed [`InBus]		in_9_9_i;
wire signed [`InBus]		in_9_10_r;
wire signed [`InBus]		in_9_10_i;
wire signed [`InBus]		in_9_11_r;
wire signed [`InBus]		in_9_11_i;
wire signed [`InBus]		in_9_12_r;
wire signed [`InBus]		in_9_12_i;
wire signed [`InBus]		in_9_13_r;
wire signed [`InBus]		in_9_13_i;
wire signed [`InBus]		in_9_14_r;
wire signed [`InBus]		in_9_14_i;
wire signed [`InBus]		in_9_15_r;
wire signed [`InBus]		in_9_15_i;
wire signed [`InBus]		in_9_16_r;
wire signed [`InBus]		in_9_16_i;
wire signed [`InBus]		in_10_1_r;
wire signed [`InBus]		in_10_1_i;
wire signed [`InBus]		in_10_2_r;
wire signed [`InBus]		in_10_2_i;
wire signed [`InBus]		in_10_3_r;
wire signed [`InBus]		in_10_3_i;
wire signed [`InBus]		in_10_4_r;
wire signed [`InBus]		in_10_4_i;
wire signed [`InBus]		in_10_5_r;
wire signed [`InBus]		in_10_5_i;
wire signed [`InBus]		in_10_6_r;
wire signed [`InBus]		in_10_6_i;
wire signed [`InBus]		in_10_7_r;
wire signed [`InBus]		in_10_7_i;
wire signed [`InBus]		in_10_8_r;
wire signed [`InBus]		in_10_8_i;
wire signed [`InBus]		in_10_9_r;
wire signed [`InBus]		in_10_9_i;
wire signed [`InBus]		in_10_10_r;
wire signed [`InBus]		in_10_10_i;
wire signed [`InBus]		in_10_11_r;
wire signed [`InBus]		in_10_11_i;
wire signed [`InBus]		in_10_12_r;
wire signed [`InBus]		in_10_12_i;
wire signed [`InBus]		in_10_13_r;
wire signed [`InBus]		in_10_13_i;
wire signed [`InBus]		in_10_14_r;
wire signed [`InBus]		in_10_14_i;
wire signed [`InBus]		in_10_15_r;
wire signed [`InBus]		in_10_15_i;
wire signed [`InBus]		in_10_16_r;
wire signed [`InBus]		in_10_16_i;
wire signed [`InBus]		in_11_1_r;
wire signed [`InBus]		in_11_1_i;
wire signed [`InBus]		in_11_2_r;
wire signed [`InBus]		in_11_2_i;
wire signed [`InBus]		in_11_3_r;
wire signed [`InBus]		in_11_3_i;
wire signed [`InBus]		in_11_4_r;
wire signed [`InBus]		in_11_4_i;
wire signed [`InBus]		in_11_5_r;
wire signed [`InBus]		in_11_5_i;
wire signed [`InBus]		in_11_6_r;
wire signed [`InBus]		in_11_6_i;
wire signed [`InBus]		in_11_7_r;
wire signed [`InBus]		in_11_7_i;
wire signed [`InBus]		in_11_8_r;
wire signed [`InBus]		in_11_8_i;
wire signed [`InBus]		in_11_9_r;
wire signed [`InBus]		in_11_9_i;
wire signed [`InBus]		in_11_10_r;
wire signed [`InBus]		in_11_10_i;
wire signed [`InBus]		in_11_11_r;
wire signed [`InBus]		in_11_11_i;
wire signed [`InBus]		in_11_12_r;
wire signed [`InBus]		in_11_12_i;
wire signed [`InBus]		in_11_13_r;
wire signed [`InBus]		in_11_13_i;
wire signed [`InBus]		in_11_14_r;
wire signed [`InBus]		in_11_14_i;
wire signed [`InBus]		in_11_15_r;
wire signed [`InBus]		in_11_15_i;
wire signed [`InBus]		in_11_16_r;
wire signed [`InBus]		in_11_16_i;
wire signed [`InBus]		in_12_1_r;
wire signed [`InBus]		in_12_1_i;
wire signed [`InBus]		in_12_2_r;
wire signed [`InBus]		in_12_2_i;
wire signed [`InBus]		in_12_3_r;
wire signed [`InBus]		in_12_3_i;
wire signed [`InBus]		in_12_4_r;
wire signed [`InBus]		in_12_4_i;
wire signed [`InBus]		in_12_5_r;
wire signed [`InBus]		in_12_5_i;
wire signed [`InBus]		in_12_6_r;
wire signed [`InBus]		in_12_6_i;
wire signed [`InBus]		in_12_7_r;
wire signed [`InBus]		in_12_7_i;
wire signed [`InBus]		in_12_8_r;
wire signed [`InBus]		in_12_8_i;
wire signed [`InBus]		in_12_9_r;
wire signed [`InBus]		in_12_9_i;
wire signed [`InBus]		in_12_10_r;
wire signed [`InBus]		in_12_10_i;
wire signed [`InBus]		in_12_11_r;
wire signed [`InBus]		in_12_11_i;
wire signed [`InBus]		in_12_12_r;
wire signed [`InBus]		in_12_12_i;
wire signed [`InBus]		in_12_13_r;
wire signed [`InBus]		in_12_13_i;
wire signed [`InBus]		in_12_14_r;
wire signed [`InBus]		in_12_14_i;
wire signed [`InBus]		in_12_15_r;
wire signed [`InBus]		in_12_15_i;
wire signed [`InBus]		in_12_16_r;
wire signed [`InBus]		in_12_16_i;
wire signed [`InBus]		in_13_1_r;
wire signed [`InBus]		in_13_1_i;
wire signed [`InBus]		in_13_2_r;
wire signed [`InBus]		in_13_2_i;
wire signed [`InBus]		in_13_3_r;
wire signed [`InBus]		in_13_3_i;
wire signed [`InBus]		in_13_4_r;
wire signed [`InBus]		in_13_4_i;
wire signed [`InBus]		in_13_5_r;
wire signed [`InBus]		in_13_5_i;
wire signed [`InBus]		in_13_6_r;
wire signed [`InBus]		in_13_6_i;
wire signed [`InBus]		in_13_7_r;
wire signed [`InBus]		in_13_7_i;
wire signed [`InBus]		in_13_8_r;
wire signed [`InBus]		in_13_8_i;
wire signed [`InBus]		in_13_9_r;
wire signed [`InBus]		in_13_9_i;
wire signed [`InBus]		in_13_10_r;
wire signed [`InBus]		in_13_10_i;
wire signed [`InBus]		in_13_11_r;
wire signed [`InBus]		in_13_11_i;
wire signed [`InBus]		in_13_12_r;
wire signed [`InBus]		in_13_12_i;
wire signed [`InBus]		in_13_13_r;
wire signed [`InBus]		in_13_13_i;
wire signed [`InBus]		in_13_14_r;
wire signed [`InBus]		in_13_14_i;
wire signed [`InBus]		in_13_15_r;
wire signed [`InBus]		in_13_15_i;
wire signed [`InBus]		in_13_16_r;
wire signed [`InBus]		in_13_16_i;
wire signed [`InBus]		in_14_1_r;
wire signed [`InBus]		in_14_1_i;
wire signed [`InBus]		in_14_2_r;
wire signed [`InBus]		in_14_2_i;
wire signed [`InBus]		in_14_3_r;
wire signed [`InBus]		in_14_3_i;
wire signed [`InBus]		in_14_4_r;
wire signed [`InBus]		in_14_4_i;
wire signed [`InBus]		in_14_5_r;
wire signed [`InBus]		in_14_5_i;
wire signed [`InBus]		in_14_6_r;
wire signed [`InBus]		in_14_6_i;
wire signed [`InBus]		in_14_7_r;
wire signed [`InBus]		in_14_7_i;
wire signed [`InBus]		in_14_8_r;
wire signed [`InBus]		in_14_8_i;
wire signed [`InBus]		in_14_9_r;
wire signed [`InBus]		in_14_9_i;
wire signed [`InBus]		in_14_10_r;
wire signed [`InBus]		in_14_10_i;
wire signed [`InBus]		in_14_11_r;
wire signed [`InBus]		in_14_11_i;
wire signed [`InBus]		in_14_12_r;
wire signed [`InBus]		in_14_12_i;
wire signed [`InBus]		in_14_13_r;
wire signed [`InBus]		in_14_13_i;
wire signed [`InBus]		in_14_14_r;
wire signed [`InBus]		in_14_14_i;
wire signed [`InBus]		in_14_15_r;
wire signed [`InBus]		in_14_15_i;
wire signed [`InBus]		in_14_16_r;
wire signed [`InBus]		in_14_16_i;
wire signed [`InBus]		in_15_1_r;
wire signed [`InBus]		in_15_1_i;
wire signed [`InBus]		in_15_2_r;
wire signed [`InBus]		in_15_2_i;
wire signed [`InBus]		in_15_3_r;
wire signed [`InBus]		in_15_3_i;
wire signed [`InBus]		in_15_4_r;
wire signed [`InBus]		in_15_4_i;
wire signed [`InBus]		in_15_5_r;
wire signed [`InBus]		in_15_5_i;
wire signed [`InBus]		in_15_6_r;
wire signed [`InBus]		in_15_6_i;
wire signed [`InBus]		in_15_7_r;
wire signed [`InBus]		in_15_7_i;
wire signed [`InBus]		in_15_8_r;
wire signed [`InBus]		in_15_8_i;
wire signed [`InBus]		in_15_9_r;
wire signed [`InBus]		in_15_9_i;
wire signed [`InBus]		in_15_10_r;
wire signed [`InBus]		in_15_10_i;
wire signed [`InBus]		in_15_11_r;
wire signed [`InBus]		in_15_11_i;
wire signed [`InBus]		in_15_12_r;
wire signed [`InBus]		in_15_12_i;
wire signed [`InBus]		in_15_13_r;
wire signed [`InBus]		in_15_13_i;
wire signed [`InBus]		in_15_14_r;
wire signed [`InBus]		in_15_14_i;
wire signed [`InBus]		in_15_15_r;
wire signed [`InBus]		in_15_15_i;
wire signed [`InBus]		in_15_16_r;
wire signed [`InBus]		in_15_16_i;
wire signed [`InBus]		in_16_1_r;
wire signed [`InBus]		in_16_1_i;
wire signed [`InBus]		in_16_2_r;
wire signed [`InBus]		in_16_2_i;
wire signed [`InBus]		in_16_3_r;
wire signed [`InBus]		in_16_3_i;
wire signed [`InBus]		in_16_4_r;
wire signed [`InBus]		in_16_4_i;
wire signed [`InBus]		in_16_5_r;
wire signed [`InBus]		in_16_5_i;
wire signed [`InBus]		in_16_6_r;
wire signed [`InBus]		in_16_6_i;
wire signed [`InBus]		in_16_7_r;
wire signed [`InBus]		in_16_7_i;
wire signed [`InBus]		in_16_8_r;
wire signed [`InBus]		in_16_8_i;
wire signed [`InBus]		in_16_9_r;
wire signed [`InBus]		in_16_9_i;
wire signed [`InBus]		in_16_10_r;
wire signed [`InBus]		in_16_10_i;
wire signed [`InBus]		in_16_11_r;
wire signed [`InBus]		in_16_11_i;
wire signed [`InBus]		in_16_12_r;
wire signed [`InBus]		in_16_12_i;
wire signed [`InBus]		in_16_13_r;
wire signed [`InBus]		in_16_13_i;
wire signed [`InBus]		in_16_14_r;
wire signed [`InBus]		in_16_14_i;
wire signed [`InBus]		in_16_15_r;
wire signed [`InBus]		in_16_15_i;
wire signed [`InBus]		in_16_16_r;
wire signed [`InBus]		in_16_16_i;

wire signed [`OutBus]		out_1_1_r;
wire signed [`OutBus]		out_1_1_i;
wire signed [`OutBus]		out_1_2_r;
wire signed [`OutBus]		out_1_2_i;
wire signed [`OutBus]		out_1_3_r;
wire signed [`OutBus]		out_1_3_i;
wire signed [`OutBus]		out_1_4_r;
wire signed [`OutBus]		out_1_4_i;
wire signed [`OutBus]		out_1_5_r;
wire signed [`OutBus]		out_1_5_i;
wire signed [`OutBus]		out_1_6_r;
wire signed [`OutBus]		out_1_6_i;
wire signed [`OutBus]		out_1_7_r;
wire signed [`OutBus]		out_1_7_i;
wire signed [`OutBus]		out_1_8_r;
wire signed [`OutBus]		out_1_8_i;
wire signed [`OutBus]		out_1_9_r;
wire signed [`OutBus]		out_1_9_i;
wire signed [`OutBus]		out_1_10_r;
wire signed [`OutBus]		out_1_10_i;
wire signed [`OutBus]		out_1_11_r;
wire signed [`OutBus]		out_1_11_i;
wire signed [`OutBus]		out_1_12_r;
wire signed [`OutBus]		out_1_12_i;
wire signed [`OutBus]		out_1_13_r;
wire signed [`OutBus]		out_1_13_i;
wire signed [`OutBus]		out_1_14_r;
wire signed [`OutBus]		out_1_14_i;
wire signed [`OutBus]		out_1_15_r;
wire signed [`OutBus]		out_1_15_i;
wire signed [`OutBus]		out_1_16_r;
wire signed [`OutBus]		out_1_16_i;
wire signed [`OutBus]		out_2_1_r;
wire signed [`OutBus]		out_2_1_i;
wire signed [`OutBus]		out_2_2_r;
wire signed [`OutBus]		out_2_2_i;
wire signed [`OutBus]		out_2_3_r;
wire signed [`OutBus]		out_2_3_i;
wire signed [`OutBus]		out_2_4_r;
wire signed [`OutBus]		out_2_4_i;
wire signed [`OutBus]		out_2_5_r;
wire signed [`OutBus]		out_2_5_i;
wire signed [`OutBus]		out_2_6_r;
wire signed [`OutBus]		out_2_6_i;
wire signed [`OutBus]		out_2_7_r;
wire signed [`OutBus]		out_2_7_i;
wire signed [`OutBus]		out_2_8_r;
wire signed [`OutBus]		out_2_8_i;
wire signed [`OutBus]		out_2_9_r;
wire signed [`OutBus]		out_2_9_i;
wire signed [`OutBus]		out_2_10_r;
wire signed [`OutBus]		out_2_10_i;
wire signed [`OutBus]		out_2_11_r;
wire signed [`OutBus]		out_2_11_i;
wire signed [`OutBus]		out_2_12_r;
wire signed [`OutBus]		out_2_12_i;
wire signed [`OutBus]		out_2_13_r;
wire signed [`OutBus]		out_2_13_i;
wire signed [`OutBus]		out_2_14_r;
wire signed [`OutBus]		out_2_14_i;
wire signed [`OutBus]		out_2_15_r;
wire signed [`OutBus]		out_2_15_i;
wire signed [`OutBus]		out_2_16_r;
wire signed [`OutBus]		out_2_16_i;
wire signed [`OutBus]		out_3_1_r;
wire signed [`OutBus]		out_3_1_i;
wire signed [`OutBus]		out_3_2_r;
wire signed [`OutBus]		out_3_2_i;
wire signed [`OutBus]		out_3_3_r;
wire signed [`OutBus]		out_3_3_i;
wire signed [`OutBus]		out_3_4_r;
wire signed [`OutBus]		out_3_4_i;
wire signed [`OutBus]		out_3_5_r;
wire signed [`OutBus]		out_3_5_i;
wire signed [`OutBus]		out_3_6_r;
wire signed [`OutBus]		out_3_6_i;
wire signed [`OutBus]		out_3_7_r;
wire signed [`OutBus]		out_3_7_i;
wire signed [`OutBus]		out_3_8_r;
wire signed [`OutBus]		out_3_8_i;
wire signed [`OutBus]		out_3_9_r;
wire signed [`OutBus]		out_3_9_i;
wire signed [`OutBus]		out_3_10_r;
wire signed [`OutBus]		out_3_10_i;
wire signed [`OutBus]		out_3_11_r;
wire signed [`OutBus]		out_3_11_i;
wire signed [`OutBus]		out_3_12_r;
wire signed [`OutBus]		out_3_12_i;
wire signed [`OutBus]		out_3_13_r;
wire signed [`OutBus]		out_3_13_i;
wire signed [`OutBus]		out_3_14_r;
wire signed [`OutBus]		out_3_14_i;
wire signed [`OutBus]		out_3_15_r;
wire signed [`OutBus]		out_3_15_i;
wire signed [`OutBus]		out_3_16_r;
wire signed [`OutBus]		out_3_16_i;
wire signed [`OutBus]		out_4_1_r;
wire signed [`OutBus]		out_4_1_i;
wire signed [`OutBus]		out_4_2_r;
wire signed [`OutBus]		out_4_2_i;
wire signed [`OutBus]		out_4_3_r;
wire signed [`OutBus]		out_4_3_i;
wire signed [`OutBus]		out_4_4_r;
wire signed [`OutBus]		out_4_4_i;
wire signed [`OutBus]		out_4_5_r;
wire signed [`OutBus]		out_4_5_i;
wire signed [`OutBus]		out_4_6_r;
wire signed [`OutBus]		out_4_6_i;
wire signed [`OutBus]		out_4_7_r;
wire signed [`OutBus]		out_4_7_i;
wire signed [`OutBus]		out_4_8_r;
wire signed [`OutBus]		out_4_8_i;
wire signed [`OutBus]		out_4_9_r;
wire signed [`OutBus]		out_4_9_i;
wire signed [`OutBus]		out_4_10_r;
wire signed [`OutBus]		out_4_10_i;
wire signed [`OutBus]		out_4_11_r;
wire signed [`OutBus]		out_4_11_i;
wire signed [`OutBus]		out_4_12_r;
wire signed [`OutBus]		out_4_12_i;
wire signed [`OutBus]		out_4_13_r;
wire signed [`OutBus]		out_4_13_i;
wire signed [`OutBus]		out_4_14_r;
wire signed [`OutBus]		out_4_14_i;
wire signed [`OutBus]		out_4_15_r;
wire signed [`OutBus]		out_4_15_i;
wire signed [`OutBus]		out_4_16_r;
wire signed [`OutBus]		out_4_16_i;
wire signed [`OutBus]		out_5_1_r;
wire signed [`OutBus]		out_5_1_i;
wire signed [`OutBus]		out_5_2_r;
wire signed [`OutBus]		out_5_2_i;
wire signed [`OutBus]		out_5_3_r;
wire signed [`OutBus]		out_5_3_i;
wire signed [`OutBus]		out_5_4_r;
wire signed [`OutBus]		out_5_4_i;
wire signed [`OutBus]		out_5_5_r;
wire signed [`OutBus]		out_5_5_i;
wire signed [`OutBus]		out_5_6_r;
wire signed [`OutBus]		out_5_6_i;
wire signed [`OutBus]		out_5_7_r;
wire signed [`OutBus]		out_5_7_i;
wire signed [`OutBus]		out_5_8_r;
wire signed [`OutBus]		out_5_8_i;
wire signed [`OutBus]		out_5_9_r;
wire signed [`OutBus]		out_5_9_i;
wire signed [`OutBus]		out_5_10_r;
wire signed [`OutBus]		out_5_10_i;
wire signed [`OutBus]		out_5_11_r;
wire signed [`OutBus]		out_5_11_i;
wire signed [`OutBus]		out_5_12_r;
wire signed [`OutBus]		out_5_12_i;
wire signed [`OutBus]		out_5_13_r;
wire signed [`OutBus]		out_5_13_i;
wire signed [`OutBus]		out_5_14_r;
wire signed [`OutBus]		out_5_14_i;
wire signed [`OutBus]		out_5_15_r;
wire signed [`OutBus]		out_5_15_i;
wire signed [`OutBus]		out_5_16_r;
wire signed [`OutBus]		out_5_16_i;
wire signed [`OutBus]		out_6_1_r;
wire signed [`OutBus]		out_6_1_i;
wire signed [`OutBus]		out_6_2_r;
wire signed [`OutBus]		out_6_2_i;
wire signed [`OutBus]		out_6_3_r;
wire signed [`OutBus]		out_6_3_i;
wire signed [`OutBus]		out_6_4_r;
wire signed [`OutBus]		out_6_4_i;
wire signed [`OutBus]		out_6_5_r;
wire signed [`OutBus]		out_6_5_i;
wire signed [`OutBus]		out_6_6_r;
wire signed [`OutBus]		out_6_6_i;
wire signed [`OutBus]		out_6_7_r;
wire signed [`OutBus]		out_6_7_i;
wire signed [`OutBus]		out_6_8_r;
wire signed [`OutBus]		out_6_8_i;
wire signed [`OutBus]		out_6_9_r;
wire signed [`OutBus]		out_6_9_i;
wire signed [`OutBus]		out_6_10_r;
wire signed [`OutBus]		out_6_10_i;
wire signed [`OutBus]		out_6_11_r;
wire signed [`OutBus]		out_6_11_i;
wire signed [`OutBus]		out_6_12_r;
wire signed [`OutBus]		out_6_12_i;
wire signed [`OutBus]		out_6_13_r;
wire signed [`OutBus]		out_6_13_i;
wire signed [`OutBus]		out_6_14_r;
wire signed [`OutBus]		out_6_14_i;
wire signed [`OutBus]		out_6_15_r;
wire signed [`OutBus]		out_6_15_i;
wire signed [`OutBus]		out_6_16_r;
wire signed [`OutBus]		out_6_16_i;
wire signed [`OutBus]		out_7_1_r;
wire signed [`OutBus]		out_7_1_i;
wire signed [`OutBus]		out_7_2_r;
wire signed [`OutBus]		out_7_2_i;
wire signed [`OutBus]		out_7_3_r;
wire signed [`OutBus]		out_7_3_i;
wire signed [`OutBus]		out_7_4_r;
wire signed [`OutBus]		out_7_4_i;
wire signed [`OutBus]		out_7_5_r;
wire signed [`OutBus]		out_7_5_i;
wire signed [`OutBus]		out_7_6_r;
wire signed [`OutBus]		out_7_6_i;
wire signed [`OutBus]		out_7_7_r;
wire signed [`OutBus]		out_7_7_i;
wire signed [`OutBus]		out_7_8_r;
wire signed [`OutBus]		out_7_8_i;
wire signed [`OutBus]		out_7_9_r;
wire signed [`OutBus]		out_7_9_i;
wire signed [`OutBus]		out_7_10_r;
wire signed [`OutBus]		out_7_10_i;
wire signed [`OutBus]		out_7_11_r;
wire signed [`OutBus]		out_7_11_i;
wire signed [`OutBus]		out_7_12_r;
wire signed [`OutBus]		out_7_12_i;
wire signed [`OutBus]		out_7_13_r;
wire signed [`OutBus]		out_7_13_i;
wire signed [`OutBus]		out_7_14_r;
wire signed [`OutBus]		out_7_14_i;
wire signed [`OutBus]		out_7_15_r;
wire signed [`OutBus]		out_7_15_i;
wire signed [`OutBus]		out_7_16_r;
wire signed [`OutBus]		out_7_16_i;
wire signed [`OutBus]		out_8_1_r;
wire signed [`OutBus]		out_8_1_i;
wire signed [`OutBus]		out_8_2_r;
wire signed [`OutBus]		out_8_2_i;
wire signed [`OutBus]		out_8_3_r;
wire signed [`OutBus]		out_8_3_i;
wire signed [`OutBus]		out_8_4_r;
wire signed [`OutBus]		out_8_4_i;
wire signed [`OutBus]		out_8_5_r;
wire signed [`OutBus]		out_8_5_i;
wire signed [`OutBus]		out_8_6_r;
wire signed [`OutBus]		out_8_6_i;
wire signed [`OutBus]		out_8_7_r;
wire signed [`OutBus]		out_8_7_i;
wire signed [`OutBus]		out_8_8_r;
wire signed [`OutBus]		out_8_8_i;
wire signed [`OutBus]		out_8_9_r;
wire signed [`OutBus]		out_8_9_i;
wire signed [`OutBus]		out_8_10_r;
wire signed [`OutBus]		out_8_10_i;
wire signed [`OutBus]		out_8_11_r;
wire signed [`OutBus]		out_8_11_i;
wire signed [`OutBus]		out_8_12_r;
wire signed [`OutBus]		out_8_12_i;
wire signed [`OutBus]		out_8_13_r;
wire signed [`OutBus]		out_8_13_i;
wire signed [`OutBus]		out_8_14_r;
wire signed [`OutBus]		out_8_14_i;
wire signed [`OutBus]		out_8_15_r;
wire signed [`OutBus]		out_8_15_i;
wire signed [`OutBus]		out_8_16_r;
wire signed [`OutBus]		out_8_16_i;
wire signed [`OutBus]		out_9_1_r;
wire signed [`OutBus]		out_9_1_i;
wire signed [`OutBus]		out_9_2_r;
wire signed [`OutBus]		out_9_2_i;
wire signed [`OutBus]		out_9_3_r;
wire signed [`OutBus]		out_9_3_i;
wire signed [`OutBus]		out_9_4_r;
wire signed [`OutBus]		out_9_4_i;
wire signed [`OutBus]		out_9_5_r;
wire signed [`OutBus]		out_9_5_i;
wire signed [`OutBus]		out_9_6_r;
wire signed [`OutBus]		out_9_6_i;
wire signed [`OutBus]		out_9_7_r;
wire signed [`OutBus]		out_9_7_i;
wire signed [`OutBus]		out_9_8_r;
wire signed [`OutBus]		out_9_8_i;
wire signed [`OutBus]		out_9_9_r;
wire signed [`OutBus]		out_9_9_i;
wire signed [`OutBus]		out_9_10_r;
wire signed [`OutBus]		out_9_10_i;
wire signed [`OutBus]		out_9_11_r;
wire signed [`OutBus]		out_9_11_i;
wire signed [`OutBus]		out_9_12_r;
wire signed [`OutBus]		out_9_12_i;
wire signed [`OutBus]		out_9_13_r;
wire signed [`OutBus]		out_9_13_i;
wire signed [`OutBus]		out_9_14_r;
wire signed [`OutBus]		out_9_14_i;
wire signed [`OutBus]		out_9_15_r;
wire signed [`OutBus]		out_9_15_i;
wire signed [`OutBus]		out_9_16_r;
wire signed [`OutBus]		out_9_16_i;
wire signed [`OutBus]		out_10_1_r;
wire signed [`OutBus]		out_10_1_i;
wire signed [`OutBus]		out_10_2_r;
wire signed [`OutBus]		out_10_2_i;
wire signed [`OutBus]		out_10_3_r;
wire signed [`OutBus]		out_10_3_i;
wire signed [`OutBus]		out_10_4_r;
wire signed [`OutBus]		out_10_4_i;
wire signed [`OutBus]		out_10_5_r;
wire signed [`OutBus]		out_10_5_i;
wire signed [`OutBus]		out_10_6_r;
wire signed [`OutBus]		out_10_6_i;
wire signed [`OutBus]		out_10_7_r;
wire signed [`OutBus]		out_10_7_i;
wire signed [`OutBus]		out_10_8_r;
wire signed [`OutBus]		out_10_8_i;
wire signed [`OutBus]		out_10_9_r;
wire signed [`OutBus]		out_10_9_i;
wire signed [`OutBus]		out_10_10_r;
wire signed [`OutBus]		out_10_10_i;
wire signed [`OutBus]		out_10_11_r;
wire signed [`OutBus]		out_10_11_i;
wire signed [`OutBus]		out_10_12_r;
wire signed [`OutBus]		out_10_12_i;
wire signed [`OutBus]		out_10_13_r;
wire signed [`OutBus]		out_10_13_i;
wire signed [`OutBus]		out_10_14_r;
wire signed [`OutBus]		out_10_14_i;
wire signed [`OutBus]		out_10_15_r;
wire signed [`OutBus]		out_10_15_i;
wire signed [`OutBus]		out_10_16_r;
wire signed [`OutBus]		out_10_16_i;
wire signed [`OutBus]		out_11_1_r;
wire signed [`OutBus]		out_11_1_i;
wire signed [`OutBus]		out_11_2_r;
wire signed [`OutBus]		out_11_2_i;
wire signed [`OutBus]		out_11_3_r;
wire signed [`OutBus]		out_11_3_i;
wire signed [`OutBus]		out_11_4_r;
wire signed [`OutBus]		out_11_4_i;
wire signed [`OutBus]		out_11_5_r;
wire signed [`OutBus]		out_11_5_i;
wire signed [`OutBus]		out_11_6_r;
wire signed [`OutBus]		out_11_6_i;
wire signed [`OutBus]		out_11_7_r;
wire signed [`OutBus]		out_11_7_i;
wire signed [`OutBus]		out_11_8_r;
wire signed [`OutBus]		out_11_8_i;
wire signed [`OutBus]		out_11_9_r;
wire signed [`OutBus]		out_11_9_i;
wire signed [`OutBus]		out_11_10_r;
wire signed [`OutBus]		out_11_10_i;
wire signed [`OutBus]		out_11_11_r;
wire signed [`OutBus]		out_11_11_i;
wire signed [`OutBus]		out_11_12_r;
wire signed [`OutBus]		out_11_12_i;
wire signed [`OutBus]		out_11_13_r;
wire signed [`OutBus]		out_11_13_i;
wire signed [`OutBus]		out_11_14_r;
wire signed [`OutBus]		out_11_14_i;
wire signed [`OutBus]		out_11_15_r;
wire signed [`OutBus]		out_11_15_i;
wire signed [`OutBus]		out_11_16_r;
wire signed [`OutBus]		out_11_16_i;
wire signed [`OutBus]		out_12_1_r;
wire signed [`OutBus]		out_12_1_i;
wire signed [`OutBus]		out_12_2_r;
wire signed [`OutBus]		out_12_2_i;
wire signed [`OutBus]		out_12_3_r;
wire signed [`OutBus]		out_12_3_i;
wire signed [`OutBus]		out_12_4_r;
wire signed [`OutBus]		out_12_4_i;
wire signed [`OutBus]		out_12_5_r;
wire signed [`OutBus]		out_12_5_i;
wire signed [`OutBus]		out_12_6_r;
wire signed [`OutBus]		out_12_6_i;
wire signed [`OutBus]		out_12_7_r;
wire signed [`OutBus]		out_12_7_i;
wire signed [`OutBus]		out_12_8_r;
wire signed [`OutBus]		out_12_8_i;
wire signed [`OutBus]		out_12_9_r;
wire signed [`OutBus]		out_12_9_i;
wire signed [`OutBus]		out_12_10_r;
wire signed [`OutBus]		out_12_10_i;
wire signed [`OutBus]		out_12_11_r;
wire signed [`OutBus]		out_12_11_i;
wire signed [`OutBus]		out_12_12_r;
wire signed [`OutBus]		out_12_12_i;
wire signed [`OutBus]		out_12_13_r;
wire signed [`OutBus]		out_12_13_i;
wire signed [`OutBus]		out_12_14_r;
wire signed [`OutBus]		out_12_14_i;
wire signed [`OutBus]		out_12_15_r;
wire signed [`OutBus]		out_12_15_i;
wire signed [`OutBus]		out_12_16_r;
wire signed [`OutBus]		out_12_16_i;
wire signed [`OutBus]		out_13_1_r;
wire signed [`OutBus]		out_13_1_i;
wire signed [`OutBus]		out_13_2_r;
wire signed [`OutBus]		out_13_2_i;
wire signed [`OutBus]		out_13_3_r;
wire signed [`OutBus]		out_13_3_i;
wire signed [`OutBus]		out_13_4_r;
wire signed [`OutBus]		out_13_4_i;
wire signed [`OutBus]		out_13_5_r;
wire signed [`OutBus]		out_13_5_i;
wire signed [`OutBus]		out_13_6_r;
wire signed [`OutBus]		out_13_6_i;
wire signed [`OutBus]		out_13_7_r;
wire signed [`OutBus]		out_13_7_i;
wire signed [`OutBus]		out_13_8_r;
wire signed [`OutBus]		out_13_8_i;
wire signed [`OutBus]		out_13_9_r;
wire signed [`OutBus]		out_13_9_i;
wire signed [`OutBus]		out_13_10_r;
wire signed [`OutBus]		out_13_10_i;
wire signed [`OutBus]		out_13_11_r;
wire signed [`OutBus]		out_13_11_i;
wire signed [`OutBus]		out_13_12_r;
wire signed [`OutBus]		out_13_12_i;
wire signed [`OutBus]		out_13_13_r;
wire signed [`OutBus]		out_13_13_i;
wire signed [`OutBus]		out_13_14_r;
wire signed [`OutBus]		out_13_14_i;
wire signed [`OutBus]		out_13_15_r;
wire signed [`OutBus]		out_13_15_i;
wire signed [`OutBus]		out_13_16_r;
wire signed [`OutBus]		out_13_16_i;
wire signed [`OutBus]		out_14_1_r;
wire signed [`OutBus]		out_14_1_i;
wire signed [`OutBus]		out_14_2_r;
wire signed [`OutBus]		out_14_2_i;
wire signed [`OutBus]		out_14_3_r;
wire signed [`OutBus]		out_14_3_i;
wire signed [`OutBus]		out_14_4_r;
wire signed [`OutBus]		out_14_4_i;
wire signed [`OutBus]		out_14_5_r;
wire signed [`OutBus]		out_14_5_i;
wire signed [`OutBus]		out_14_6_r;
wire signed [`OutBus]		out_14_6_i;
wire signed [`OutBus]		out_14_7_r;
wire signed [`OutBus]		out_14_7_i;
wire signed [`OutBus]		out_14_8_r;
wire signed [`OutBus]		out_14_8_i;
wire signed [`OutBus]		out_14_9_r;
wire signed [`OutBus]		out_14_9_i;
wire signed [`OutBus]		out_14_10_r;
wire signed [`OutBus]		out_14_10_i;
wire signed [`OutBus]		out_14_11_r;
wire signed [`OutBus]		out_14_11_i;
wire signed [`OutBus]		out_14_12_r;
wire signed [`OutBus]		out_14_12_i;
wire signed [`OutBus]		out_14_13_r;
wire signed [`OutBus]		out_14_13_i;
wire signed [`OutBus]		out_14_14_r;
wire signed [`OutBus]		out_14_14_i;
wire signed [`OutBus]		out_14_15_r;
wire signed [`OutBus]		out_14_15_i;
wire signed [`OutBus]		out_14_16_r;
wire signed [`OutBus]		out_14_16_i;
wire signed [`OutBus]		out_15_1_r;
wire signed [`OutBus]		out_15_1_i;
wire signed [`OutBus]		out_15_2_r;
wire signed [`OutBus]		out_15_2_i;
wire signed [`OutBus]		out_15_3_r;
wire signed [`OutBus]		out_15_3_i;
wire signed [`OutBus]		out_15_4_r;
wire signed [`OutBus]		out_15_4_i;
wire signed [`OutBus]		out_15_5_r;
wire signed [`OutBus]		out_15_5_i;
wire signed [`OutBus]		out_15_6_r;
wire signed [`OutBus]		out_15_6_i;
wire signed [`OutBus]		out_15_7_r;
wire signed [`OutBus]		out_15_7_i;
wire signed [`OutBus]		out_15_8_r;
wire signed [`OutBus]		out_15_8_i;
wire signed [`OutBus]		out_15_9_r;
wire signed [`OutBus]		out_15_9_i;
wire signed [`OutBus]		out_15_10_r;
wire signed [`OutBus]		out_15_10_i;
wire signed [`OutBus]		out_15_11_r;
wire signed [`OutBus]		out_15_11_i;
wire signed [`OutBus]		out_15_12_r;
wire signed [`OutBus]		out_15_12_i;
wire signed [`OutBus]		out_15_13_r;
wire signed [`OutBus]		out_15_13_i;
wire signed [`OutBus]		out_15_14_r;
wire signed [`OutBus]		out_15_14_i;
wire signed [`OutBus]		out_15_15_r;
wire signed [`OutBus]		out_15_15_i;
wire signed [`OutBus]		out_15_16_r;
wire signed [`OutBus]		out_15_16_i;
wire signed [`OutBus]		out_16_1_r;
wire signed [`OutBus]		out_16_1_i;
wire signed [`OutBus]		out_16_2_r;
wire signed [`OutBus]		out_16_2_i;
wire signed [`OutBus]		out_16_3_r;
wire signed [`OutBus]		out_16_3_i;
wire signed [`OutBus]		out_16_4_r;
wire signed [`OutBus]		out_16_4_i;
wire signed [`OutBus]		out_16_5_r;
wire signed [`OutBus]		out_16_5_i;
wire signed [`OutBus]		out_16_6_r;
wire signed [`OutBus]		out_16_6_i;
wire signed [`OutBus]		out_16_7_r;
wire signed [`OutBus]		out_16_7_i;
wire signed [`OutBus]		out_16_8_r;
wire signed [`OutBus]		out_16_8_i;
wire signed [`OutBus]		out_16_9_r;
wire signed [`OutBus]		out_16_9_i;
wire signed [`OutBus]		out_16_10_r;
wire signed [`OutBus]		out_16_10_i;
wire signed [`OutBus]		out_16_11_r;
wire signed [`OutBus]		out_16_11_i;
wire signed [`OutBus]		out_16_12_r;
wire signed [`OutBus]		out_16_12_i;
wire signed [`OutBus]		out_16_13_r;
wire signed [`OutBus]		out_16_13_i;
wire signed [`OutBus]		out_16_14_r;
wire signed [`OutBus]		out_16_14_i;
wire signed [`OutBus]		out_16_15_r;
wire signed [`OutBus]		out_16_15_i;
wire signed [`OutBus]		out_16_16_r;
wire signed [`OutBus]		out_16_16_i;

/************************temp MUX butterfly***********************/
wire signed [`CalcTempBus]          temp_m1_1_1_r;
wire signed [`CalcTempBus]          temp_m1_1_1_i;
wire signed [`CalcTempBus]          temp_m1_1_2_r;
wire signed [`CalcTempBus]          temp_m1_1_2_i;
wire signed [`CalcTempBus]          temp_m1_1_3_r;
wire signed [`CalcTempBus]          temp_m1_1_3_i;
wire signed [`CalcTempBus]          temp_m1_1_4_r;
wire signed [`CalcTempBus]          temp_m1_1_4_i;
wire signed [`CalcTempBus]          temp_m1_1_5_r;
wire signed [`CalcTempBus]          temp_m1_1_5_i;
wire signed [`CalcTempBus]          temp_m1_1_6_r;
wire signed [`CalcTempBus]          temp_m1_1_6_i;
wire signed [`CalcTempBus]          temp_m1_1_7_r;
wire signed [`CalcTempBus]          temp_m1_1_7_i;
wire signed [`CalcTempBus]          temp_m1_1_8_r;
wire signed [`CalcTempBus]          temp_m1_1_8_i;
wire signed [`CalcTempBus]          temp_m1_1_9_r;
wire signed [`CalcTempBus]          temp_m1_1_9_i;
wire signed [`CalcTempBus]          temp_m1_1_10_r;
wire signed [`CalcTempBus]          temp_m1_1_10_i;
wire signed [`CalcTempBus]          temp_m1_1_11_r;
wire signed [`CalcTempBus]          temp_m1_1_11_i;
wire signed [`CalcTempBus]          temp_m1_1_12_r;
wire signed [`CalcTempBus]          temp_m1_1_12_i;
wire signed [`CalcTempBus]          temp_m1_1_13_r;
wire signed [`CalcTempBus]          temp_m1_1_13_i;
wire signed [`CalcTempBus]          temp_m1_1_14_r;
wire signed [`CalcTempBus]          temp_m1_1_14_i;
wire signed [`CalcTempBus]          temp_m1_1_15_r;
wire signed [`CalcTempBus]          temp_m1_1_15_i;
wire signed [`CalcTempBus]          temp_m1_1_16_r;
wire signed [`CalcTempBus]          temp_m1_1_16_i;
wire signed [`CalcTempBus]          temp_m1_2_1_r;
wire signed [`CalcTempBus]          temp_m1_2_1_i;
wire signed [`CalcTempBus]          temp_m1_2_2_r;
wire signed [`CalcTempBus]          temp_m1_2_2_i;
wire signed [`CalcTempBus]          temp_m1_2_3_r;
wire signed [`CalcTempBus]          temp_m1_2_3_i;
wire signed [`CalcTempBus]          temp_m1_2_4_r;
wire signed [`CalcTempBus]          temp_m1_2_4_i;
wire signed [`CalcTempBus]          temp_m1_2_5_r;
wire signed [`CalcTempBus]          temp_m1_2_5_i;
wire signed [`CalcTempBus]          temp_m1_2_6_r;
wire signed [`CalcTempBus]          temp_m1_2_6_i;
wire signed [`CalcTempBus]          temp_m1_2_7_r;
wire signed [`CalcTempBus]          temp_m1_2_7_i;
wire signed [`CalcTempBus]          temp_m1_2_8_r;
wire signed [`CalcTempBus]          temp_m1_2_8_i;
wire signed [`CalcTempBus]          temp_m1_2_9_r;
wire signed [`CalcTempBus]          temp_m1_2_9_i;
wire signed [`CalcTempBus]          temp_m1_2_10_r;
wire signed [`CalcTempBus]          temp_m1_2_10_i;
wire signed [`CalcTempBus]          temp_m1_2_11_r;
wire signed [`CalcTempBus]          temp_m1_2_11_i;
wire signed [`CalcTempBus]          temp_m1_2_12_r;
wire signed [`CalcTempBus]          temp_m1_2_12_i;
wire signed [`CalcTempBus]          temp_m1_2_13_r;
wire signed [`CalcTempBus]          temp_m1_2_13_i;
wire signed [`CalcTempBus]          temp_m1_2_14_r;
wire signed [`CalcTempBus]          temp_m1_2_14_i;
wire signed [`CalcTempBus]          temp_m1_2_15_r;
wire signed [`CalcTempBus]          temp_m1_2_15_i;
wire signed [`CalcTempBus]          temp_m1_2_16_r;
wire signed [`CalcTempBus]          temp_m1_2_16_i;
wire signed [`CalcTempBus]          temp_m1_3_1_r;
wire signed [`CalcTempBus]          temp_m1_3_1_i;
wire signed [`CalcTempBus]          temp_m1_3_2_r;
wire signed [`CalcTempBus]          temp_m1_3_2_i;
wire signed [`CalcTempBus]          temp_m1_3_3_r;
wire signed [`CalcTempBus]          temp_m1_3_3_i;
wire signed [`CalcTempBus]          temp_m1_3_4_r;
wire signed [`CalcTempBus]          temp_m1_3_4_i;
wire signed [`CalcTempBus]          temp_m1_3_5_r;
wire signed [`CalcTempBus]          temp_m1_3_5_i;
wire signed [`CalcTempBus]          temp_m1_3_6_r;
wire signed [`CalcTempBus]          temp_m1_3_6_i;
wire signed [`CalcTempBus]          temp_m1_3_7_r;
wire signed [`CalcTempBus]          temp_m1_3_7_i;
wire signed [`CalcTempBus]          temp_m1_3_8_r;
wire signed [`CalcTempBus]          temp_m1_3_8_i;
wire signed [`CalcTempBus]          temp_m1_3_9_r;
wire signed [`CalcTempBus]          temp_m1_3_9_i;
wire signed [`CalcTempBus]          temp_m1_3_10_r;
wire signed [`CalcTempBus]          temp_m1_3_10_i;
wire signed [`CalcTempBus]          temp_m1_3_11_r;
wire signed [`CalcTempBus]          temp_m1_3_11_i;
wire signed [`CalcTempBus]          temp_m1_3_12_r;
wire signed [`CalcTempBus]          temp_m1_3_12_i;
wire signed [`CalcTempBus]          temp_m1_3_13_r;
wire signed [`CalcTempBus]          temp_m1_3_13_i;
wire signed [`CalcTempBus]          temp_m1_3_14_r;
wire signed [`CalcTempBus]          temp_m1_3_14_i;
wire signed [`CalcTempBus]          temp_m1_3_15_r;
wire signed [`CalcTempBus]          temp_m1_3_15_i;
wire signed [`CalcTempBus]          temp_m1_3_16_r;
wire signed [`CalcTempBus]          temp_m1_3_16_i;
wire signed [`CalcTempBus]          temp_m1_4_1_r;
wire signed [`CalcTempBus]          temp_m1_4_1_i;
wire signed [`CalcTempBus]          temp_m1_4_2_r;
wire signed [`CalcTempBus]          temp_m1_4_2_i;
wire signed [`CalcTempBus]          temp_m1_4_3_r;
wire signed [`CalcTempBus]          temp_m1_4_3_i;
wire signed [`CalcTempBus]          temp_m1_4_4_r;
wire signed [`CalcTempBus]          temp_m1_4_4_i;
wire signed [`CalcTempBus]          temp_m1_4_5_r;
wire signed [`CalcTempBus]          temp_m1_4_5_i;
wire signed [`CalcTempBus]          temp_m1_4_6_r;
wire signed [`CalcTempBus]          temp_m1_4_6_i;
wire signed [`CalcTempBus]          temp_m1_4_7_r;
wire signed [`CalcTempBus]          temp_m1_4_7_i;
wire signed [`CalcTempBus]          temp_m1_4_8_r;
wire signed [`CalcTempBus]          temp_m1_4_8_i;
wire signed [`CalcTempBus]          temp_m1_4_9_r;
wire signed [`CalcTempBus]          temp_m1_4_9_i;
wire signed [`CalcTempBus]          temp_m1_4_10_r;
wire signed [`CalcTempBus]          temp_m1_4_10_i;
wire signed [`CalcTempBus]          temp_m1_4_11_r;
wire signed [`CalcTempBus]          temp_m1_4_11_i;
wire signed [`CalcTempBus]          temp_m1_4_12_r;
wire signed [`CalcTempBus]          temp_m1_4_12_i;
wire signed [`CalcTempBus]          temp_m1_4_13_r;
wire signed [`CalcTempBus]          temp_m1_4_13_i;
wire signed [`CalcTempBus]          temp_m1_4_14_r;
wire signed [`CalcTempBus]          temp_m1_4_14_i;
wire signed [`CalcTempBus]          temp_m1_4_15_r;
wire signed [`CalcTempBus]          temp_m1_4_15_i;
wire signed [`CalcTempBus]          temp_m1_4_16_r;
wire signed [`CalcTempBus]          temp_m1_4_16_i;
wire signed [`CalcTempBus]          temp_m1_5_1_r;
wire signed [`CalcTempBus]          temp_m1_5_1_i;
wire signed [`CalcTempBus]          temp_m1_5_2_r;
wire signed [`CalcTempBus]          temp_m1_5_2_i;
wire signed [`CalcTempBus]          temp_m1_5_3_r;
wire signed [`CalcTempBus]          temp_m1_5_3_i;
wire signed [`CalcTempBus]          temp_m1_5_4_r;
wire signed [`CalcTempBus]          temp_m1_5_4_i;
wire signed [`CalcTempBus]          temp_m1_5_5_r;
wire signed [`CalcTempBus]          temp_m1_5_5_i;
wire signed [`CalcTempBus]          temp_m1_5_6_r;
wire signed [`CalcTempBus]          temp_m1_5_6_i;
wire signed [`CalcTempBus]          temp_m1_5_7_r;
wire signed [`CalcTempBus]          temp_m1_5_7_i;
wire signed [`CalcTempBus]          temp_m1_5_8_r;
wire signed [`CalcTempBus]          temp_m1_5_8_i;
wire signed [`CalcTempBus]          temp_m1_5_9_r;
wire signed [`CalcTempBus]          temp_m1_5_9_i;
wire signed [`CalcTempBus]          temp_m1_5_10_r;
wire signed [`CalcTempBus]          temp_m1_5_10_i;
wire signed [`CalcTempBus]          temp_m1_5_11_r;
wire signed [`CalcTempBus]          temp_m1_5_11_i;
wire signed [`CalcTempBus]          temp_m1_5_12_r;
wire signed [`CalcTempBus]          temp_m1_5_12_i;
wire signed [`CalcTempBus]          temp_m1_5_13_r;
wire signed [`CalcTempBus]          temp_m1_5_13_i;
wire signed [`CalcTempBus]          temp_m1_5_14_r;
wire signed [`CalcTempBus]          temp_m1_5_14_i;
wire signed [`CalcTempBus]          temp_m1_5_15_r;
wire signed [`CalcTempBus]          temp_m1_5_15_i;
wire signed [`CalcTempBus]          temp_m1_5_16_r;
wire signed [`CalcTempBus]          temp_m1_5_16_i;
wire signed [`CalcTempBus]          temp_m1_6_1_r;
wire signed [`CalcTempBus]          temp_m1_6_1_i;
wire signed [`CalcTempBus]          temp_m1_6_2_r;
wire signed [`CalcTempBus]          temp_m1_6_2_i;
wire signed [`CalcTempBus]          temp_m1_6_3_r;
wire signed [`CalcTempBus]          temp_m1_6_3_i;
wire signed [`CalcTempBus]          temp_m1_6_4_r;
wire signed [`CalcTempBus]          temp_m1_6_4_i;
wire signed [`CalcTempBus]          temp_m1_6_5_r;
wire signed [`CalcTempBus]          temp_m1_6_5_i;
wire signed [`CalcTempBus]          temp_m1_6_6_r;
wire signed [`CalcTempBus]          temp_m1_6_6_i;
wire signed [`CalcTempBus]          temp_m1_6_7_r;
wire signed [`CalcTempBus]          temp_m1_6_7_i;
wire signed [`CalcTempBus]          temp_m1_6_8_r;
wire signed [`CalcTempBus]          temp_m1_6_8_i;
wire signed [`CalcTempBus]          temp_m1_6_9_r;
wire signed [`CalcTempBus]          temp_m1_6_9_i;
wire signed [`CalcTempBus]          temp_m1_6_10_r;
wire signed [`CalcTempBus]          temp_m1_6_10_i;
wire signed [`CalcTempBus]          temp_m1_6_11_r;
wire signed [`CalcTempBus]          temp_m1_6_11_i;
wire signed [`CalcTempBus]          temp_m1_6_12_r;
wire signed [`CalcTempBus]          temp_m1_6_12_i;
wire signed [`CalcTempBus]          temp_m1_6_13_r;
wire signed [`CalcTempBus]          temp_m1_6_13_i;
wire signed [`CalcTempBus]          temp_m1_6_14_r;
wire signed [`CalcTempBus]          temp_m1_6_14_i;
wire signed [`CalcTempBus]          temp_m1_6_15_r;
wire signed [`CalcTempBus]          temp_m1_6_15_i;
wire signed [`CalcTempBus]          temp_m1_6_16_r;
wire signed [`CalcTempBus]          temp_m1_6_16_i;
wire signed [`CalcTempBus]          temp_m1_7_1_r;
wire signed [`CalcTempBus]          temp_m1_7_1_i;
wire signed [`CalcTempBus]          temp_m1_7_2_r;
wire signed [`CalcTempBus]          temp_m1_7_2_i;
wire signed [`CalcTempBus]          temp_m1_7_3_r;
wire signed [`CalcTempBus]          temp_m1_7_3_i;
wire signed [`CalcTempBus]          temp_m1_7_4_r;
wire signed [`CalcTempBus]          temp_m1_7_4_i;
wire signed [`CalcTempBus]          temp_m1_7_5_r;
wire signed [`CalcTempBus]          temp_m1_7_5_i;
wire signed [`CalcTempBus]          temp_m1_7_6_r;
wire signed [`CalcTempBus]          temp_m1_7_6_i;
wire signed [`CalcTempBus]          temp_m1_7_7_r;
wire signed [`CalcTempBus]          temp_m1_7_7_i;
wire signed [`CalcTempBus]          temp_m1_7_8_r;
wire signed [`CalcTempBus]          temp_m1_7_8_i;
wire signed [`CalcTempBus]          temp_m1_7_9_r;
wire signed [`CalcTempBus]          temp_m1_7_9_i;
wire signed [`CalcTempBus]          temp_m1_7_10_r;
wire signed [`CalcTempBus]          temp_m1_7_10_i;
wire signed [`CalcTempBus]          temp_m1_7_11_r;
wire signed [`CalcTempBus]          temp_m1_7_11_i;
wire signed [`CalcTempBus]          temp_m1_7_12_r;
wire signed [`CalcTempBus]          temp_m1_7_12_i;
wire signed [`CalcTempBus]          temp_m1_7_13_r;
wire signed [`CalcTempBus]          temp_m1_7_13_i;
wire signed [`CalcTempBus]          temp_m1_7_14_r;
wire signed [`CalcTempBus]          temp_m1_7_14_i;
wire signed [`CalcTempBus]          temp_m1_7_15_r;
wire signed [`CalcTempBus]          temp_m1_7_15_i;
wire signed [`CalcTempBus]          temp_m1_7_16_r;
wire signed [`CalcTempBus]          temp_m1_7_16_i;
wire signed [`CalcTempBus]          temp_m1_8_1_r;
wire signed [`CalcTempBus]          temp_m1_8_1_i;
wire signed [`CalcTempBus]          temp_m1_8_2_r;
wire signed [`CalcTempBus]          temp_m1_8_2_i;
wire signed [`CalcTempBus]          temp_m1_8_3_r;
wire signed [`CalcTempBus]          temp_m1_8_3_i;
wire signed [`CalcTempBus]          temp_m1_8_4_r;
wire signed [`CalcTempBus]          temp_m1_8_4_i;
wire signed [`CalcTempBus]          temp_m1_8_5_r;
wire signed [`CalcTempBus]          temp_m1_8_5_i;
wire signed [`CalcTempBus]          temp_m1_8_6_r;
wire signed [`CalcTempBus]          temp_m1_8_6_i;
wire signed [`CalcTempBus]          temp_m1_8_7_r;
wire signed [`CalcTempBus]          temp_m1_8_7_i;
wire signed [`CalcTempBus]          temp_m1_8_8_r;
wire signed [`CalcTempBus]          temp_m1_8_8_i;
wire signed [`CalcTempBus]          temp_m1_8_9_r;
wire signed [`CalcTempBus]          temp_m1_8_9_i;
wire signed [`CalcTempBus]          temp_m1_8_10_r;
wire signed [`CalcTempBus]          temp_m1_8_10_i;
wire signed [`CalcTempBus]          temp_m1_8_11_r;
wire signed [`CalcTempBus]          temp_m1_8_11_i;
wire signed [`CalcTempBus]          temp_m1_8_12_r;
wire signed [`CalcTempBus]          temp_m1_8_12_i;
wire signed [`CalcTempBus]          temp_m1_8_13_r;
wire signed [`CalcTempBus]          temp_m1_8_13_i;
wire signed [`CalcTempBus]          temp_m1_8_14_r;
wire signed [`CalcTempBus]          temp_m1_8_14_i;
wire signed [`CalcTempBus]          temp_m1_8_15_r;
wire signed [`CalcTempBus]          temp_m1_8_15_i;
wire signed [`CalcTempBus]          temp_m1_8_16_r;
wire signed [`CalcTempBus]          temp_m1_8_16_i;
wire signed [`CalcTempBus]          temp_m1_9_1_r;
wire signed [`CalcTempBus]          temp_m1_9_1_i;
wire signed [`CalcTempBus]          temp_m1_9_2_r;
wire signed [`CalcTempBus]          temp_m1_9_2_i;
wire signed [`CalcTempBus]          temp_m1_9_3_r;
wire signed [`CalcTempBus]          temp_m1_9_3_i;
wire signed [`CalcTempBus]          temp_m1_9_4_r;
wire signed [`CalcTempBus]          temp_m1_9_4_i;
wire signed [`CalcTempBus]          temp_m1_9_5_r;
wire signed [`CalcTempBus]          temp_m1_9_5_i;
wire signed [`CalcTempBus]          temp_m1_9_6_r;
wire signed [`CalcTempBus]          temp_m1_9_6_i;
wire signed [`CalcTempBus]          temp_m1_9_7_r;
wire signed [`CalcTempBus]          temp_m1_9_7_i;
wire signed [`CalcTempBus]          temp_m1_9_8_r;
wire signed [`CalcTempBus]          temp_m1_9_8_i;
wire signed [`CalcTempBus]          temp_m1_9_9_r;
wire signed [`CalcTempBus]          temp_m1_9_9_i;
wire signed [`CalcTempBus]          temp_m1_9_10_r;
wire signed [`CalcTempBus]          temp_m1_9_10_i;
wire signed [`CalcTempBus]          temp_m1_9_11_r;
wire signed [`CalcTempBus]          temp_m1_9_11_i;
wire signed [`CalcTempBus]          temp_m1_9_12_r;
wire signed [`CalcTempBus]          temp_m1_9_12_i;
wire signed [`CalcTempBus]          temp_m1_9_13_r;
wire signed [`CalcTempBus]          temp_m1_9_13_i;
wire signed [`CalcTempBus]          temp_m1_9_14_r;
wire signed [`CalcTempBus]          temp_m1_9_14_i;
wire signed [`CalcTempBus]          temp_m1_9_15_r;
wire signed [`CalcTempBus]          temp_m1_9_15_i;
wire signed [`CalcTempBus]          temp_m1_9_16_r;
wire signed [`CalcTempBus]          temp_m1_9_16_i;
wire signed [`CalcTempBus]          temp_m1_10_1_r;
wire signed [`CalcTempBus]          temp_m1_10_1_i;
wire signed [`CalcTempBus]          temp_m1_10_2_r;
wire signed [`CalcTempBus]          temp_m1_10_2_i;
wire signed [`CalcTempBus]          temp_m1_10_3_r;
wire signed [`CalcTempBus]          temp_m1_10_3_i;
wire signed [`CalcTempBus]          temp_m1_10_4_r;
wire signed [`CalcTempBus]          temp_m1_10_4_i;
wire signed [`CalcTempBus]          temp_m1_10_5_r;
wire signed [`CalcTempBus]          temp_m1_10_5_i;
wire signed [`CalcTempBus]          temp_m1_10_6_r;
wire signed [`CalcTempBus]          temp_m1_10_6_i;
wire signed [`CalcTempBus]          temp_m1_10_7_r;
wire signed [`CalcTempBus]          temp_m1_10_7_i;
wire signed [`CalcTempBus]          temp_m1_10_8_r;
wire signed [`CalcTempBus]          temp_m1_10_8_i;
wire signed [`CalcTempBus]          temp_m1_10_9_r;
wire signed [`CalcTempBus]          temp_m1_10_9_i;
wire signed [`CalcTempBus]          temp_m1_10_10_r;
wire signed [`CalcTempBus]          temp_m1_10_10_i;
wire signed [`CalcTempBus]          temp_m1_10_11_r;
wire signed [`CalcTempBus]          temp_m1_10_11_i;
wire signed [`CalcTempBus]          temp_m1_10_12_r;
wire signed [`CalcTempBus]          temp_m1_10_12_i;
wire signed [`CalcTempBus]          temp_m1_10_13_r;
wire signed [`CalcTempBus]          temp_m1_10_13_i;
wire signed [`CalcTempBus]          temp_m1_10_14_r;
wire signed [`CalcTempBus]          temp_m1_10_14_i;
wire signed [`CalcTempBus]          temp_m1_10_15_r;
wire signed [`CalcTempBus]          temp_m1_10_15_i;
wire signed [`CalcTempBus]          temp_m1_10_16_r;
wire signed [`CalcTempBus]          temp_m1_10_16_i;
wire signed [`CalcTempBus]          temp_m1_11_1_r;
wire signed [`CalcTempBus]          temp_m1_11_1_i;
wire signed [`CalcTempBus]          temp_m1_11_2_r;
wire signed [`CalcTempBus]          temp_m1_11_2_i;
wire signed [`CalcTempBus]          temp_m1_11_3_r;
wire signed [`CalcTempBus]          temp_m1_11_3_i;
wire signed [`CalcTempBus]          temp_m1_11_4_r;
wire signed [`CalcTempBus]          temp_m1_11_4_i;
wire signed [`CalcTempBus]          temp_m1_11_5_r;
wire signed [`CalcTempBus]          temp_m1_11_5_i;
wire signed [`CalcTempBus]          temp_m1_11_6_r;
wire signed [`CalcTempBus]          temp_m1_11_6_i;
wire signed [`CalcTempBus]          temp_m1_11_7_r;
wire signed [`CalcTempBus]          temp_m1_11_7_i;
wire signed [`CalcTempBus]          temp_m1_11_8_r;
wire signed [`CalcTempBus]          temp_m1_11_8_i;
wire signed [`CalcTempBus]          temp_m1_11_9_r;
wire signed [`CalcTempBus]          temp_m1_11_9_i;
wire signed [`CalcTempBus]          temp_m1_11_10_r;
wire signed [`CalcTempBus]          temp_m1_11_10_i;
wire signed [`CalcTempBus]          temp_m1_11_11_r;
wire signed [`CalcTempBus]          temp_m1_11_11_i;
wire signed [`CalcTempBus]          temp_m1_11_12_r;
wire signed [`CalcTempBus]          temp_m1_11_12_i;
wire signed [`CalcTempBus]          temp_m1_11_13_r;
wire signed [`CalcTempBus]          temp_m1_11_13_i;
wire signed [`CalcTempBus]          temp_m1_11_14_r;
wire signed [`CalcTempBus]          temp_m1_11_14_i;
wire signed [`CalcTempBus]          temp_m1_11_15_r;
wire signed [`CalcTempBus]          temp_m1_11_15_i;
wire signed [`CalcTempBus]          temp_m1_11_16_r;
wire signed [`CalcTempBus]          temp_m1_11_16_i;
wire signed [`CalcTempBus]          temp_m1_12_1_r;
wire signed [`CalcTempBus]          temp_m1_12_1_i;
wire signed [`CalcTempBus]          temp_m1_12_2_r;
wire signed [`CalcTempBus]          temp_m1_12_2_i;
wire signed [`CalcTempBus]          temp_m1_12_3_r;
wire signed [`CalcTempBus]          temp_m1_12_3_i;
wire signed [`CalcTempBus]          temp_m1_12_4_r;
wire signed [`CalcTempBus]          temp_m1_12_4_i;
wire signed [`CalcTempBus]          temp_m1_12_5_r;
wire signed [`CalcTempBus]          temp_m1_12_5_i;
wire signed [`CalcTempBus]          temp_m1_12_6_r;
wire signed [`CalcTempBus]          temp_m1_12_6_i;
wire signed [`CalcTempBus]          temp_m1_12_7_r;
wire signed [`CalcTempBus]          temp_m1_12_7_i;
wire signed [`CalcTempBus]          temp_m1_12_8_r;
wire signed [`CalcTempBus]          temp_m1_12_8_i;
wire signed [`CalcTempBus]          temp_m1_12_9_r;
wire signed [`CalcTempBus]          temp_m1_12_9_i;
wire signed [`CalcTempBus]          temp_m1_12_10_r;
wire signed [`CalcTempBus]          temp_m1_12_10_i;
wire signed [`CalcTempBus]          temp_m1_12_11_r;
wire signed [`CalcTempBus]          temp_m1_12_11_i;
wire signed [`CalcTempBus]          temp_m1_12_12_r;
wire signed [`CalcTempBus]          temp_m1_12_12_i;
wire signed [`CalcTempBus]          temp_m1_12_13_r;
wire signed [`CalcTempBus]          temp_m1_12_13_i;
wire signed [`CalcTempBus]          temp_m1_12_14_r;
wire signed [`CalcTempBus]          temp_m1_12_14_i;
wire signed [`CalcTempBus]          temp_m1_12_15_r;
wire signed [`CalcTempBus]          temp_m1_12_15_i;
wire signed [`CalcTempBus]          temp_m1_12_16_r;
wire signed [`CalcTempBus]          temp_m1_12_16_i;
wire signed [`CalcTempBus]          temp_m1_13_1_r;
wire signed [`CalcTempBus]          temp_m1_13_1_i;
wire signed [`CalcTempBus]          temp_m1_13_2_r;
wire signed [`CalcTempBus]          temp_m1_13_2_i;
wire signed [`CalcTempBus]          temp_m1_13_3_r;
wire signed [`CalcTempBus]          temp_m1_13_3_i;
wire signed [`CalcTempBus]          temp_m1_13_4_r;
wire signed [`CalcTempBus]          temp_m1_13_4_i;
wire signed [`CalcTempBus]          temp_m1_13_5_r;
wire signed [`CalcTempBus]          temp_m1_13_5_i;
wire signed [`CalcTempBus]          temp_m1_13_6_r;
wire signed [`CalcTempBus]          temp_m1_13_6_i;
wire signed [`CalcTempBus]          temp_m1_13_7_r;
wire signed [`CalcTempBus]          temp_m1_13_7_i;
wire signed [`CalcTempBus]          temp_m1_13_8_r;
wire signed [`CalcTempBus]          temp_m1_13_8_i;
wire signed [`CalcTempBus]          temp_m1_13_9_r;
wire signed [`CalcTempBus]          temp_m1_13_9_i;
wire signed [`CalcTempBus]          temp_m1_13_10_r;
wire signed [`CalcTempBus]          temp_m1_13_10_i;
wire signed [`CalcTempBus]          temp_m1_13_11_r;
wire signed [`CalcTempBus]          temp_m1_13_11_i;
wire signed [`CalcTempBus]          temp_m1_13_12_r;
wire signed [`CalcTempBus]          temp_m1_13_12_i;
wire signed [`CalcTempBus]          temp_m1_13_13_r;
wire signed [`CalcTempBus]          temp_m1_13_13_i;
wire signed [`CalcTempBus]          temp_m1_13_14_r;
wire signed [`CalcTempBus]          temp_m1_13_14_i;
wire signed [`CalcTempBus]          temp_m1_13_15_r;
wire signed [`CalcTempBus]          temp_m1_13_15_i;
wire signed [`CalcTempBus]          temp_m1_13_16_r;
wire signed [`CalcTempBus]          temp_m1_13_16_i;
wire signed [`CalcTempBus]          temp_m1_14_1_r;
wire signed [`CalcTempBus]          temp_m1_14_1_i;
wire signed [`CalcTempBus]          temp_m1_14_2_r;
wire signed [`CalcTempBus]          temp_m1_14_2_i;
wire signed [`CalcTempBus]          temp_m1_14_3_r;
wire signed [`CalcTempBus]          temp_m1_14_3_i;
wire signed [`CalcTempBus]          temp_m1_14_4_r;
wire signed [`CalcTempBus]          temp_m1_14_4_i;
wire signed [`CalcTempBus]          temp_m1_14_5_r;
wire signed [`CalcTempBus]          temp_m1_14_5_i;
wire signed [`CalcTempBus]          temp_m1_14_6_r;
wire signed [`CalcTempBus]          temp_m1_14_6_i;
wire signed [`CalcTempBus]          temp_m1_14_7_r;
wire signed [`CalcTempBus]          temp_m1_14_7_i;
wire signed [`CalcTempBus]          temp_m1_14_8_r;
wire signed [`CalcTempBus]          temp_m1_14_8_i;
wire signed [`CalcTempBus]          temp_m1_14_9_r;
wire signed [`CalcTempBus]          temp_m1_14_9_i;
wire signed [`CalcTempBus]          temp_m1_14_10_r;
wire signed [`CalcTempBus]          temp_m1_14_10_i;
wire signed [`CalcTempBus]          temp_m1_14_11_r;
wire signed [`CalcTempBus]          temp_m1_14_11_i;
wire signed [`CalcTempBus]          temp_m1_14_12_r;
wire signed [`CalcTempBus]          temp_m1_14_12_i;
wire signed [`CalcTempBus]          temp_m1_14_13_r;
wire signed [`CalcTempBus]          temp_m1_14_13_i;
wire signed [`CalcTempBus]          temp_m1_14_14_r;
wire signed [`CalcTempBus]          temp_m1_14_14_i;
wire signed [`CalcTempBus]          temp_m1_14_15_r;
wire signed [`CalcTempBus]          temp_m1_14_15_i;
wire signed [`CalcTempBus]          temp_m1_14_16_r;
wire signed [`CalcTempBus]          temp_m1_14_16_i;
wire signed [`CalcTempBus]          temp_m1_15_1_r;
wire signed [`CalcTempBus]          temp_m1_15_1_i;
wire signed [`CalcTempBus]          temp_m1_15_2_r;
wire signed [`CalcTempBus]          temp_m1_15_2_i;
wire signed [`CalcTempBus]          temp_m1_15_3_r;
wire signed [`CalcTempBus]          temp_m1_15_3_i;
wire signed [`CalcTempBus]          temp_m1_15_4_r;
wire signed [`CalcTempBus]          temp_m1_15_4_i;
wire signed [`CalcTempBus]          temp_m1_15_5_r;
wire signed [`CalcTempBus]          temp_m1_15_5_i;
wire signed [`CalcTempBus]          temp_m1_15_6_r;
wire signed [`CalcTempBus]          temp_m1_15_6_i;
wire signed [`CalcTempBus]          temp_m1_15_7_r;
wire signed [`CalcTempBus]          temp_m1_15_7_i;
wire signed [`CalcTempBus]          temp_m1_15_8_r;
wire signed [`CalcTempBus]          temp_m1_15_8_i;
wire signed [`CalcTempBus]          temp_m1_15_9_r;
wire signed [`CalcTempBus]          temp_m1_15_9_i;
wire signed [`CalcTempBus]          temp_m1_15_10_r;
wire signed [`CalcTempBus]          temp_m1_15_10_i;
wire signed [`CalcTempBus]          temp_m1_15_11_r;
wire signed [`CalcTempBus]          temp_m1_15_11_i;
wire signed [`CalcTempBus]          temp_m1_15_12_r;
wire signed [`CalcTempBus]          temp_m1_15_12_i;
wire signed [`CalcTempBus]          temp_m1_15_13_r;
wire signed [`CalcTempBus]          temp_m1_15_13_i;
wire signed [`CalcTempBus]          temp_m1_15_14_r;
wire signed [`CalcTempBus]          temp_m1_15_14_i;
wire signed [`CalcTempBus]          temp_m1_15_15_r;
wire signed [`CalcTempBus]          temp_m1_15_15_i;
wire signed [`CalcTempBus]          temp_m1_15_16_r;
wire signed [`CalcTempBus]          temp_m1_15_16_i;
wire signed [`CalcTempBus]          temp_m1_16_1_r;
wire signed [`CalcTempBus]          temp_m1_16_1_i;
wire signed [`CalcTempBus]          temp_m1_16_2_r;
wire signed [`CalcTempBus]          temp_m1_16_2_i;
wire signed [`CalcTempBus]          temp_m1_16_3_r;
wire signed [`CalcTempBus]          temp_m1_16_3_i;
wire signed [`CalcTempBus]          temp_m1_16_4_r;
wire signed [`CalcTempBus]          temp_m1_16_4_i;
wire signed [`CalcTempBus]          temp_m1_16_5_r;
wire signed [`CalcTempBus]          temp_m1_16_5_i;
wire signed [`CalcTempBus]          temp_m1_16_6_r;
wire signed [`CalcTempBus]          temp_m1_16_6_i;
wire signed [`CalcTempBus]          temp_m1_16_7_r;
wire signed [`CalcTempBus]          temp_m1_16_7_i;
wire signed [`CalcTempBus]          temp_m1_16_8_r;
wire signed [`CalcTempBus]          temp_m1_16_8_i;
wire signed [`CalcTempBus]          temp_m1_16_9_r;
wire signed [`CalcTempBus]          temp_m1_16_9_i;
wire signed [`CalcTempBus]          temp_m1_16_10_r;
wire signed [`CalcTempBus]          temp_m1_16_10_i;
wire signed [`CalcTempBus]          temp_m1_16_11_r;
wire signed [`CalcTempBus]          temp_m1_16_11_i;
wire signed [`CalcTempBus]          temp_m1_16_12_r;
wire signed [`CalcTempBus]          temp_m1_16_12_i;
wire signed [`CalcTempBus]          temp_m1_16_13_r;
wire signed [`CalcTempBus]          temp_m1_16_13_i;
wire signed [`CalcTempBus]          temp_m1_16_14_r;
wire signed [`CalcTempBus]          temp_m1_16_14_i;
wire signed [`CalcTempBus]          temp_m1_16_15_r;
wire signed [`CalcTempBus]          temp_m1_16_15_i;
wire signed [`CalcTempBus]          temp_m1_16_16_r;
wire signed [`CalcTempBus]          temp_m1_16_16_i;
wire signed [`CalcTempBus]          temp_m2_1_1_r;
wire signed [`CalcTempBus]          temp_m2_1_1_i;
wire signed [`CalcTempBus]          temp_m2_1_2_r;
wire signed [`CalcTempBus]          temp_m2_1_2_i;
wire signed [`CalcTempBus]          temp_m2_1_3_r;
wire signed [`CalcTempBus]          temp_m2_1_3_i;
wire signed [`CalcTempBus]          temp_m2_1_4_r;
wire signed [`CalcTempBus]          temp_m2_1_4_i;
wire signed [`CalcTempBus]          temp_m2_1_5_r;
wire signed [`CalcTempBus]          temp_m2_1_5_i;
wire signed [`CalcTempBus]          temp_m2_1_6_r;
wire signed [`CalcTempBus]          temp_m2_1_6_i;
wire signed [`CalcTempBus]          temp_m2_1_7_r;
wire signed [`CalcTempBus]          temp_m2_1_7_i;
wire signed [`CalcTempBus]          temp_m2_1_8_r;
wire signed [`CalcTempBus]          temp_m2_1_8_i;
wire signed [`CalcTempBus]          temp_m2_1_9_r;
wire signed [`CalcTempBus]          temp_m2_1_9_i;
wire signed [`CalcTempBus]          temp_m2_1_10_r;
wire signed [`CalcTempBus]          temp_m2_1_10_i;
wire signed [`CalcTempBus]          temp_m2_1_11_r;
wire signed [`CalcTempBus]          temp_m2_1_11_i;
wire signed [`CalcTempBus]          temp_m2_1_12_r;
wire signed [`CalcTempBus]          temp_m2_1_12_i;
wire signed [`CalcTempBus]          temp_m2_1_13_r;
wire signed [`CalcTempBus]          temp_m2_1_13_i;
wire signed [`CalcTempBus]          temp_m2_1_14_r;
wire signed [`CalcTempBus]          temp_m2_1_14_i;
wire signed [`CalcTempBus]          temp_m2_1_15_r;
wire signed [`CalcTempBus]          temp_m2_1_15_i;
wire signed [`CalcTempBus]          temp_m2_1_16_r;
wire signed [`CalcTempBus]          temp_m2_1_16_i;
wire signed [`CalcTempBus]          temp_m2_2_1_r;
wire signed [`CalcTempBus]          temp_m2_2_1_i;
wire signed [`CalcTempBus]          temp_m2_2_2_r;
wire signed [`CalcTempBus]          temp_m2_2_2_i;
wire signed [`CalcTempBus]          temp_m2_2_3_r;
wire signed [`CalcTempBus]          temp_m2_2_3_i;
wire signed [`CalcTempBus]          temp_m2_2_4_r;
wire signed [`CalcTempBus]          temp_m2_2_4_i;
wire signed [`CalcTempBus]          temp_m2_2_5_r;
wire signed [`CalcTempBus]          temp_m2_2_5_i;
wire signed [`CalcTempBus]          temp_m2_2_6_r;
wire signed [`CalcTempBus]          temp_m2_2_6_i;
wire signed [`CalcTempBus]          temp_m2_2_7_r;
wire signed [`CalcTempBus]          temp_m2_2_7_i;
wire signed [`CalcTempBus]          temp_m2_2_8_r;
wire signed [`CalcTempBus]          temp_m2_2_8_i;
wire signed [`CalcTempBus]          temp_m2_2_9_r;
wire signed [`CalcTempBus]          temp_m2_2_9_i;
wire signed [`CalcTempBus]          temp_m2_2_10_r;
wire signed [`CalcTempBus]          temp_m2_2_10_i;
wire signed [`CalcTempBus]          temp_m2_2_11_r;
wire signed [`CalcTempBus]          temp_m2_2_11_i;
wire signed [`CalcTempBus]          temp_m2_2_12_r;
wire signed [`CalcTempBus]          temp_m2_2_12_i;
wire signed [`CalcTempBus]          temp_m2_2_13_r;
wire signed [`CalcTempBus]          temp_m2_2_13_i;
wire signed [`CalcTempBus]          temp_m2_2_14_r;
wire signed [`CalcTempBus]          temp_m2_2_14_i;
wire signed [`CalcTempBus]          temp_m2_2_15_r;
wire signed [`CalcTempBus]          temp_m2_2_15_i;
wire signed [`CalcTempBus]          temp_m2_2_16_r;
wire signed [`CalcTempBus]          temp_m2_2_16_i;
wire signed [`CalcTempBus]          temp_m2_3_1_r;
wire signed [`CalcTempBus]          temp_m2_3_1_i;
wire signed [`CalcTempBus]          temp_m2_3_2_r;
wire signed [`CalcTempBus]          temp_m2_3_2_i;
wire signed [`CalcTempBus]          temp_m2_3_3_r;
wire signed [`CalcTempBus]          temp_m2_3_3_i;
wire signed [`CalcTempBus]          temp_m2_3_4_r;
wire signed [`CalcTempBus]          temp_m2_3_4_i;
wire signed [`CalcTempBus]          temp_m2_3_5_r;
wire signed [`CalcTempBus]          temp_m2_3_5_i;
wire signed [`CalcTempBus]          temp_m2_3_6_r;
wire signed [`CalcTempBus]          temp_m2_3_6_i;
wire signed [`CalcTempBus]          temp_m2_3_7_r;
wire signed [`CalcTempBus]          temp_m2_3_7_i;
wire signed [`CalcTempBus]          temp_m2_3_8_r;
wire signed [`CalcTempBus]          temp_m2_3_8_i;
wire signed [`CalcTempBus]          temp_m2_3_9_r;
wire signed [`CalcTempBus]          temp_m2_3_9_i;
wire signed [`CalcTempBus]          temp_m2_3_10_r;
wire signed [`CalcTempBus]          temp_m2_3_10_i;
wire signed [`CalcTempBus]          temp_m2_3_11_r;
wire signed [`CalcTempBus]          temp_m2_3_11_i;
wire signed [`CalcTempBus]          temp_m2_3_12_r;
wire signed [`CalcTempBus]          temp_m2_3_12_i;
wire signed [`CalcTempBus]          temp_m2_3_13_r;
wire signed [`CalcTempBus]          temp_m2_3_13_i;
wire signed [`CalcTempBus]          temp_m2_3_14_r;
wire signed [`CalcTempBus]          temp_m2_3_14_i;
wire signed [`CalcTempBus]          temp_m2_3_15_r;
wire signed [`CalcTempBus]          temp_m2_3_15_i;
wire signed [`CalcTempBus]          temp_m2_3_16_r;
wire signed [`CalcTempBus]          temp_m2_3_16_i;
wire signed [`CalcTempBus]          temp_m2_4_1_r;
wire signed [`CalcTempBus]          temp_m2_4_1_i;
wire signed [`CalcTempBus]          temp_m2_4_2_r;
wire signed [`CalcTempBus]          temp_m2_4_2_i;
wire signed [`CalcTempBus]          temp_m2_4_3_r;
wire signed [`CalcTempBus]          temp_m2_4_3_i;
wire signed [`CalcTempBus]          temp_m2_4_4_r;
wire signed [`CalcTempBus]          temp_m2_4_4_i;
wire signed [`CalcTempBus]          temp_m2_4_5_r;
wire signed [`CalcTempBus]          temp_m2_4_5_i;
wire signed [`CalcTempBus]          temp_m2_4_6_r;
wire signed [`CalcTempBus]          temp_m2_4_6_i;
wire signed [`CalcTempBus]          temp_m2_4_7_r;
wire signed [`CalcTempBus]          temp_m2_4_7_i;
wire signed [`CalcTempBus]          temp_m2_4_8_r;
wire signed [`CalcTempBus]          temp_m2_4_8_i;
wire signed [`CalcTempBus]          temp_m2_4_9_r;
wire signed [`CalcTempBus]          temp_m2_4_9_i;
wire signed [`CalcTempBus]          temp_m2_4_10_r;
wire signed [`CalcTempBus]          temp_m2_4_10_i;
wire signed [`CalcTempBus]          temp_m2_4_11_r;
wire signed [`CalcTempBus]          temp_m2_4_11_i;
wire signed [`CalcTempBus]          temp_m2_4_12_r;
wire signed [`CalcTempBus]          temp_m2_4_12_i;
wire signed [`CalcTempBus]          temp_m2_4_13_r;
wire signed [`CalcTempBus]          temp_m2_4_13_i;
wire signed [`CalcTempBus]          temp_m2_4_14_r;
wire signed [`CalcTempBus]          temp_m2_4_14_i;
wire signed [`CalcTempBus]          temp_m2_4_15_r;
wire signed [`CalcTempBus]          temp_m2_4_15_i;
wire signed [`CalcTempBus]          temp_m2_4_16_r;
wire signed [`CalcTempBus]          temp_m2_4_16_i;
wire signed [`CalcTempBus]          temp_m2_5_1_r;
wire signed [`CalcTempBus]          temp_m2_5_1_i;
wire signed [`CalcTempBus]          temp_m2_5_2_r;
wire signed [`CalcTempBus]          temp_m2_5_2_i;
wire signed [`CalcTempBus]          temp_m2_5_3_r;
wire signed [`CalcTempBus]          temp_m2_5_3_i;
wire signed [`CalcTempBus]          temp_m2_5_4_r;
wire signed [`CalcTempBus]          temp_m2_5_4_i;
wire signed [`CalcTempBus]          temp_m2_5_5_r;
wire signed [`CalcTempBus]          temp_m2_5_5_i;
wire signed [`CalcTempBus]          temp_m2_5_6_r;
wire signed [`CalcTempBus]          temp_m2_5_6_i;
wire signed [`CalcTempBus]          temp_m2_5_7_r;
wire signed [`CalcTempBus]          temp_m2_5_7_i;
wire signed [`CalcTempBus]          temp_m2_5_8_r;
wire signed [`CalcTempBus]          temp_m2_5_8_i;
wire signed [`CalcTempBus]          temp_m2_5_9_r;
wire signed [`CalcTempBus]          temp_m2_5_9_i;
wire signed [`CalcTempBus]          temp_m2_5_10_r;
wire signed [`CalcTempBus]          temp_m2_5_10_i;
wire signed [`CalcTempBus]          temp_m2_5_11_r;
wire signed [`CalcTempBus]          temp_m2_5_11_i;
wire signed [`CalcTempBus]          temp_m2_5_12_r;
wire signed [`CalcTempBus]          temp_m2_5_12_i;
wire signed [`CalcTempBus]          temp_m2_5_13_r;
wire signed [`CalcTempBus]          temp_m2_5_13_i;
wire signed [`CalcTempBus]          temp_m2_5_14_r;
wire signed [`CalcTempBus]          temp_m2_5_14_i;
wire signed [`CalcTempBus]          temp_m2_5_15_r;
wire signed [`CalcTempBus]          temp_m2_5_15_i;
wire signed [`CalcTempBus]          temp_m2_5_16_r;
wire signed [`CalcTempBus]          temp_m2_5_16_i;
wire signed [`CalcTempBus]          temp_m2_6_1_r;
wire signed [`CalcTempBus]          temp_m2_6_1_i;
wire signed [`CalcTempBus]          temp_m2_6_2_r;
wire signed [`CalcTempBus]          temp_m2_6_2_i;
wire signed [`CalcTempBus]          temp_m2_6_3_r;
wire signed [`CalcTempBus]          temp_m2_6_3_i;
wire signed [`CalcTempBus]          temp_m2_6_4_r;
wire signed [`CalcTempBus]          temp_m2_6_4_i;
wire signed [`CalcTempBus]          temp_m2_6_5_r;
wire signed [`CalcTempBus]          temp_m2_6_5_i;
wire signed [`CalcTempBus]          temp_m2_6_6_r;
wire signed [`CalcTempBus]          temp_m2_6_6_i;
wire signed [`CalcTempBus]          temp_m2_6_7_r;
wire signed [`CalcTempBus]          temp_m2_6_7_i;
wire signed [`CalcTempBus]          temp_m2_6_8_r;
wire signed [`CalcTempBus]          temp_m2_6_8_i;
wire signed [`CalcTempBus]          temp_m2_6_9_r;
wire signed [`CalcTempBus]          temp_m2_6_9_i;
wire signed [`CalcTempBus]          temp_m2_6_10_r;
wire signed [`CalcTempBus]          temp_m2_6_10_i;
wire signed [`CalcTempBus]          temp_m2_6_11_r;
wire signed [`CalcTempBus]          temp_m2_6_11_i;
wire signed [`CalcTempBus]          temp_m2_6_12_r;
wire signed [`CalcTempBus]          temp_m2_6_12_i;
wire signed [`CalcTempBus]          temp_m2_6_13_r;
wire signed [`CalcTempBus]          temp_m2_6_13_i;
wire signed [`CalcTempBus]          temp_m2_6_14_r;
wire signed [`CalcTempBus]          temp_m2_6_14_i;
wire signed [`CalcTempBus]          temp_m2_6_15_r;
wire signed [`CalcTempBus]          temp_m2_6_15_i;
wire signed [`CalcTempBus]          temp_m2_6_16_r;
wire signed [`CalcTempBus]          temp_m2_6_16_i;
wire signed [`CalcTempBus]          temp_m2_7_1_r;
wire signed [`CalcTempBus]          temp_m2_7_1_i;
wire signed [`CalcTempBus]          temp_m2_7_2_r;
wire signed [`CalcTempBus]          temp_m2_7_2_i;
wire signed [`CalcTempBus]          temp_m2_7_3_r;
wire signed [`CalcTempBus]          temp_m2_7_3_i;
wire signed [`CalcTempBus]          temp_m2_7_4_r;
wire signed [`CalcTempBus]          temp_m2_7_4_i;
wire signed [`CalcTempBus]          temp_m2_7_5_r;
wire signed [`CalcTempBus]          temp_m2_7_5_i;
wire signed [`CalcTempBus]          temp_m2_7_6_r;
wire signed [`CalcTempBus]          temp_m2_7_6_i;
wire signed [`CalcTempBus]          temp_m2_7_7_r;
wire signed [`CalcTempBus]          temp_m2_7_7_i;
wire signed [`CalcTempBus]          temp_m2_7_8_r;
wire signed [`CalcTempBus]          temp_m2_7_8_i;
wire signed [`CalcTempBus]          temp_m2_7_9_r;
wire signed [`CalcTempBus]          temp_m2_7_9_i;
wire signed [`CalcTempBus]          temp_m2_7_10_r;
wire signed [`CalcTempBus]          temp_m2_7_10_i;
wire signed [`CalcTempBus]          temp_m2_7_11_r;
wire signed [`CalcTempBus]          temp_m2_7_11_i;
wire signed [`CalcTempBus]          temp_m2_7_12_r;
wire signed [`CalcTempBus]          temp_m2_7_12_i;
wire signed [`CalcTempBus]          temp_m2_7_13_r;
wire signed [`CalcTempBus]          temp_m2_7_13_i;
wire signed [`CalcTempBus]          temp_m2_7_14_r;
wire signed [`CalcTempBus]          temp_m2_7_14_i;
wire signed [`CalcTempBus]          temp_m2_7_15_r;
wire signed [`CalcTempBus]          temp_m2_7_15_i;
wire signed [`CalcTempBus]          temp_m2_7_16_r;
wire signed [`CalcTempBus]          temp_m2_7_16_i;
wire signed [`CalcTempBus]          temp_m2_8_1_r;
wire signed [`CalcTempBus]          temp_m2_8_1_i;
wire signed [`CalcTempBus]          temp_m2_8_2_r;
wire signed [`CalcTempBus]          temp_m2_8_2_i;
wire signed [`CalcTempBus]          temp_m2_8_3_r;
wire signed [`CalcTempBus]          temp_m2_8_3_i;
wire signed [`CalcTempBus]          temp_m2_8_4_r;
wire signed [`CalcTempBus]          temp_m2_8_4_i;
wire signed [`CalcTempBus]          temp_m2_8_5_r;
wire signed [`CalcTempBus]          temp_m2_8_5_i;
wire signed [`CalcTempBus]          temp_m2_8_6_r;
wire signed [`CalcTempBus]          temp_m2_8_6_i;
wire signed [`CalcTempBus]          temp_m2_8_7_r;
wire signed [`CalcTempBus]          temp_m2_8_7_i;
wire signed [`CalcTempBus]          temp_m2_8_8_r;
wire signed [`CalcTempBus]          temp_m2_8_8_i;
wire signed [`CalcTempBus]          temp_m2_8_9_r;
wire signed [`CalcTempBus]          temp_m2_8_9_i;
wire signed [`CalcTempBus]          temp_m2_8_10_r;
wire signed [`CalcTempBus]          temp_m2_8_10_i;
wire signed [`CalcTempBus]          temp_m2_8_11_r;
wire signed [`CalcTempBus]          temp_m2_8_11_i;
wire signed [`CalcTempBus]          temp_m2_8_12_r;
wire signed [`CalcTempBus]          temp_m2_8_12_i;
wire signed [`CalcTempBus]          temp_m2_8_13_r;
wire signed [`CalcTempBus]          temp_m2_8_13_i;
wire signed [`CalcTempBus]          temp_m2_8_14_r;
wire signed [`CalcTempBus]          temp_m2_8_14_i;
wire signed [`CalcTempBus]          temp_m2_8_15_r;
wire signed [`CalcTempBus]          temp_m2_8_15_i;
wire signed [`CalcTempBus]          temp_m2_8_16_r;
wire signed [`CalcTempBus]          temp_m2_8_16_i;
wire signed [`CalcTempBus]          temp_m2_9_1_r;
wire signed [`CalcTempBus]          temp_m2_9_1_i;
wire signed [`CalcTempBus]          temp_m2_9_2_r;
wire signed [`CalcTempBus]          temp_m2_9_2_i;
wire signed [`CalcTempBus]          temp_m2_9_3_r;
wire signed [`CalcTempBus]          temp_m2_9_3_i;
wire signed [`CalcTempBus]          temp_m2_9_4_r;
wire signed [`CalcTempBus]          temp_m2_9_4_i;
wire signed [`CalcTempBus]          temp_m2_9_5_r;
wire signed [`CalcTempBus]          temp_m2_9_5_i;
wire signed [`CalcTempBus]          temp_m2_9_6_r;
wire signed [`CalcTempBus]          temp_m2_9_6_i;
wire signed [`CalcTempBus]          temp_m2_9_7_r;
wire signed [`CalcTempBus]          temp_m2_9_7_i;
wire signed [`CalcTempBus]          temp_m2_9_8_r;
wire signed [`CalcTempBus]          temp_m2_9_8_i;
wire signed [`CalcTempBus]          temp_m2_9_9_r;
wire signed [`CalcTempBus]          temp_m2_9_9_i;
wire signed [`CalcTempBus]          temp_m2_9_10_r;
wire signed [`CalcTempBus]          temp_m2_9_10_i;
wire signed [`CalcTempBus]          temp_m2_9_11_r;
wire signed [`CalcTempBus]          temp_m2_9_11_i;
wire signed [`CalcTempBus]          temp_m2_9_12_r;
wire signed [`CalcTempBus]          temp_m2_9_12_i;
wire signed [`CalcTempBus]          temp_m2_9_13_r;
wire signed [`CalcTempBus]          temp_m2_9_13_i;
wire signed [`CalcTempBus]          temp_m2_9_14_r;
wire signed [`CalcTempBus]          temp_m2_9_14_i;
wire signed [`CalcTempBus]          temp_m2_9_15_r;
wire signed [`CalcTempBus]          temp_m2_9_15_i;
wire signed [`CalcTempBus]          temp_m2_9_16_r;
wire signed [`CalcTempBus]          temp_m2_9_16_i;
wire signed [`CalcTempBus]          temp_m2_10_1_r;
wire signed [`CalcTempBus]          temp_m2_10_1_i;
wire signed [`CalcTempBus]          temp_m2_10_2_r;
wire signed [`CalcTempBus]          temp_m2_10_2_i;
wire signed [`CalcTempBus]          temp_m2_10_3_r;
wire signed [`CalcTempBus]          temp_m2_10_3_i;
wire signed [`CalcTempBus]          temp_m2_10_4_r;
wire signed [`CalcTempBus]          temp_m2_10_4_i;
wire signed [`CalcTempBus]          temp_m2_10_5_r;
wire signed [`CalcTempBus]          temp_m2_10_5_i;
wire signed [`CalcTempBus]          temp_m2_10_6_r;
wire signed [`CalcTempBus]          temp_m2_10_6_i;
wire signed [`CalcTempBus]          temp_m2_10_7_r;
wire signed [`CalcTempBus]          temp_m2_10_7_i;
wire signed [`CalcTempBus]          temp_m2_10_8_r;
wire signed [`CalcTempBus]          temp_m2_10_8_i;
wire signed [`CalcTempBus]          temp_m2_10_9_r;
wire signed [`CalcTempBus]          temp_m2_10_9_i;
wire signed [`CalcTempBus]          temp_m2_10_10_r;
wire signed [`CalcTempBus]          temp_m2_10_10_i;
wire signed [`CalcTempBus]          temp_m2_10_11_r;
wire signed [`CalcTempBus]          temp_m2_10_11_i;
wire signed [`CalcTempBus]          temp_m2_10_12_r;
wire signed [`CalcTempBus]          temp_m2_10_12_i;
wire signed [`CalcTempBus]          temp_m2_10_13_r;
wire signed [`CalcTempBus]          temp_m2_10_13_i;
wire signed [`CalcTempBus]          temp_m2_10_14_r;
wire signed [`CalcTempBus]          temp_m2_10_14_i;
wire signed [`CalcTempBus]          temp_m2_10_15_r;
wire signed [`CalcTempBus]          temp_m2_10_15_i;
wire signed [`CalcTempBus]          temp_m2_10_16_r;
wire signed [`CalcTempBus]          temp_m2_10_16_i;
wire signed [`CalcTempBus]          temp_m2_11_1_r;
wire signed [`CalcTempBus]          temp_m2_11_1_i;
wire signed [`CalcTempBus]          temp_m2_11_2_r;
wire signed [`CalcTempBus]          temp_m2_11_2_i;
wire signed [`CalcTempBus]          temp_m2_11_3_r;
wire signed [`CalcTempBus]          temp_m2_11_3_i;
wire signed [`CalcTempBus]          temp_m2_11_4_r;
wire signed [`CalcTempBus]          temp_m2_11_4_i;
wire signed [`CalcTempBus]          temp_m2_11_5_r;
wire signed [`CalcTempBus]          temp_m2_11_5_i;
wire signed [`CalcTempBus]          temp_m2_11_6_r;
wire signed [`CalcTempBus]          temp_m2_11_6_i;
wire signed [`CalcTempBus]          temp_m2_11_7_r;
wire signed [`CalcTempBus]          temp_m2_11_7_i;
wire signed [`CalcTempBus]          temp_m2_11_8_r;
wire signed [`CalcTempBus]          temp_m2_11_8_i;
wire signed [`CalcTempBus]          temp_m2_11_9_r;
wire signed [`CalcTempBus]          temp_m2_11_9_i;
wire signed [`CalcTempBus]          temp_m2_11_10_r;
wire signed [`CalcTempBus]          temp_m2_11_10_i;
wire signed [`CalcTempBus]          temp_m2_11_11_r;
wire signed [`CalcTempBus]          temp_m2_11_11_i;
wire signed [`CalcTempBus]          temp_m2_11_12_r;
wire signed [`CalcTempBus]          temp_m2_11_12_i;
wire signed [`CalcTempBus]          temp_m2_11_13_r;
wire signed [`CalcTempBus]          temp_m2_11_13_i;
wire signed [`CalcTempBus]          temp_m2_11_14_r;
wire signed [`CalcTempBus]          temp_m2_11_14_i;
wire signed [`CalcTempBus]          temp_m2_11_15_r;
wire signed [`CalcTempBus]          temp_m2_11_15_i;
wire signed [`CalcTempBus]          temp_m2_11_16_r;
wire signed [`CalcTempBus]          temp_m2_11_16_i;
wire signed [`CalcTempBus]          temp_m2_12_1_r;
wire signed [`CalcTempBus]          temp_m2_12_1_i;
wire signed [`CalcTempBus]          temp_m2_12_2_r;
wire signed [`CalcTempBus]          temp_m2_12_2_i;
wire signed [`CalcTempBus]          temp_m2_12_3_r;
wire signed [`CalcTempBus]          temp_m2_12_3_i;
wire signed [`CalcTempBus]          temp_m2_12_4_r;
wire signed [`CalcTempBus]          temp_m2_12_4_i;
wire signed [`CalcTempBus]          temp_m2_12_5_r;
wire signed [`CalcTempBus]          temp_m2_12_5_i;
wire signed [`CalcTempBus]          temp_m2_12_6_r;
wire signed [`CalcTempBus]          temp_m2_12_6_i;
wire signed [`CalcTempBus]          temp_m2_12_7_r;
wire signed [`CalcTempBus]          temp_m2_12_7_i;
wire signed [`CalcTempBus]          temp_m2_12_8_r;
wire signed [`CalcTempBus]          temp_m2_12_8_i;
wire signed [`CalcTempBus]          temp_m2_12_9_r;
wire signed [`CalcTempBus]          temp_m2_12_9_i;
wire signed [`CalcTempBus]          temp_m2_12_10_r;
wire signed [`CalcTempBus]          temp_m2_12_10_i;
wire signed [`CalcTempBus]          temp_m2_12_11_r;
wire signed [`CalcTempBus]          temp_m2_12_11_i;
wire signed [`CalcTempBus]          temp_m2_12_12_r;
wire signed [`CalcTempBus]          temp_m2_12_12_i;
wire signed [`CalcTempBus]          temp_m2_12_13_r;
wire signed [`CalcTempBus]          temp_m2_12_13_i;
wire signed [`CalcTempBus]          temp_m2_12_14_r;
wire signed [`CalcTempBus]          temp_m2_12_14_i;
wire signed [`CalcTempBus]          temp_m2_12_15_r;
wire signed [`CalcTempBus]          temp_m2_12_15_i;
wire signed [`CalcTempBus]          temp_m2_12_16_r;
wire signed [`CalcTempBus]          temp_m2_12_16_i;
wire signed [`CalcTempBus]          temp_m2_13_1_r;
wire signed [`CalcTempBus]          temp_m2_13_1_i;
wire signed [`CalcTempBus]          temp_m2_13_2_r;
wire signed [`CalcTempBus]          temp_m2_13_2_i;
wire signed [`CalcTempBus]          temp_m2_13_3_r;
wire signed [`CalcTempBus]          temp_m2_13_3_i;
wire signed [`CalcTempBus]          temp_m2_13_4_r;
wire signed [`CalcTempBus]          temp_m2_13_4_i;
wire signed [`CalcTempBus]          temp_m2_13_5_r;
wire signed [`CalcTempBus]          temp_m2_13_5_i;
wire signed [`CalcTempBus]          temp_m2_13_6_r;
wire signed [`CalcTempBus]          temp_m2_13_6_i;
wire signed [`CalcTempBus]          temp_m2_13_7_r;
wire signed [`CalcTempBus]          temp_m2_13_7_i;
wire signed [`CalcTempBus]          temp_m2_13_8_r;
wire signed [`CalcTempBus]          temp_m2_13_8_i;
wire signed [`CalcTempBus]          temp_m2_13_9_r;
wire signed [`CalcTempBus]          temp_m2_13_9_i;
wire signed [`CalcTempBus]          temp_m2_13_10_r;
wire signed [`CalcTempBus]          temp_m2_13_10_i;
wire signed [`CalcTempBus]          temp_m2_13_11_r;
wire signed [`CalcTempBus]          temp_m2_13_11_i;
wire signed [`CalcTempBus]          temp_m2_13_12_r;
wire signed [`CalcTempBus]          temp_m2_13_12_i;
wire signed [`CalcTempBus]          temp_m2_13_13_r;
wire signed [`CalcTempBus]          temp_m2_13_13_i;
wire signed [`CalcTempBus]          temp_m2_13_14_r;
wire signed [`CalcTempBus]          temp_m2_13_14_i;
wire signed [`CalcTempBus]          temp_m2_13_15_r;
wire signed [`CalcTempBus]          temp_m2_13_15_i;
wire signed [`CalcTempBus]          temp_m2_13_16_r;
wire signed [`CalcTempBus]          temp_m2_13_16_i;
wire signed [`CalcTempBus]          temp_m2_14_1_r;
wire signed [`CalcTempBus]          temp_m2_14_1_i;
wire signed [`CalcTempBus]          temp_m2_14_2_r;
wire signed [`CalcTempBus]          temp_m2_14_2_i;
wire signed [`CalcTempBus]          temp_m2_14_3_r;
wire signed [`CalcTempBus]          temp_m2_14_3_i;
wire signed [`CalcTempBus]          temp_m2_14_4_r;
wire signed [`CalcTempBus]          temp_m2_14_4_i;
wire signed [`CalcTempBus]          temp_m2_14_5_r;
wire signed [`CalcTempBus]          temp_m2_14_5_i;
wire signed [`CalcTempBus]          temp_m2_14_6_r;
wire signed [`CalcTempBus]          temp_m2_14_6_i;
wire signed [`CalcTempBus]          temp_m2_14_7_r;
wire signed [`CalcTempBus]          temp_m2_14_7_i;
wire signed [`CalcTempBus]          temp_m2_14_8_r;
wire signed [`CalcTempBus]          temp_m2_14_8_i;
wire signed [`CalcTempBus]          temp_m2_14_9_r;
wire signed [`CalcTempBus]          temp_m2_14_9_i;
wire signed [`CalcTempBus]          temp_m2_14_10_r;
wire signed [`CalcTempBus]          temp_m2_14_10_i;
wire signed [`CalcTempBus]          temp_m2_14_11_r;
wire signed [`CalcTempBus]          temp_m2_14_11_i;
wire signed [`CalcTempBus]          temp_m2_14_12_r;
wire signed [`CalcTempBus]          temp_m2_14_12_i;
wire signed [`CalcTempBus]          temp_m2_14_13_r;
wire signed [`CalcTempBus]          temp_m2_14_13_i;
wire signed [`CalcTempBus]          temp_m2_14_14_r;
wire signed [`CalcTempBus]          temp_m2_14_14_i;
wire signed [`CalcTempBus]          temp_m2_14_15_r;
wire signed [`CalcTempBus]          temp_m2_14_15_i;
wire signed [`CalcTempBus]          temp_m2_14_16_r;
wire signed [`CalcTempBus]          temp_m2_14_16_i;
wire signed [`CalcTempBus]          temp_m2_15_1_r;
wire signed [`CalcTempBus]          temp_m2_15_1_i;
wire signed [`CalcTempBus]          temp_m2_15_2_r;
wire signed [`CalcTempBus]          temp_m2_15_2_i;
wire signed [`CalcTempBus]          temp_m2_15_3_r;
wire signed [`CalcTempBus]          temp_m2_15_3_i;
wire signed [`CalcTempBus]          temp_m2_15_4_r;
wire signed [`CalcTempBus]          temp_m2_15_4_i;
wire signed [`CalcTempBus]          temp_m2_15_5_r;
wire signed [`CalcTempBus]          temp_m2_15_5_i;
wire signed [`CalcTempBus]          temp_m2_15_6_r;
wire signed [`CalcTempBus]          temp_m2_15_6_i;
wire signed [`CalcTempBus]          temp_m2_15_7_r;
wire signed [`CalcTempBus]          temp_m2_15_7_i;
wire signed [`CalcTempBus]          temp_m2_15_8_r;
wire signed [`CalcTempBus]          temp_m2_15_8_i;
wire signed [`CalcTempBus]          temp_m2_15_9_r;
wire signed [`CalcTempBus]          temp_m2_15_9_i;
wire signed [`CalcTempBus]          temp_m2_15_10_r;
wire signed [`CalcTempBus]          temp_m2_15_10_i;
wire signed [`CalcTempBus]          temp_m2_15_11_r;
wire signed [`CalcTempBus]          temp_m2_15_11_i;
wire signed [`CalcTempBus]          temp_m2_15_12_r;
wire signed [`CalcTempBus]          temp_m2_15_12_i;
wire signed [`CalcTempBus]          temp_m2_15_13_r;
wire signed [`CalcTempBus]          temp_m2_15_13_i;
wire signed [`CalcTempBus]          temp_m2_15_14_r;
wire signed [`CalcTempBus]          temp_m2_15_14_i;
wire signed [`CalcTempBus]          temp_m2_15_15_r;
wire signed [`CalcTempBus]          temp_m2_15_15_i;
wire signed [`CalcTempBus]          temp_m2_15_16_r;
wire signed [`CalcTempBus]          temp_m2_15_16_i;
wire signed [`CalcTempBus]          temp_m2_16_1_r;
wire signed [`CalcTempBus]          temp_m2_16_1_i;
wire signed [`CalcTempBus]          temp_m2_16_2_r;
wire signed [`CalcTempBus]          temp_m2_16_2_i;
wire signed [`CalcTempBus]          temp_m2_16_3_r;
wire signed [`CalcTempBus]          temp_m2_16_3_i;
wire signed [`CalcTempBus]          temp_m2_16_4_r;
wire signed [`CalcTempBus]          temp_m2_16_4_i;
wire signed [`CalcTempBus]          temp_m2_16_5_r;
wire signed [`CalcTempBus]          temp_m2_16_5_i;
wire signed [`CalcTempBus]          temp_m2_16_6_r;
wire signed [`CalcTempBus]          temp_m2_16_6_i;
wire signed [`CalcTempBus]          temp_m2_16_7_r;
wire signed [`CalcTempBus]          temp_m2_16_7_i;
wire signed [`CalcTempBus]          temp_m2_16_8_r;
wire signed [`CalcTempBus]          temp_m2_16_8_i;
wire signed [`CalcTempBus]          temp_m2_16_9_r;
wire signed [`CalcTempBus]          temp_m2_16_9_i;
wire signed [`CalcTempBus]          temp_m2_16_10_r;
wire signed [`CalcTempBus]          temp_m2_16_10_i;
wire signed [`CalcTempBus]          temp_m2_16_11_r;
wire signed [`CalcTempBus]          temp_m2_16_11_i;
wire signed [`CalcTempBus]          temp_m2_16_12_r;
wire signed [`CalcTempBus]          temp_m2_16_12_i;
wire signed [`CalcTempBus]          temp_m2_16_13_r;
wire signed [`CalcTempBus]          temp_m2_16_13_i;
wire signed [`CalcTempBus]          temp_m2_16_14_r;
wire signed [`CalcTempBus]          temp_m2_16_14_i;
wire signed [`CalcTempBus]          temp_m2_16_15_r;
wire signed [`CalcTempBus]          temp_m2_16_15_i;
wire signed [`CalcTempBus]          temp_m2_16_16_r;
wire signed [`CalcTempBus]          temp_m2_16_16_i;
wire signed [`CalcTempBus]          temp_m3_1_1_r;
wire signed [`CalcTempBus]          temp_m3_1_1_i;
wire signed [`CalcTempBus]          temp_m3_1_2_r;
wire signed [`CalcTempBus]          temp_m3_1_2_i;
wire signed [`CalcTempBus]          temp_m3_1_3_r;
wire signed [`CalcTempBus]          temp_m3_1_3_i;
wire signed [`CalcTempBus]          temp_m3_1_4_r;
wire signed [`CalcTempBus]          temp_m3_1_4_i;
wire signed [`CalcTempBus]          temp_m3_1_5_r;
wire signed [`CalcTempBus]          temp_m3_1_5_i;
wire signed [`CalcTempBus]          temp_m3_1_6_r;
wire signed [`CalcTempBus]          temp_m3_1_6_i;
wire signed [`CalcTempBus]          temp_m3_1_7_r;
wire signed [`CalcTempBus]          temp_m3_1_7_i;
wire signed [`CalcTempBus]          temp_m3_1_8_r;
wire signed [`CalcTempBus]          temp_m3_1_8_i;
wire signed [`CalcTempBus]          temp_m3_1_9_r;
wire signed [`CalcTempBus]          temp_m3_1_9_i;
wire signed [`CalcTempBus]          temp_m3_1_10_r;
wire signed [`CalcTempBus]          temp_m3_1_10_i;
wire signed [`CalcTempBus]          temp_m3_1_11_r;
wire signed [`CalcTempBus]          temp_m3_1_11_i;
wire signed [`CalcTempBus]          temp_m3_1_12_r;
wire signed [`CalcTempBus]          temp_m3_1_12_i;
wire signed [`CalcTempBus]          temp_m3_1_13_r;
wire signed [`CalcTempBus]          temp_m3_1_13_i;
wire signed [`CalcTempBus]          temp_m3_1_14_r;
wire signed [`CalcTempBus]          temp_m3_1_14_i;
wire signed [`CalcTempBus]          temp_m3_1_15_r;
wire signed [`CalcTempBus]          temp_m3_1_15_i;
wire signed [`CalcTempBus]          temp_m3_1_16_r;
wire signed [`CalcTempBus]          temp_m3_1_16_i;
wire signed [`CalcTempBus]          temp_m3_2_1_r;
wire signed [`CalcTempBus]          temp_m3_2_1_i;
wire signed [`CalcTempBus]          temp_m3_2_2_r;
wire signed [`CalcTempBus]          temp_m3_2_2_i;
wire signed [`CalcTempBus]          temp_m3_2_3_r;
wire signed [`CalcTempBus]          temp_m3_2_3_i;
wire signed [`CalcTempBus]          temp_m3_2_4_r;
wire signed [`CalcTempBus]          temp_m3_2_4_i;
wire signed [`CalcTempBus]          temp_m3_2_5_r;
wire signed [`CalcTempBus]          temp_m3_2_5_i;
wire signed [`CalcTempBus]          temp_m3_2_6_r;
wire signed [`CalcTempBus]          temp_m3_2_6_i;
wire signed [`CalcTempBus]          temp_m3_2_7_r;
wire signed [`CalcTempBus]          temp_m3_2_7_i;
wire signed [`CalcTempBus]          temp_m3_2_8_r;
wire signed [`CalcTempBus]          temp_m3_2_8_i;
wire signed [`CalcTempBus]          temp_m3_2_9_r;
wire signed [`CalcTempBus]          temp_m3_2_9_i;
wire signed [`CalcTempBus]          temp_m3_2_10_r;
wire signed [`CalcTempBus]          temp_m3_2_10_i;
wire signed [`CalcTempBus]          temp_m3_2_11_r;
wire signed [`CalcTempBus]          temp_m3_2_11_i;
wire signed [`CalcTempBus]          temp_m3_2_12_r;
wire signed [`CalcTempBus]          temp_m3_2_12_i;
wire signed [`CalcTempBus]          temp_m3_2_13_r;
wire signed [`CalcTempBus]          temp_m3_2_13_i;
wire signed [`CalcTempBus]          temp_m3_2_14_r;
wire signed [`CalcTempBus]          temp_m3_2_14_i;
wire signed [`CalcTempBus]          temp_m3_2_15_r;
wire signed [`CalcTempBus]          temp_m3_2_15_i;
wire signed [`CalcTempBus]          temp_m3_2_16_r;
wire signed [`CalcTempBus]          temp_m3_2_16_i;
wire signed [`CalcTempBus]          temp_m3_3_1_r;
wire signed [`CalcTempBus]          temp_m3_3_1_i;
wire signed [`CalcTempBus]          temp_m3_3_2_r;
wire signed [`CalcTempBus]          temp_m3_3_2_i;
wire signed [`CalcTempBus]          temp_m3_3_3_r;
wire signed [`CalcTempBus]          temp_m3_3_3_i;
wire signed [`CalcTempBus]          temp_m3_3_4_r;
wire signed [`CalcTempBus]          temp_m3_3_4_i;
wire signed [`CalcTempBus]          temp_m3_3_5_r;
wire signed [`CalcTempBus]          temp_m3_3_5_i;
wire signed [`CalcTempBus]          temp_m3_3_6_r;
wire signed [`CalcTempBus]          temp_m3_3_6_i;
wire signed [`CalcTempBus]          temp_m3_3_7_r;
wire signed [`CalcTempBus]          temp_m3_3_7_i;
wire signed [`CalcTempBus]          temp_m3_3_8_r;
wire signed [`CalcTempBus]          temp_m3_3_8_i;
wire signed [`CalcTempBus]          temp_m3_3_9_r;
wire signed [`CalcTempBus]          temp_m3_3_9_i;
wire signed [`CalcTempBus]          temp_m3_3_10_r;
wire signed [`CalcTempBus]          temp_m3_3_10_i;
wire signed [`CalcTempBus]          temp_m3_3_11_r;
wire signed [`CalcTempBus]          temp_m3_3_11_i;
wire signed [`CalcTempBus]          temp_m3_3_12_r;
wire signed [`CalcTempBus]          temp_m3_3_12_i;
wire signed [`CalcTempBus]          temp_m3_3_13_r;
wire signed [`CalcTempBus]          temp_m3_3_13_i;
wire signed [`CalcTempBus]          temp_m3_3_14_r;
wire signed [`CalcTempBus]          temp_m3_3_14_i;
wire signed [`CalcTempBus]          temp_m3_3_15_r;
wire signed [`CalcTempBus]          temp_m3_3_15_i;
wire signed [`CalcTempBus]          temp_m3_3_16_r;
wire signed [`CalcTempBus]          temp_m3_3_16_i;
wire signed [`CalcTempBus]          temp_m3_4_1_r;
wire signed [`CalcTempBus]          temp_m3_4_1_i;
wire signed [`CalcTempBus]          temp_m3_4_2_r;
wire signed [`CalcTempBus]          temp_m3_4_2_i;
wire signed [`CalcTempBus]          temp_m3_4_3_r;
wire signed [`CalcTempBus]          temp_m3_4_3_i;
wire signed [`CalcTempBus]          temp_m3_4_4_r;
wire signed [`CalcTempBus]          temp_m3_4_4_i;
wire signed [`CalcTempBus]          temp_m3_4_5_r;
wire signed [`CalcTempBus]          temp_m3_4_5_i;
wire signed [`CalcTempBus]          temp_m3_4_6_r;
wire signed [`CalcTempBus]          temp_m3_4_6_i;
wire signed [`CalcTempBus]          temp_m3_4_7_r;
wire signed [`CalcTempBus]          temp_m3_4_7_i;
wire signed [`CalcTempBus]          temp_m3_4_8_r;
wire signed [`CalcTempBus]          temp_m3_4_8_i;
wire signed [`CalcTempBus]          temp_m3_4_9_r;
wire signed [`CalcTempBus]          temp_m3_4_9_i;
wire signed [`CalcTempBus]          temp_m3_4_10_r;
wire signed [`CalcTempBus]          temp_m3_4_10_i;
wire signed [`CalcTempBus]          temp_m3_4_11_r;
wire signed [`CalcTempBus]          temp_m3_4_11_i;
wire signed [`CalcTempBus]          temp_m3_4_12_r;
wire signed [`CalcTempBus]          temp_m3_4_12_i;
wire signed [`CalcTempBus]          temp_m3_4_13_r;
wire signed [`CalcTempBus]          temp_m3_4_13_i;
wire signed [`CalcTempBus]          temp_m3_4_14_r;
wire signed [`CalcTempBus]          temp_m3_4_14_i;
wire signed [`CalcTempBus]          temp_m3_4_15_r;
wire signed [`CalcTempBus]          temp_m3_4_15_i;
wire signed [`CalcTempBus]          temp_m3_4_16_r;
wire signed [`CalcTempBus]          temp_m3_4_16_i;
wire signed [`CalcTempBus]          temp_m3_5_1_r;
wire signed [`CalcTempBus]          temp_m3_5_1_i;
wire signed [`CalcTempBus]          temp_m3_5_2_r;
wire signed [`CalcTempBus]          temp_m3_5_2_i;
wire signed [`CalcTempBus]          temp_m3_5_3_r;
wire signed [`CalcTempBus]          temp_m3_5_3_i;
wire signed [`CalcTempBus]          temp_m3_5_4_r;
wire signed [`CalcTempBus]          temp_m3_5_4_i;
wire signed [`CalcTempBus]          temp_m3_5_5_r;
wire signed [`CalcTempBus]          temp_m3_5_5_i;
wire signed [`CalcTempBus]          temp_m3_5_6_r;
wire signed [`CalcTempBus]          temp_m3_5_6_i;
wire signed [`CalcTempBus]          temp_m3_5_7_r;
wire signed [`CalcTempBus]          temp_m3_5_7_i;
wire signed [`CalcTempBus]          temp_m3_5_8_r;
wire signed [`CalcTempBus]          temp_m3_5_8_i;
wire signed [`CalcTempBus]          temp_m3_5_9_r;
wire signed [`CalcTempBus]          temp_m3_5_9_i;
wire signed [`CalcTempBus]          temp_m3_5_10_r;
wire signed [`CalcTempBus]          temp_m3_5_10_i;
wire signed [`CalcTempBus]          temp_m3_5_11_r;
wire signed [`CalcTempBus]          temp_m3_5_11_i;
wire signed [`CalcTempBus]          temp_m3_5_12_r;
wire signed [`CalcTempBus]          temp_m3_5_12_i;
wire signed [`CalcTempBus]          temp_m3_5_13_r;
wire signed [`CalcTempBus]          temp_m3_5_13_i;
wire signed [`CalcTempBus]          temp_m3_5_14_r;
wire signed [`CalcTempBus]          temp_m3_5_14_i;
wire signed [`CalcTempBus]          temp_m3_5_15_r;
wire signed [`CalcTempBus]          temp_m3_5_15_i;
wire signed [`CalcTempBus]          temp_m3_5_16_r;
wire signed [`CalcTempBus]          temp_m3_5_16_i;
wire signed [`CalcTempBus]          temp_m3_6_1_r;
wire signed [`CalcTempBus]          temp_m3_6_1_i;
wire signed [`CalcTempBus]          temp_m3_6_2_r;
wire signed [`CalcTempBus]          temp_m3_6_2_i;
wire signed [`CalcTempBus]          temp_m3_6_3_r;
wire signed [`CalcTempBus]          temp_m3_6_3_i;
wire signed [`CalcTempBus]          temp_m3_6_4_r;
wire signed [`CalcTempBus]          temp_m3_6_4_i;
wire signed [`CalcTempBus]          temp_m3_6_5_r;
wire signed [`CalcTempBus]          temp_m3_6_5_i;
wire signed [`CalcTempBus]          temp_m3_6_6_r;
wire signed [`CalcTempBus]          temp_m3_6_6_i;
wire signed [`CalcTempBus]          temp_m3_6_7_r;
wire signed [`CalcTempBus]          temp_m3_6_7_i;
wire signed [`CalcTempBus]          temp_m3_6_8_r;
wire signed [`CalcTempBus]          temp_m3_6_8_i;
wire signed [`CalcTempBus]          temp_m3_6_9_r;
wire signed [`CalcTempBus]          temp_m3_6_9_i;
wire signed [`CalcTempBus]          temp_m3_6_10_r;
wire signed [`CalcTempBus]          temp_m3_6_10_i;
wire signed [`CalcTempBus]          temp_m3_6_11_r;
wire signed [`CalcTempBus]          temp_m3_6_11_i;
wire signed [`CalcTempBus]          temp_m3_6_12_r;
wire signed [`CalcTempBus]          temp_m3_6_12_i;
wire signed [`CalcTempBus]          temp_m3_6_13_r;
wire signed [`CalcTempBus]          temp_m3_6_13_i;
wire signed [`CalcTempBus]          temp_m3_6_14_r;
wire signed [`CalcTempBus]          temp_m3_6_14_i;
wire signed [`CalcTempBus]          temp_m3_6_15_r;
wire signed [`CalcTempBus]          temp_m3_6_15_i;
wire signed [`CalcTempBus]          temp_m3_6_16_r;
wire signed [`CalcTempBus]          temp_m3_6_16_i;
wire signed [`CalcTempBus]          temp_m3_7_1_r;
wire signed [`CalcTempBus]          temp_m3_7_1_i;
wire signed [`CalcTempBus]          temp_m3_7_2_r;
wire signed [`CalcTempBus]          temp_m3_7_2_i;
wire signed [`CalcTempBus]          temp_m3_7_3_r;
wire signed [`CalcTempBus]          temp_m3_7_3_i;
wire signed [`CalcTempBus]          temp_m3_7_4_r;
wire signed [`CalcTempBus]          temp_m3_7_4_i;
wire signed [`CalcTempBus]          temp_m3_7_5_r;
wire signed [`CalcTempBus]          temp_m3_7_5_i;
wire signed [`CalcTempBus]          temp_m3_7_6_r;
wire signed [`CalcTempBus]          temp_m3_7_6_i;
wire signed [`CalcTempBus]          temp_m3_7_7_r;
wire signed [`CalcTempBus]          temp_m3_7_7_i;
wire signed [`CalcTempBus]          temp_m3_7_8_r;
wire signed [`CalcTempBus]          temp_m3_7_8_i;
wire signed [`CalcTempBus]          temp_m3_7_9_r;
wire signed [`CalcTempBus]          temp_m3_7_9_i;
wire signed [`CalcTempBus]          temp_m3_7_10_r;
wire signed [`CalcTempBus]          temp_m3_7_10_i;
wire signed [`CalcTempBus]          temp_m3_7_11_r;
wire signed [`CalcTempBus]          temp_m3_7_11_i;
wire signed [`CalcTempBus]          temp_m3_7_12_r;
wire signed [`CalcTempBus]          temp_m3_7_12_i;
wire signed [`CalcTempBus]          temp_m3_7_13_r;
wire signed [`CalcTempBus]          temp_m3_7_13_i;
wire signed [`CalcTempBus]          temp_m3_7_14_r;
wire signed [`CalcTempBus]          temp_m3_7_14_i;
wire signed [`CalcTempBus]          temp_m3_7_15_r;
wire signed [`CalcTempBus]          temp_m3_7_15_i;
wire signed [`CalcTempBus]          temp_m3_7_16_r;
wire signed [`CalcTempBus]          temp_m3_7_16_i;
wire signed [`CalcTempBus]          temp_m3_8_1_r;
wire signed [`CalcTempBus]          temp_m3_8_1_i;
wire signed [`CalcTempBus]          temp_m3_8_2_r;
wire signed [`CalcTempBus]          temp_m3_8_2_i;
wire signed [`CalcTempBus]          temp_m3_8_3_r;
wire signed [`CalcTempBus]          temp_m3_8_3_i;
wire signed [`CalcTempBus]          temp_m3_8_4_r;
wire signed [`CalcTempBus]          temp_m3_8_4_i;
wire signed [`CalcTempBus]          temp_m3_8_5_r;
wire signed [`CalcTempBus]          temp_m3_8_5_i;
wire signed [`CalcTempBus]          temp_m3_8_6_r;
wire signed [`CalcTempBus]          temp_m3_8_6_i;
wire signed [`CalcTempBus]          temp_m3_8_7_r;
wire signed [`CalcTempBus]          temp_m3_8_7_i;
wire signed [`CalcTempBus]          temp_m3_8_8_r;
wire signed [`CalcTempBus]          temp_m3_8_8_i;
wire signed [`CalcTempBus]          temp_m3_8_9_r;
wire signed [`CalcTempBus]          temp_m3_8_9_i;
wire signed [`CalcTempBus]          temp_m3_8_10_r;
wire signed [`CalcTempBus]          temp_m3_8_10_i;
wire signed [`CalcTempBus]          temp_m3_8_11_r;
wire signed [`CalcTempBus]          temp_m3_8_11_i;
wire signed [`CalcTempBus]          temp_m3_8_12_r;
wire signed [`CalcTempBus]          temp_m3_8_12_i;
wire signed [`CalcTempBus]          temp_m3_8_13_r;
wire signed [`CalcTempBus]          temp_m3_8_13_i;
wire signed [`CalcTempBus]          temp_m3_8_14_r;
wire signed [`CalcTempBus]          temp_m3_8_14_i;
wire signed [`CalcTempBus]          temp_m3_8_15_r;
wire signed [`CalcTempBus]          temp_m3_8_15_i;
wire signed [`CalcTempBus]          temp_m3_8_16_r;
wire signed [`CalcTempBus]          temp_m3_8_16_i;
wire signed [`CalcTempBus]          temp_m3_9_1_r;
wire signed [`CalcTempBus]          temp_m3_9_1_i;
wire signed [`CalcTempBus]          temp_m3_9_2_r;
wire signed [`CalcTempBus]          temp_m3_9_2_i;
wire signed [`CalcTempBus]          temp_m3_9_3_r;
wire signed [`CalcTempBus]          temp_m3_9_3_i;
wire signed [`CalcTempBus]          temp_m3_9_4_r;
wire signed [`CalcTempBus]          temp_m3_9_4_i;
wire signed [`CalcTempBus]          temp_m3_9_5_r;
wire signed [`CalcTempBus]          temp_m3_9_5_i;
wire signed [`CalcTempBus]          temp_m3_9_6_r;
wire signed [`CalcTempBus]          temp_m3_9_6_i;
wire signed [`CalcTempBus]          temp_m3_9_7_r;
wire signed [`CalcTempBus]          temp_m3_9_7_i;
wire signed [`CalcTempBus]          temp_m3_9_8_r;
wire signed [`CalcTempBus]          temp_m3_9_8_i;
wire signed [`CalcTempBus]          temp_m3_9_9_r;
wire signed [`CalcTempBus]          temp_m3_9_9_i;
wire signed [`CalcTempBus]          temp_m3_9_10_r;
wire signed [`CalcTempBus]          temp_m3_9_10_i;
wire signed [`CalcTempBus]          temp_m3_9_11_r;
wire signed [`CalcTempBus]          temp_m3_9_11_i;
wire signed [`CalcTempBus]          temp_m3_9_12_r;
wire signed [`CalcTempBus]          temp_m3_9_12_i;
wire signed [`CalcTempBus]          temp_m3_9_13_r;
wire signed [`CalcTempBus]          temp_m3_9_13_i;
wire signed [`CalcTempBus]          temp_m3_9_14_r;
wire signed [`CalcTempBus]          temp_m3_9_14_i;
wire signed [`CalcTempBus]          temp_m3_9_15_r;
wire signed [`CalcTempBus]          temp_m3_9_15_i;
wire signed [`CalcTempBus]          temp_m3_9_16_r;
wire signed [`CalcTempBus]          temp_m3_9_16_i;
wire signed [`CalcTempBus]          temp_m3_10_1_r;
wire signed [`CalcTempBus]          temp_m3_10_1_i;
wire signed [`CalcTempBus]          temp_m3_10_2_r;
wire signed [`CalcTempBus]          temp_m3_10_2_i;
wire signed [`CalcTempBus]          temp_m3_10_3_r;
wire signed [`CalcTempBus]          temp_m3_10_3_i;
wire signed [`CalcTempBus]          temp_m3_10_4_r;
wire signed [`CalcTempBus]          temp_m3_10_4_i;
wire signed [`CalcTempBus]          temp_m3_10_5_r;
wire signed [`CalcTempBus]          temp_m3_10_5_i;
wire signed [`CalcTempBus]          temp_m3_10_6_r;
wire signed [`CalcTempBus]          temp_m3_10_6_i;
wire signed [`CalcTempBus]          temp_m3_10_7_r;
wire signed [`CalcTempBus]          temp_m3_10_7_i;
wire signed [`CalcTempBus]          temp_m3_10_8_r;
wire signed [`CalcTempBus]          temp_m3_10_8_i;
wire signed [`CalcTempBus]          temp_m3_10_9_r;
wire signed [`CalcTempBus]          temp_m3_10_9_i;
wire signed [`CalcTempBus]          temp_m3_10_10_r;
wire signed [`CalcTempBus]          temp_m3_10_10_i;
wire signed [`CalcTempBus]          temp_m3_10_11_r;
wire signed [`CalcTempBus]          temp_m3_10_11_i;
wire signed [`CalcTempBus]          temp_m3_10_12_r;
wire signed [`CalcTempBus]          temp_m3_10_12_i;
wire signed [`CalcTempBus]          temp_m3_10_13_r;
wire signed [`CalcTempBus]          temp_m3_10_13_i;
wire signed [`CalcTempBus]          temp_m3_10_14_r;
wire signed [`CalcTempBus]          temp_m3_10_14_i;
wire signed [`CalcTempBus]          temp_m3_10_15_r;
wire signed [`CalcTempBus]          temp_m3_10_15_i;
wire signed [`CalcTempBus]          temp_m3_10_16_r;
wire signed [`CalcTempBus]          temp_m3_10_16_i;
wire signed [`CalcTempBus]          temp_m3_11_1_r;
wire signed [`CalcTempBus]          temp_m3_11_1_i;
wire signed [`CalcTempBus]          temp_m3_11_2_r;
wire signed [`CalcTempBus]          temp_m3_11_2_i;
wire signed [`CalcTempBus]          temp_m3_11_3_r;
wire signed [`CalcTempBus]          temp_m3_11_3_i;
wire signed [`CalcTempBus]          temp_m3_11_4_r;
wire signed [`CalcTempBus]          temp_m3_11_4_i;
wire signed [`CalcTempBus]          temp_m3_11_5_r;
wire signed [`CalcTempBus]          temp_m3_11_5_i;
wire signed [`CalcTempBus]          temp_m3_11_6_r;
wire signed [`CalcTempBus]          temp_m3_11_6_i;
wire signed [`CalcTempBus]          temp_m3_11_7_r;
wire signed [`CalcTempBus]          temp_m3_11_7_i;
wire signed [`CalcTempBus]          temp_m3_11_8_r;
wire signed [`CalcTempBus]          temp_m3_11_8_i;
wire signed [`CalcTempBus]          temp_m3_11_9_r;
wire signed [`CalcTempBus]          temp_m3_11_9_i;
wire signed [`CalcTempBus]          temp_m3_11_10_r;
wire signed [`CalcTempBus]          temp_m3_11_10_i;
wire signed [`CalcTempBus]          temp_m3_11_11_r;
wire signed [`CalcTempBus]          temp_m3_11_11_i;
wire signed [`CalcTempBus]          temp_m3_11_12_r;
wire signed [`CalcTempBus]          temp_m3_11_12_i;
wire signed [`CalcTempBus]          temp_m3_11_13_r;
wire signed [`CalcTempBus]          temp_m3_11_13_i;
wire signed [`CalcTempBus]          temp_m3_11_14_r;
wire signed [`CalcTempBus]          temp_m3_11_14_i;
wire signed [`CalcTempBus]          temp_m3_11_15_r;
wire signed [`CalcTempBus]          temp_m3_11_15_i;
wire signed [`CalcTempBus]          temp_m3_11_16_r;
wire signed [`CalcTempBus]          temp_m3_11_16_i;
wire signed [`CalcTempBus]          temp_m3_12_1_r;
wire signed [`CalcTempBus]          temp_m3_12_1_i;
wire signed [`CalcTempBus]          temp_m3_12_2_r;
wire signed [`CalcTempBus]          temp_m3_12_2_i;
wire signed [`CalcTempBus]          temp_m3_12_3_r;
wire signed [`CalcTempBus]          temp_m3_12_3_i;
wire signed [`CalcTempBus]          temp_m3_12_4_r;
wire signed [`CalcTempBus]          temp_m3_12_4_i;
wire signed [`CalcTempBus]          temp_m3_12_5_r;
wire signed [`CalcTempBus]          temp_m3_12_5_i;
wire signed [`CalcTempBus]          temp_m3_12_6_r;
wire signed [`CalcTempBus]          temp_m3_12_6_i;
wire signed [`CalcTempBus]          temp_m3_12_7_r;
wire signed [`CalcTempBus]          temp_m3_12_7_i;
wire signed [`CalcTempBus]          temp_m3_12_8_r;
wire signed [`CalcTempBus]          temp_m3_12_8_i;
wire signed [`CalcTempBus]          temp_m3_12_9_r;
wire signed [`CalcTempBus]          temp_m3_12_9_i;
wire signed [`CalcTempBus]          temp_m3_12_10_r;
wire signed [`CalcTempBus]          temp_m3_12_10_i;
wire signed [`CalcTempBus]          temp_m3_12_11_r;
wire signed [`CalcTempBus]          temp_m3_12_11_i;
wire signed [`CalcTempBus]          temp_m3_12_12_r;
wire signed [`CalcTempBus]          temp_m3_12_12_i;
wire signed [`CalcTempBus]          temp_m3_12_13_r;
wire signed [`CalcTempBus]          temp_m3_12_13_i;
wire signed [`CalcTempBus]          temp_m3_12_14_r;
wire signed [`CalcTempBus]          temp_m3_12_14_i;
wire signed [`CalcTempBus]          temp_m3_12_15_r;
wire signed [`CalcTempBus]          temp_m3_12_15_i;
wire signed [`CalcTempBus]          temp_m3_12_16_r;
wire signed [`CalcTempBus]          temp_m3_12_16_i;
wire signed [`CalcTempBus]          temp_m3_13_1_r;
wire signed [`CalcTempBus]          temp_m3_13_1_i;
wire signed [`CalcTempBus]          temp_m3_13_2_r;
wire signed [`CalcTempBus]          temp_m3_13_2_i;
wire signed [`CalcTempBus]          temp_m3_13_3_r;
wire signed [`CalcTempBus]          temp_m3_13_3_i;
wire signed [`CalcTempBus]          temp_m3_13_4_r;
wire signed [`CalcTempBus]          temp_m3_13_4_i;
wire signed [`CalcTempBus]          temp_m3_13_5_r;
wire signed [`CalcTempBus]          temp_m3_13_5_i;
wire signed [`CalcTempBus]          temp_m3_13_6_r;
wire signed [`CalcTempBus]          temp_m3_13_6_i;
wire signed [`CalcTempBus]          temp_m3_13_7_r;
wire signed [`CalcTempBus]          temp_m3_13_7_i;
wire signed [`CalcTempBus]          temp_m3_13_8_r;
wire signed [`CalcTempBus]          temp_m3_13_8_i;
wire signed [`CalcTempBus]          temp_m3_13_9_r;
wire signed [`CalcTempBus]          temp_m3_13_9_i;
wire signed [`CalcTempBus]          temp_m3_13_10_r;
wire signed [`CalcTempBus]          temp_m3_13_10_i;
wire signed [`CalcTempBus]          temp_m3_13_11_r;
wire signed [`CalcTempBus]          temp_m3_13_11_i;
wire signed [`CalcTempBus]          temp_m3_13_12_r;
wire signed [`CalcTempBus]          temp_m3_13_12_i;
wire signed [`CalcTempBus]          temp_m3_13_13_r;
wire signed [`CalcTempBus]          temp_m3_13_13_i;
wire signed [`CalcTempBus]          temp_m3_13_14_r;
wire signed [`CalcTempBus]          temp_m3_13_14_i;
wire signed [`CalcTempBus]          temp_m3_13_15_r;
wire signed [`CalcTempBus]          temp_m3_13_15_i;
wire signed [`CalcTempBus]          temp_m3_13_16_r;
wire signed [`CalcTempBus]          temp_m3_13_16_i;
wire signed [`CalcTempBus]          temp_m3_14_1_r;
wire signed [`CalcTempBus]          temp_m3_14_1_i;
wire signed [`CalcTempBus]          temp_m3_14_2_r;
wire signed [`CalcTempBus]          temp_m3_14_2_i;
wire signed [`CalcTempBus]          temp_m3_14_3_r;
wire signed [`CalcTempBus]          temp_m3_14_3_i;
wire signed [`CalcTempBus]          temp_m3_14_4_r;
wire signed [`CalcTempBus]          temp_m3_14_4_i;
wire signed [`CalcTempBus]          temp_m3_14_5_r;
wire signed [`CalcTempBus]          temp_m3_14_5_i;
wire signed [`CalcTempBus]          temp_m3_14_6_r;
wire signed [`CalcTempBus]          temp_m3_14_6_i;
wire signed [`CalcTempBus]          temp_m3_14_7_r;
wire signed [`CalcTempBus]          temp_m3_14_7_i;
wire signed [`CalcTempBus]          temp_m3_14_8_r;
wire signed [`CalcTempBus]          temp_m3_14_8_i;
wire signed [`CalcTempBus]          temp_m3_14_9_r;
wire signed [`CalcTempBus]          temp_m3_14_9_i;
wire signed [`CalcTempBus]          temp_m3_14_10_r;
wire signed [`CalcTempBus]          temp_m3_14_10_i;
wire signed [`CalcTempBus]          temp_m3_14_11_r;
wire signed [`CalcTempBus]          temp_m3_14_11_i;
wire signed [`CalcTempBus]          temp_m3_14_12_r;
wire signed [`CalcTempBus]          temp_m3_14_12_i;
wire signed [`CalcTempBus]          temp_m3_14_13_r;
wire signed [`CalcTempBus]          temp_m3_14_13_i;
wire signed [`CalcTempBus]          temp_m3_14_14_r;
wire signed [`CalcTempBus]          temp_m3_14_14_i;
wire signed [`CalcTempBus]          temp_m3_14_15_r;
wire signed [`CalcTempBus]          temp_m3_14_15_i;
wire signed [`CalcTempBus]          temp_m3_14_16_r;
wire signed [`CalcTempBus]          temp_m3_14_16_i;
wire signed [`CalcTempBus]          temp_m3_15_1_r;
wire signed [`CalcTempBus]          temp_m3_15_1_i;
wire signed [`CalcTempBus]          temp_m3_15_2_r;
wire signed [`CalcTempBus]          temp_m3_15_2_i;
wire signed [`CalcTempBus]          temp_m3_15_3_r;
wire signed [`CalcTempBus]          temp_m3_15_3_i;
wire signed [`CalcTempBus]          temp_m3_15_4_r;
wire signed [`CalcTempBus]          temp_m3_15_4_i;
wire signed [`CalcTempBus]          temp_m3_15_5_r;
wire signed [`CalcTempBus]          temp_m3_15_5_i;
wire signed [`CalcTempBus]          temp_m3_15_6_r;
wire signed [`CalcTempBus]          temp_m3_15_6_i;
wire signed [`CalcTempBus]          temp_m3_15_7_r;
wire signed [`CalcTempBus]          temp_m3_15_7_i;
wire signed [`CalcTempBus]          temp_m3_15_8_r;
wire signed [`CalcTempBus]          temp_m3_15_8_i;
wire signed [`CalcTempBus]          temp_m3_15_9_r;
wire signed [`CalcTempBus]          temp_m3_15_9_i;
wire signed [`CalcTempBus]          temp_m3_15_10_r;
wire signed [`CalcTempBus]          temp_m3_15_10_i;
wire signed [`CalcTempBus]          temp_m3_15_11_r;
wire signed [`CalcTempBus]          temp_m3_15_11_i;
wire signed [`CalcTempBus]          temp_m3_15_12_r;
wire signed [`CalcTempBus]          temp_m3_15_12_i;
wire signed [`CalcTempBus]          temp_m3_15_13_r;
wire signed [`CalcTempBus]          temp_m3_15_13_i;
wire signed [`CalcTempBus]          temp_m3_15_14_r;
wire signed [`CalcTempBus]          temp_m3_15_14_i;
wire signed [`CalcTempBus]          temp_m3_15_15_r;
wire signed [`CalcTempBus]          temp_m3_15_15_i;
wire signed [`CalcTempBus]          temp_m3_15_16_r;
wire signed [`CalcTempBus]          temp_m3_15_16_i;
wire signed [`CalcTempBus]          temp_m3_16_1_r;
wire signed [`CalcTempBus]          temp_m3_16_1_i;
wire signed [`CalcTempBus]          temp_m3_16_2_r;
wire signed [`CalcTempBus]          temp_m3_16_2_i;
wire signed [`CalcTempBus]          temp_m3_16_3_r;
wire signed [`CalcTempBus]          temp_m3_16_3_i;
wire signed [`CalcTempBus]          temp_m3_16_4_r;
wire signed [`CalcTempBus]          temp_m3_16_4_i;
wire signed [`CalcTempBus]          temp_m3_16_5_r;
wire signed [`CalcTempBus]          temp_m3_16_5_i;
wire signed [`CalcTempBus]          temp_m3_16_6_r;
wire signed [`CalcTempBus]          temp_m3_16_6_i;
wire signed [`CalcTempBus]          temp_m3_16_7_r;
wire signed [`CalcTempBus]          temp_m3_16_7_i;
wire signed [`CalcTempBus]          temp_m3_16_8_r;
wire signed [`CalcTempBus]          temp_m3_16_8_i;
wire signed [`CalcTempBus]          temp_m3_16_9_r;
wire signed [`CalcTempBus]          temp_m3_16_9_i;
wire signed [`CalcTempBus]          temp_m3_16_10_r;
wire signed [`CalcTempBus]          temp_m3_16_10_i;
wire signed [`CalcTempBus]          temp_m3_16_11_r;
wire signed [`CalcTempBus]          temp_m3_16_11_i;
wire signed [`CalcTempBus]          temp_m3_16_12_r;
wire signed [`CalcTempBus]          temp_m3_16_12_i;
wire signed [`CalcTempBus]          temp_m3_16_13_r;
wire signed [`CalcTempBus]          temp_m3_16_13_i;
wire signed [`CalcTempBus]          temp_m3_16_14_r;
wire signed [`CalcTempBus]          temp_m3_16_14_i;
wire signed [`CalcTempBus]          temp_m3_16_15_r;
wire signed [`CalcTempBus]          temp_m3_16_15_i;
wire signed [`CalcTempBus]          temp_m3_16_16_r;
wire signed [`CalcTempBus]          temp_m3_16_16_i;
wire signed [`CalcTempBus]          temp_m4_1_1_r;
wire signed [`CalcTempBus]          temp_m4_1_1_i;
wire signed [`CalcTempBus]          temp_m4_1_2_r;
wire signed [`CalcTempBus]          temp_m4_1_2_i;
wire signed [`CalcTempBus]          temp_m4_1_3_r;
wire signed [`CalcTempBus]          temp_m4_1_3_i;
wire signed [`CalcTempBus]          temp_m4_1_4_r;
wire signed [`CalcTempBus]          temp_m4_1_4_i;
wire signed [`CalcTempBus]          temp_m4_1_5_r;
wire signed [`CalcTempBus]          temp_m4_1_5_i;
wire signed [`CalcTempBus]          temp_m4_1_6_r;
wire signed [`CalcTempBus]          temp_m4_1_6_i;
wire signed [`CalcTempBus]          temp_m4_1_7_r;
wire signed [`CalcTempBus]          temp_m4_1_7_i;
wire signed [`CalcTempBus]          temp_m4_1_8_r;
wire signed [`CalcTempBus]          temp_m4_1_8_i;
wire signed [`CalcTempBus]          temp_m4_1_9_r;
wire signed [`CalcTempBus]          temp_m4_1_9_i;
wire signed [`CalcTempBus]          temp_m4_1_10_r;
wire signed [`CalcTempBus]          temp_m4_1_10_i;
wire signed [`CalcTempBus]          temp_m4_1_11_r;
wire signed [`CalcTempBus]          temp_m4_1_11_i;
wire signed [`CalcTempBus]          temp_m4_1_12_r;
wire signed [`CalcTempBus]          temp_m4_1_12_i;
wire signed [`CalcTempBus]          temp_m4_1_13_r;
wire signed [`CalcTempBus]          temp_m4_1_13_i;
wire signed [`CalcTempBus]          temp_m4_1_14_r;
wire signed [`CalcTempBus]          temp_m4_1_14_i;
wire signed [`CalcTempBus]          temp_m4_1_15_r;
wire signed [`CalcTempBus]          temp_m4_1_15_i;
wire signed [`CalcTempBus]          temp_m4_1_16_r;
wire signed [`CalcTempBus]          temp_m4_1_16_i;
wire signed [`CalcTempBus]          temp_m4_2_1_r;
wire signed [`CalcTempBus]          temp_m4_2_1_i;
wire signed [`CalcTempBus]          temp_m4_2_2_r;
wire signed [`CalcTempBus]          temp_m4_2_2_i;
wire signed [`CalcTempBus]          temp_m4_2_3_r;
wire signed [`CalcTempBus]          temp_m4_2_3_i;
wire signed [`CalcTempBus]          temp_m4_2_4_r;
wire signed [`CalcTempBus]          temp_m4_2_4_i;
wire signed [`CalcTempBus]          temp_m4_2_5_r;
wire signed [`CalcTempBus]          temp_m4_2_5_i;
wire signed [`CalcTempBus]          temp_m4_2_6_r;
wire signed [`CalcTempBus]          temp_m4_2_6_i;
wire signed [`CalcTempBus]          temp_m4_2_7_r;
wire signed [`CalcTempBus]          temp_m4_2_7_i;
wire signed [`CalcTempBus]          temp_m4_2_8_r;
wire signed [`CalcTempBus]          temp_m4_2_8_i;
wire signed [`CalcTempBus]          temp_m4_2_9_r;
wire signed [`CalcTempBus]          temp_m4_2_9_i;
wire signed [`CalcTempBus]          temp_m4_2_10_r;
wire signed [`CalcTempBus]          temp_m4_2_10_i;
wire signed [`CalcTempBus]          temp_m4_2_11_r;
wire signed [`CalcTempBus]          temp_m4_2_11_i;
wire signed [`CalcTempBus]          temp_m4_2_12_r;
wire signed [`CalcTempBus]          temp_m4_2_12_i;
wire signed [`CalcTempBus]          temp_m4_2_13_r;
wire signed [`CalcTempBus]          temp_m4_2_13_i;
wire signed [`CalcTempBus]          temp_m4_2_14_r;
wire signed [`CalcTempBus]          temp_m4_2_14_i;
wire signed [`CalcTempBus]          temp_m4_2_15_r;
wire signed [`CalcTempBus]          temp_m4_2_15_i;
wire signed [`CalcTempBus]          temp_m4_2_16_r;
wire signed [`CalcTempBus]          temp_m4_2_16_i;
wire signed [`CalcTempBus]          temp_m4_3_1_r;
wire signed [`CalcTempBus]          temp_m4_3_1_i;
wire signed [`CalcTempBus]          temp_m4_3_2_r;
wire signed [`CalcTempBus]          temp_m4_3_2_i;
wire signed [`CalcTempBus]          temp_m4_3_3_r;
wire signed [`CalcTempBus]          temp_m4_3_3_i;
wire signed [`CalcTempBus]          temp_m4_3_4_r;
wire signed [`CalcTempBus]          temp_m4_3_4_i;
wire signed [`CalcTempBus]          temp_m4_3_5_r;
wire signed [`CalcTempBus]          temp_m4_3_5_i;
wire signed [`CalcTempBus]          temp_m4_3_6_r;
wire signed [`CalcTempBus]          temp_m4_3_6_i;
wire signed [`CalcTempBus]          temp_m4_3_7_r;
wire signed [`CalcTempBus]          temp_m4_3_7_i;
wire signed [`CalcTempBus]          temp_m4_3_8_r;
wire signed [`CalcTempBus]          temp_m4_3_8_i;
wire signed [`CalcTempBus]          temp_m4_3_9_r;
wire signed [`CalcTempBus]          temp_m4_3_9_i;
wire signed [`CalcTempBus]          temp_m4_3_10_r;
wire signed [`CalcTempBus]          temp_m4_3_10_i;
wire signed [`CalcTempBus]          temp_m4_3_11_r;
wire signed [`CalcTempBus]          temp_m4_3_11_i;
wire signed [`CalcTempBus]          temp_m4_3_12_r;
wire signed [`CalcTempBus]          temp_m4_3_12_i;
wire signed [`CalcTempBus]          temp_m4_3_13_r;
wire signed [`CalcTempBus]          temp_m4_3_13_i;
wire signed [`CalcTempBus]          temp_m4_3_14_r;
wire signed [`CalcTempBus]          temp_m4_3_14_i;
wire signed [`CalcTempBus]          temp_m4_3_15_r;
wire signed [`CalcTempBus]          temp_m4_3_15_i;
wire signed [`CalcTempBus]          temp_m4_3_16_r;
wire signed [`CalcTempBus]          temp_m4_3_16_i;
wire signed [`CalcTempBus]          temp_m4_4_1_r;
wire signed [`CalcTempBus]          temp_m4_4_1_i;
wire signed [`CalcTempBus]          temp_m4_4_2_r;
wire signed [`CalcTempBus]          temp_m4_4_2_i;
wire signed [`CalcTempBus]          temp_m4_4_3_r;
wire signed [`CalcTempBus]          temp_m4_4_3_i;
wire signed [`CalcTempBus]          temp_m4_4_4_r;
wire signed [`CalcTempBus]          temp_m4_4_4_i;
wire signed [`CalcTempBus]          temp_m4_4_5_r;
wire signed [`CalcTempBus]          temp_m4_4_5_i;
wire signed [`CalcTempBus]          temp_m4_4_6_r;
wire signed [`CalcTempBus]          temp_m4_4_6_i;
wire signed [`CalcTempBus]          temp_m4_4_7_r;
wire signed [`CalcTempBus]          temp_m4_4_7_i;
wire signed [`CalcTempBus]          temp_m4_4_8_r;
wire signed [`CalcTempBus]          temp_m4_4_8_i;
wire signed [`CalcTempBus]          temp_m4_4_9_r;
wire signed [`CalcTempBus]          temp_m4_4_9_i;
wire signed [`CalcTempBus]          temp_m4_4_10_r;
wire signed [`CalcTempBus]          temp_m4_4_10_i;
wire signed [`CalcTempBus]          temp_m4_4_11_r;
wire signed [`CalcTempBus]          temp_m4_4_11_i;
wire signed [`CalcTempBus]          temp_m4_4_12_r;
wire signed [`CalcTempBus]          temp_m4_4_12_i;
wire signed [`CalcTempBus]          temp_m4_4_13_r;
wire signed [`CalcTempBus]          temp_m4_4_13_i;
wire signed [`CalcTempBus]          temp_m4_4_14_r;
wire signed [`CalcTempBus]          temp_m4_4_14_i;
wire signed [`CalcTempBus]          temp_m4_4_15_r;
wire signed [`CalcTempBus]          temp_m4_4_15_i;
wire signed [`CalcTempBus]          temp_m4_4_16_r;
wire signed [`CalcTempBus]          temp_m4_4_16_i;
wire signed [`CalcTempBus]          temp_m4_5_1_r;
wire signed [`CalcTempBus]          temp_m4_5_1_i;
wire signed [`CalcTempBus]          temp_m4_5_2_r;
wire signed [`CalcTempBus]          temp_m4_5_2_i;
wire signed [`CalcTempBus]          temp_m4_5_3_r;
wire signed [`CalcTempBus]          temp_m4_5_3_i;
wire signed [`CalcTempBus]          temp_m4_5_4_r;
wire signed [`CalcTempBus]          temp_m4_5_4_i;
wire signed [`CalcTempBus]          temp_m4_5_5_r;
wire signed [`CalcTempBus]          temp_m4_5_5_i;
wire signed [`CalcTempBus]          temp_m4_5_6_r;
wire signed [`CalcTempBus]          temp_m4_5_6_i;
wire signed [`CalcTempBus]          temp_m4_5_7_r;
wire signed [`CalcTempBus]          temp_m4_5_7_i;
wire signed [`CalcTempBus]          temp_m4_5_8_r;
wire signed [`CalcTempBus]          temp_m4_5_8_i;
wire signed [`CalcTempBus]          temp_m4_5_9_r;
wire signed [`CalcTempBus]          temp_m4_5_9_i;
wire signed [`CalcTempBus]          temp_m4_5_10_r;
wire signed [`CalcTempBus]          temp_m4_5_10_i;
wire signed [`CalcTempBus]          temp_m4_5_11_r;
wire signed [`CalcTempBus]          temp_m4_5_11_i;
wire signed [`CalcTempBus]          temp_m4_5_12_r;
wire signed [`CalcTempBus]          temp_m4_5_12_i;
wire signed [`CalcTempBus]          temp_m4_5_13_r;
wire signed [`CalcTempBus]          temp_m4_5_13_i;
wire signed [`CalcTempBus]          temp_m4_5_14_r;
wire signed [`CalcTempBus]          temp_m4_5_14_i;
wire signed [`CalcTempBus]          temp_m4_5_15_r;
wire signed [`CalcTempBus]          temp_m4_5_15_i;
wire signed [`CalcTempBus]          temp_m4_5_16_r;
wire signed [`CalcTempBus]          temp_m4_5_16_i;
wire signed [`CalcTempBus]          temp_m4_6_1_r;
wire signed [`CalcTempBus]          temp_m4_6_1_i;
wire signed [`CalcTempBus]          temp_m4_6_2_r;
wire signed [`CalcTempBus]          temp_m4_6_2_i;
wire signed [`CalcTempBus]          temp_m4_6_3_r;
wire signed [`CalcTempBus]          temp_m4_6_3_i;
wire signed [`CalcTempBus]          temp_m4_6_4_r;
wire signed [`CalcTempBus]          temp_m4_6_4_i;
wire signed [`CalcTempBus]          temp_m4_6_5_r;
wire signed [`CalcTempBus]          temp_m4_6_5_i;
wire signed [`CalcTempBus]          temp_m4_6_6_r;
wire signed [`CalcTempBus]          temp_m4_6_6_i;
wire signed [`CalcTempBus]          temp_m4_6_7_r;
wire signed [`CalcTempBus]          temp_m4_6_7_i;
wire signed [`CalcTempBus]          temp_m4_6_8_r;
wire signed [`CalcTempBus]          temp_m4_6_8_i;
wire signed [`CalcTempBus]          temp_m4_6_9_r;
wire signed [`CalcTempBus]          temp_m4_6_9_i;
wire signed [`CalcTempBus]          temp_m4_6_10_r;
wire signed [`CalcTempBus]          temp_m4_6_10_i;
wire signed [`CalcTempBus]          temp_m4_6_11_r;
wire signed [`CalcTempBus]          temp_m4_6_11_i;
wire signed [`CalcTempBus]          temp_m4_6_12_r;
wire signed [`CalcTempBus]          temp_m4_6_12_i;
wire signed [`CalcTempBus]          temp_m4_6_13_r;
wire signed [`CalcTempBus]          temp_m4_6_13_i;
wire signed [`CalcTempBus]          temp_m4_6_14_r;
wire signed [`CalcTempBus]          temp_m4_6_14_i;
wire signed [`CalcTempBus]          temp_m4_6_15_r;
wire signed [`CalcTempBus]          temp_m4_6_15_i;
wire signed [`CalcTempBus]          temp_m4_6_16_r;
wire signed [`CalcTempBus]          temp_m4_6_16_i;
wire signed [`CalcTempBus]          temp_m4_7_1_r;
wire signed [`CalcTempBus]          temp_m4_7_1_i;
wire signed [`CalcTempBus]          temp_m4_7_2_r;
wire signed [`CalcTempBus]          temp_m4_7_2_i;
wire signed [`CalcTempBus]          temp_m4_7_3_r;
wire signed [`CalcTempBus]          temp_m4_7_3_i;
wire signed [`CalcTempBus]          temp_m4_7_4_r;
wire signed [`CalcTempBus]          temp_m4_7_4_i;
wire signed [`CalcTempBus]          temp_m4_7_5_r;
wire signed [`CalcTempBus]          temp_m4_7_5_i;
wire signed [`CalcTempBus]          temp_m4_7_6_r;
wire signed [`CalcTempBus]          temp_m4_7_6_i;
wire signed [`CalcTempBus]          temp_m4_7_7_r;
wire signed [`CalcTempBus]          temp_m4_7_7_i;
wire signed [`CalcTempBus]          temp_m4_7_8_r;
wire signed [`CalcTempBus]          temp_m4_7_8_i;
wire signed [`CalcTempBus]          temp_m4_7_9_r;
wire signed [`CalcTempBus]          temp_m4_7_9_i;
wire signed [`CalcTempBus]          temp_m4_7_10_r;
wire signed [`CalcTempBus]          temp_m4_7_10_i;
wire signed [`CalcTempBus]          temp_m4_7_11_r;
wire signed [`CalcTempBus]          temp_m4_7_11_i;
wire signed [`CalcTempBus]          temp_m4_7_12_r;
wire signed [`CalcTempBus]          temp_m4_7_12_i;
wire signed [`CalcTempBus]          temp_m4_7_13_r;
wire signed [`CalcTempBus]          temp_m4_7_13_i;
wire signed [`CalcTempBus]          temp_m4_7_14_r;
wire signed [`CalcTempBus]          temp_m4_7_14_i;
wire signed [`CalcTempBus]          temp_m4_7_15_r;
wire signed [`CalcTempBus]          temp_m4_7_15_i;
wire signed [`CalcTempBus]          temp_m4_7_16_r;
wire signed [`CalcTempBus]          temp_m4_7_16_i;
wire signed [`CalcTempBus]          temp_m4_8_1_r;
wire signed [`CalcTempBus]          temp_m4_8_1_i;
wire signed [`CalcTempBus]          temp_m4_8_2_r;
wire signed [`CalcTempBus]          temp_m4_8_2_i;
wire signed [`CalcTempBus]          temp_m4_8_3_r;
wire signed [`CalcTempBus]          temp_m4_8_3_i;
wire signed [`CalcTempBus]          temp_m4_8_4_r;
wire signed [`CalcTempBus]          temp_m4_8_4_i;
wire signed [`CalcTempBus]          temp_m4_8_5_r;
wire signed [`CalcTempBus]          temp_m4_8_5_i;
wire signed [`CalcTempBus]          temp_m4_8_6_r;
wire signed [`CalcTempBus]          temp_m4_8_6_i;
wire signed [`CalcTempBus]          temp_m4_8_7_r;
wire signed [`CalcTempBus]          temp_m4_8_7_i;
wire signed [`CalcTempBus]          temp_m4_8_8_r;
wire signed [`CalcTempBus]          temp_m4_8_8_i;
wire signed [`CalcTempBus]          temp_m4_8_9_r;
wire signed [`CalcTempBus]          temp_m4_8_9_i;
wire signed [`CalcTempBus]          temp_m4_8_10_r;
wire signed [`CalcTempBus]          temp_m4_8_10_i;
wire signed [`CalcTempBus]          temp_m4_8_11_r;
wire signed [`CalcTempBus]          temp_m4_8_11_i;
wire signed [`CalcTempBus]          temp_m4_8_12_r;
wire signed [`CalcTempBus]          temp_m4_8_12_i;
wire signed [`CalcTempBus]          temp_m4_8_13_r;
wire signed [`CalcTempBus]          temp_m4_8_13_i;
wire signed [`CalcTempBus]          temp_m4_8_14_r;
wire signed [`CalcTempBus]          temp_m4_8_14_i;
wire signed [`CalcTempBus]          temp_m4_8_15_r;
wire signed [`CalcTempBus]          temp_m4_8_15_i;
wire signed [`CalcTempBus]          temp_m4_8_16_r;
wire signed [`CalcTempBus]          temp_m4_8_16_i;
wire signed [`CalcTempBus]          temp_m4_9_1_r;
wire signed [`CalcTempBus]          temp_m4_9_1_i;
wire signed [`CalcTempBus]          temp_m4_9_2_r;
wire signed [`CalcTempBus]          temp_m4_9_2_i;
wire signed [`CalcTempBus]          temp_m4_9_3_r;
wire signed [`CalcTempBus]          temp_m4_9_3_i;
wire signed [`CalcTempBus]          temp_m4_9_4_r;
wire signed [`CalcTempBus]          temp_m4_9_4_i;
wire signed [`CalcTempBus]          temp_m4_9_5_r;
wire signed [`CalcTempBus]          temp_m4_9_5_i;
wire signed [`CalcTempBus]          temp_m4_9_6_r;
wire signed [`CalcTempBus]          temp_m4_9_6_i;
wire signed [`CalcTempBus]          temp_m4_9_7_r;
wire signed [`CalcTempBus]          temp_m4_9_7_i;
wire signed [`CalcTempBus]          temp_m4_9_8_r;
wire signed [`CalcTempBus]          temp_m4_9_8_i;
wire signed [`CalcTempBus]          temp_m4_9_9_r;
wire signed [`CalcTempBus]          temp_m4_9_9_i;
wire signed [`CalcTempBus]          temp_m4_9_10_r;
wire signed [`CalcTempBus]          temp_m4_9_10_i;
wire signed [`CalcTempBus]          temp_m4_9_11_r;
wire signed [`CalcTempBus]          temp_m4_9_11_i;
wire signed [`CalcTempBus]          temp_m4_9_12_r;
wire signed [`CalcTempBus]          temp_m4_9_12_i;
wire signed [`CalcTempBus]          temp_m4_9_13_r;
wire signed [`CalcTempBus]          temp_m4_9_13_i;
wire signed [`CalcTempBus]          temp_m4_9_14_r;
wire signed [`CalcTempBus]          temp_m4_9_14_i;
wire signed [`CalcTempBus]          temp_m4_9_15_r;
wire signed [`CalcTempBus]          temp_m4_9_15_i;
wire signed [`CalcTempBus]          temp_m4_9_16_r;
wire signed [`CalcTempBus]          temp_m4_9_16_i;
wire signed [`CalcTempBus]          temp_m4_10_1_r;
wire signed [`CalcTempBus]          temp_m4_10_1_i;
wire signed [`CalcTempBus]          temp_m4_10_2_r;
wire signed [`CalcTempBus]          temp_m4_10_2_i;
wire signed [`CalcTempBus]          temp_m4_10_3_r;
wire signed [`CalcTempBus]          temp_m4_10_3_i;
wire signed [`CalcTempBus]          temp_m4_10_4_r;
wire signed [`CalcTempBus]          temp_m4_10_4_i;
wire signed [`CalcTempBus]          temp_m4_10_5_r;
wire signed [`CalcTempBus]          temp_m4_10_5_i;
wire signed [`CalcTempBus]          temp_m4_10_6_r;
wire signed [`CalcTempBus]          temp_m4_10_6_i;
wire signed [`CalcTempBus]          temp_m4_10_7_r;
wire signed [`CalcTempBus]          temp_m4_10_7_i;
wire signed [`CalcTempBus]          temp_m4_10_8_r;
wire signed [`CalcTempBus]          temp_m4_10_8_i;
wire signed [`CalcTempBus]          temp_m4_10_9_r;
wire signed [`CalcTempBus]          temp_m4_10_9_i;
wire signed [`CalcTempBus]          temp_m4_10_10_r;
wire signed [`CalcTempBus]          temp_m4_10_10_i;
wire signed [`CalcTempBus]          temp_m4_10_11_r;
wire signed [`CalcTempBus]          temp_m4_10_11_i;
wire signed [`CalcTempBus]          temp_m4_10_12_r;
wire signed [`CalcTempBus]          temp_m4_10_12_i;
wire signed [`CalcTempBus]          temp_m4_10_13_r;
wire signed [`CalcTempBus]          temp_m4_10_13_i;
wire signed [`CalcTempBus]          temp_m4_10_14_r;
wire signed [`CalcTempBus]          temp_m4_10_14_i;
wire signed [`CalcTempBus]          temp_m4_10_15_r;
wire signed [`CalcTempBus]          temp_m4_10_15_i;
wire signed [`CalcTempBus]          temp_m4_10_16_r;
wire signed [`CalcTempBus]          temp_m4_10_16_i;
wire signed [`CalcTempBus]          temp_m4_11_1_r;
wire signed [`CalcTempBus]          temp_m4_11_1_i;
wire signed [`CalcTempBus]          temp_m4_11_2_r;
wire signed [`CalcTempBus]          temp_m4_11_2_i;
wire signed [`CalcTempBus]          temp_m4_11_3_r;
wire signed [`CalcTempBus]          temp_m4_11_3_i;
wire signed [`CalcTempBus]          temp_m4_11_4_r;
wire signed [`CalcTempBus]          temp_m4_11_4_i;
wire signed [`CalcTempBus]          temp_m4_11_5_r;
wire signed [`CalcTempBus]          temp_m4_11_5_i;
wire signed [`CalcTempBus]          temp_m4_11_6_r;
wire signed [`CalcTempBus]          temp_m4_11_6_i;
wire signed [`CalcTempBus]          temp_m4_11_7_r;
wire signed [`CalcTempBus]          temp_m4_11_7_i;
wire signed [`CalcTempBus]          temp_m4_11_8_r;
wire signed [`CalcTempBus]          temp_m4_11_8_i;
wire signed [`CalcTempBus]          temp_m4_11_9_r;
wire signed [`CalcTempBus]          temp_m4_11_9_i;
wire signed [`CalcTempBus]          temp_m4_11_10_r;
wire signed [`CalcTempBus]          temp_m4_11_10_i;
wire signed [`CalcTempBus]          temp_m4_11_11_r;
wire signed [`CalcTempBus]          temp_m4_11_11_i;
wire signed [`CalcTempBus]          temp_m4_11_12_r;
wire signed [`CalcTempBus]          temp_m4_11_12_i;
wire signed [`CalcTempBus]          temp_m4_11_13_r;
wire signed [`CalcTempBus]          temp_m4_11_13_i;
wire signed [`CalcTempBus]          temp_m4_11_14_r;
wire signed [`CalcTempBus]          temp_m4_11_14_i;
wire signed [`CalcTempBus]          temp_m4_11_15_r;
wire signed [`CalcTempBus]          temp_m4_11_15_i;
wire signed [`CalcTempBus]          temp_m4_11_16_r;
wire signed [`CalcTempBus]          temp_m4_11_16_i;
wire signed [`CalcTempBus]          temp_m4_12_1_r;
wire signed [`CalcTempBus]          temp_m4_12_1_i;
wire signed [`CalcTempBus]          temp_m4_12_2_r;
wire signed [`CalcTempBus]          temp_m4_12_2_i;
wire signed [`CalcTempBus]          temp_m4_12_3_r;
wire signed [`CalcTempBus]          temp_m4_12_3_i;
wire signed [`CalcTempBus]          temp_m4_12_4_r;
wire signed [`CalcTempBus]          temp_m4_12_4_i;
wire signed [`CalcTempBus]          temp_m4_12_5_r;
wire signed [`CalcTempBus]          temp_m4_12_5_i;
wire signed [`CalcTempBus]          temp_m4_12_6_r;
wire signed [`CalcTempBus]          temp_m4_12_6_i;
wire signed [`CalcTempBus]          temp_m4_12_7_r;
wire signed [`CalcTempBus]          temp_m4_12_7_i;
wire signed [`CalcTempBus]          temp_m4_12_8_r;
wire signed [`CalcTempBus]          temp_m4_12_8_i;
wire signed [`CalcTempBus]          temp_m4_12_9_r;
wire signed [`CalcTempBus]          temp_m4_12_9_i;
wire signed [`CalcTempBus]          temp_m4_12_10_r;
wire signed [`CalcTempBus]          temp_m4_12_10_i;
wire signed [`CalcTempBus]          temp_m4_12_11_r;
wire signed [`CalcTempBus]          temp_m4_12_11_i;
wire signed [`CalcTempBus]          temp_m4_12_12_r;
wire signed [`CalcTempBus]          temp_m4_12_12_i;
wire signed [`CalcTempBus]          temp_m4_12_13_r;
wire signed [`CalcTempBus]          temp_m4_12_13_i;
wire signed [`CalcTempBus]          temp_m4_12_14_r;
wire signed [`CalcTempBus]          temp_m4_12_14_i;
wire signed [`CalcTempBus]          temp_m4_12_15_r;
wire signed [`CalcTempBus]          temp_m4_12_15_i;
wire signed [`CalcTempBus]          temp_m4_12_16_r;
wire signed [`CalcTempBus]          temp_m4_12_16_i;
wire signed [`CalcTempBus]          temp_m4_13_1_r;
wire signed [`CalcTempBus]          temp_m4_13_1_i;
wire signed [`CalcTempBus]          temp_m4_13_2_r;
wire signed [`CalcTempBus]          temp_m4_13_2_i;
wire signed [`CalcTempBus]          temp_m4_13_3_r;
wire signed [`CalcTempBus]          temp_m4_13_3_i;
wire signed [`CalcTempBus]          temp_m4_13_4_r;
wire signed [`CalcTempBus]          temp_m4_13_4_i;
wire signed [`CalcTempBus]          temp_m4_13_5_r;
wire signed [`CalcTempBus]          temp_m4_13_5_i;
wire signed [`CalcTempBus]          temp_m4_13_6_r;
wire signed [`CalcTempBus]          temp_m4_13_6_i;
wire signed [`CalcTempBus]          temp_m4_13_7_r;
wire signed [`CalcTempBus]          temp_m4_13_7_i;
wire signed [`CalcTempBus]          temp_m4_13_8_r;
wire signed [`CalcTempBus]          temp_m4_13_8_i;
wire signed [`CalcTempBus]          temp_m4_13_9_r;
wire signed [`CalcTempBus]          temp_m4_13_9_i;
wire signed [`CalcTempBus]          temp_m4_13_10_r;
wire signed [`CalcTempBus]          temp_m4_13_10_i;
wire signed [`CalcTempBus]          temp_m4_13_11_r;
wire signed [`CalcTempBus]          temp_m4_13_11_i;
wire signed [`CalcTempBus]          temp_m4_13_12_r;
wire signed [`CalcTempBus]          temp_m4_13_12_i;
wire signed [`CalcTempBus]          temp_m4_13_13_r;
wire signed [`CalcTempBus]          temp_m4_13_13_i;
wire signed [`CalcTempBus]          temp_m4_13_14_r;
wire signed [`CalcTempBus]          temp_m4_13_14_i;
wire signed [`CalcTempBus]          temp_m4_13_15_r;
wire signed [`CalcTempBus]          temp_m4_13_15_i;
wire signed [`CalcTempBus]          temp_m4_13_16_r;
wire signed [`CalcTempBus]          temp_m4_13_16_i;
wire signed [`CalcTempBus]          temp_m4_14_1_r;
wire signed [`CalcTempBus]          temp_m4_14_1_i;
wire signed [`CalcTempBus]          temp_m4_14_2_r;
wire signed [`CalcTempBus]          temp_m4_14_2_i;
wire signed [`CalcTempBus]          temp_m4_14_3_r;
wire signed [`CalcTempBus]          temp_m4_14_3_i;
wire signed [`CalcTempBus]          temp_m4_14_4_r;
wire signed [`CalcTempBus]          temp_m4_14_4_i;
wire signed [`CalcTempBus]          temp_m4_14_5_r;
wire signed [`CalcTempBus]          temp_m4_14_5_i;
wire signed [`CalcTempBus]          temp_m4_14_6_r;
wire signed [`CalcTempBus]          temp_m4_14_6_i;
wire signed [`CalcTempBus]          temp_m4_14_7_r;
wire signed [`CalcTempBus]          temp_m4_14_7_i;
wire signed [`CalcTempBus]          temp_m4_14_8_r;
wire signed [`CalcTempBus]          temp_m4_14_8_i;
wire signed [`CalcTempBus]          temp_m4_14_9_r;
wire signed [`CalcTempBus]          temp_m4_14_9_i;
wire signed [`CalcTempBus]          temp_m4_14_10_r;
wire signed [`CalcTempBus]          temp_m4_14_10_i;
wire signed [`CalcTempBus]          temp_m4_14_11_r;
wire signed [`CalcTempBus]          temp_m4_14_11_i;
wire signed [`CalcTempBus]          temp_m4_14_12_r;
wire signed [`CalcTempBus]          temp_m4_14_12_i;
wire signed [`CalcTempBus]          temp_m4_14_13_r;
wire signed [`CalcTempBus]          temp_m4_14_13_i;
wire signed [`CalcTempBus]          temp_m4_14_14_r;
wire signed [`CalcTempBus]          temp_m4_14_14_i;
wire signed [`CalcTempBus]          temp_m4_14_15_r;
wire signed [`CalcTempBus]          temp_m4_14_15_i;
wire signed [`CalcTempBus]          temp_m4_14_16_r;
wire signed [`CalcTempBus]          temp_m4_14_16_i;
wire signed [`CalcTempBus]          temp_m4_15_1_r;
wire signed [`CalcTempBus]          temp_m4_15_1_i;
wire signed [`CalcTempBus]          temp_m4_15_2_r;
wire signed [`CalcTempBus]          temp_m4_15_2_i;
wire signed [`CalcTempBus]          temp_m4_15_3_r;
wire signed [`CalcTempBus]          temp_m4_15_3_i;
wire signed [`CalcTempBus]          temp_m4_15_4_r;
wire signed [`CalcTempBus]          temp_m4_15_4_i;
wire signed [`CalcTempBus]          temp_m4_15_5_r;
wire signed [`CalcTempBus]          temp_m4_15_5_i;
wire signed [`CalcTempBus]          temp_m4_15_6_r;
wire signed [`CalcTempBus]          temp_m4_15_6_i;
wire signed [`CalcTempBus]          temp_m4_15_7_r;
wire signed [`CalcTempBus]          temp_m4_15_7_i;
wire signed [`CalcTempBus]          temp_m4_15_8_r;
wire signed [`CalcTempBus]          temp_m4_15_8_i;
wire signed [`CalcTempBus]          temp_m4_15_9_r;
wire signed [`CalcTempBus]          temp_m4_15_9_i;
wire signed [`CalcTempBus]          temp_m4_15_10_r;
wire signed [`CalcTempBus]          temp_m4_15_10_i;
wire signed [`CalcTempBus]          temp_m4_15_11_r;
wire signed [`CalcTempBus]          temp_m4_15_11_i;
wire signed [`CalcTempBus]          temp_m4_15_12_r;
wire signed [`CalcTempBus]          temp_m4_15_12_i;
wire signed [`CalcTempBus]          temp_m4_15_13_r;
wire signed [`CalcTempBus]          temp_m4_15_13_i;
wire signed [`CalcTempBus]          temp_m4_15_14_r;
wire signed [`CalcTempBus]          temp_m4_15_14_i;
wire signed [`CalcTempBus]          temp_m4_15_15_r;
wire signed [`CalcTempBus]          temp_m4_15_15_i;
wire signed [`CalcTempBus]          temp_m4_15_16_r;
wire signed [`CalcTempBus]          temp_m4_15_16_i;
wire signed [`CalcTempBus]          temp_m4_16_1_r;
wire signed [`CalcTempBus]          temp_m4_16_1_i;
wire signed [`CalcTempBus]          temp_m4_16_2_r;
wire signed [`CalcTempBus]          temp_m4_16_2_i;
wire signed [`CalcTempBus]          temp_m4_16_3_r;
wire signed [`CalcTempBus]          temp_m4_16_3_i;
wire signed [`CalcTempBus]          temp_m4_16_4_r;
wire signed [`CalcTempBus]          temp_m4_16_4_i;
wire signed [`CalcTempBus]          temp_m4_16_5_r;
wire signed [`CalcTempBus]          temp_m4_16_5_i;
wire signed [`CalcTempBus]          temp_m4_16_6_r;
wire signed [`CalcTempBus]          temp_m4_16_6_i;
wire signed [`CalcTempBus]          temp_m4_16_7_r;
wire signed [`CalcTempBus]          temp_m4_16_7_i;
wire signed [`CalcTempBus]          temp_m4_16_8_r;
wire signed [`CalcTempBus]          temp_m4_16_8_i;
wire signed [`CalcTempBus]          temp_m4_16_9_r;
wire signed [`CalcTempBus]          temp_m4_16_9_i;
wire signed [`CalcTempBus]          temp_m4_16_10_r;
wire signed [`CalcTempBus]          temp_m4_16_10_i;
wire signed [`CalcTempBus]          temp_m4_16_11_r;
wire signed [`CalcTempBus]          temp_m4_16_11_i;
wire signed [`CalcTempBus]          temp_m4_16_12_r;
wire signed [`CalcTempBus]          temp_m4_16_12_i;
wire signed [`CalcTempBus]          temp_m4_16_13_r;
wire signed [`CalcTempBus]          temp_m4_16_13_i;
wire signed [`CalcTempBus]          temp_m4_16_14_r;
wire signed [`CalcTempBus]          temp_m4_16_14_i;
wire signed [`CalcTempBus]          temp_m4_16_15_r;
wire signed [`CalcTempBus]          temp_m4_16_15_i;
wire signed [`CalcTempBus]          temp_m4_16_16_r;
wire signed [`CalcTempBus]          temp_m4_16_16_i;

wire signed [`CalcTempBus]          temp_b1_1_1_r;
wire signed [`CalcTempBus]          temp_b1_1_1_i;
wire signed [`CalcTempBus]          temp_b1_1_2_r;
wire signed [`CalcTempBus]          temp_b1_1_2_i;
wire signed [`CalcTempBus]          temp_b1_1_3_r;
wire signed [`CalcTempBus]          temp_b1_1_3_i;
wire signed [`CalcTempBus]          temp_b1_1_4_r;
wire signed [`CalcTempBus]          temp_b1_1_4_i;
wire signed [`CalcTempBus]          temp_b1_1_5_r;
wire signed [`CalcTempBus]          temp_b1_1_5_i;
wire signed [`CalcTempBus]          temp_b1_1_6_r;
wire signed [`CalcTempBus]          temp_b1_1_6_i;
wire signed [`CalcTempBus]          temp_b1_1_7_r;
wire signed [`CalcTempBus]          temp_b1_1_7_i;
wire signed [`CalcTempBus]          temp_b1_1_8_r;
wire signed [`CalcTempBus]          temp_b1_1_8_i;
wire signed [`CalcTempBus]          temp_b1_1_9_r;
wire signed [`CalcTempBus]          temp_b1_1_9_i;
wire signed [`CalcTempBus]          temp_b1_1_10_r;
wire signed [`CalcTempBus]          temp_b1_1_10_i;
wire signed [`CalcTempBus]          temp_b1_1_11_r;
wire signed [`CalcTempBus]          temp_b1_1_11_i;
wire signed [`CalcTempBus]          temp_b1_1_12_r;
wire signed [`CalcTempBus]          temp_b1_1_12_i;
wire signed [`CalcTempBus]          temp_b1_1_13_r;
wire signed [`CalcTempBus]          temp_b1_1_13_i;
wire signed [`CalcTempBus]          temp_b1_1_14_r;
wire signed [`CalcTempBus]          temp_b1_1_14_i;
wire signed [`CalcTempBus]          temp_b1_1_15_r;
wire signed [`CalcTempBus]          temp_b1_1_15_i;
wire signed [`CalcTempBus]          temp_b1_1_16_r;
wire signed [`CalcTempBus]          temp_b1_1_16_i;
wire signed [`CalcTempBus]          temp_b1_2_1_r;
wire signed [`CalcTempBus]          temp_b1_2_1_i;
wire signed [`CalcTempBus]          temp_b1_2_2_r;
wire signed [`CalcTempBus]          temp_b1_2_2_i;
wire signed [`CalcTempBus]          temp_b1_2_3_r;
wire signed [`CalcTempBus]          temp_b1_2_3_i;
wire signed [`CalcTempBus]          temp_b1_2_4_r;
wire signed [`CalcTempBus]          temp_b1_2_4_i;
wire signed [`CalcTempBus]          temp_b1_2_5_r;
wire signed [`CalcTempBus]          temp_b1_2_5_i;
wire signed [`CalcTempBus]          temp_b1_2_6_r;
wire signed [`CalcTempBus]          temp_b1_2_6_i;
wire signed [`CalcTempBus]          temp_b1_2_7_r;
wire signed [`CalcTempBus]          temp_b1_2_7_i;
wire signed [`CalcTempBus]          temp_b1_2_8_r;
wire signed [`CalcTempBus]          temp_b1_2_8_i;
wire signed [`CalcTempBus]          temp_b1_2_9_r;
wire signed [`CalcTempBus]          temp_b1_2_9_i;
wire signed [`CalcTempBus]          temp_b1_2_10_r;
wire signed [`CalcTempBus]          temp_b1_2_10_i;
wire signed [`CalcTempBus]          temp_b1_2_11_r;
wire signed [`CalcTempBus]          temp_b1_2_11_i;
wire signed [`CalcTempBus]          temp_b1_2_12_r;
wire signed [`CalcTempBus]          temp_b1_2_12_i;
wire signed [`CalcTempBus]          temp_b1_2_13_r;
wire signed [`CalcTempBus]          temp_b1_2_13_i;
wire signed [`CalcTempBus]          temp_b1_2_14_r;
wire signed [`CalcTempBus]          temp_b1_2_14_i;
wire signed [`CalcTempBus]          temp_b1_2_15_r;
wire signed [`CalcTempBus]          temp_b1_2_15_i;
wire signed [`CalcTempBus]          temp_b1_2_16_r;
wire signed [`CalcTempBus]          temp_b1_2_16_i;
wire signed [`CalcTempBus]          temp_b1_3_1_r;
wire signed [`CalcTempBus]          temp_b1_3_1_i;
wire signed [`CalcTempBus]          temp_b1_3_2_r;
wire signed [`CalcTempBus]          temp_b1_3_2_i;
wire signed [`CalcTempBus]          temp_b1_3_3_r;
wire signed [`CalcTempBus]          temp_b1_3_3_i;
wire signed [`CalcTempBus]          temp_b1_3_4_r;
wire signed [`CalcTempBus]          temp_b1_3_4_i;
wire signed [`CalcTempBus]          temp_b1_3_5_r;
wire signed [`CalcTempBus]          temp_b1_3_5_i;
wire signed [`CalcTempBus]          temp_b1_3_6_r;
wire signed [`CalcTempBus]          temp_b1_3_6_i;
wire signed [`CalcTempBus]          temp_b1_3_7_r;
wire signed [`CalcTempBus]          temp_b1_3_7_i;
wire signed [`CalcTempBus]          temp_b1_3_8_r;
wire signed [`CalcTempBus]          temp_b1_3_8_i;
wire signed [`CalcTempBus]          temp_b1_3_9_r;
wire signed [`CalcTempBus]          temp_b1_3_9_i;
wire signed [`CalcTempBus]          temp_b1_3_10_r;
wire signed [`CalcTempBus]          temp_b1_3_10_i;
wire signed [`CalcTempBus]          temp_b1_3_11_r;
wire signed [`CalcTempBus]          temp_b1_3_11_i;
wire signed [`CalcTempBus]          temp_b1_3_12_r;
wire signed [`CalcTempBus]          temp_b1_3_12_i;
wire signed [`CalcTempBus]          temp_b1_3_13_r;
wire signed [`CalcTempBus]          temp_b1_3_13_i;
wire signed [`CalcTempBus]          temp_b1_3_14_r;
wire signed [`CalcTempBus]          temp_b1_3_14_i;
wire signed [`CalcTempBus]          temp_b1_3_15_r;
wire signed [`CalcTempBus]          temp_b1_3_15_i;
wire signed [`CalcTempBus]          temp_b1_3_16_r;
wire signed [`CalcTempBus]          temp_b1_3_16_i;
wire signed [`CalcTempBus]          temp_b1_4_1_r;
wire signed [`CalcTempBus]          temp_b1_4_1_i;
wire signed [`CalcTempBus]          temp_b1_4_2_r;
wire signed [`CalcTempBus]          temp_b1_4_2_i;
wire signed [`CalcTempBus]          temp_b1_4_3_r;
wire signed [`CalcTempBus]          temp_b1_4_3_i;
wire signed [`CalcTempBus]          temp_b1_4_4_r;
wire signed [`CalcTempBus]          temp_b1_4_4_i;
wire signed [`CalcTempBus]          temp_b1_4_5_r;
wire signed [`CalcTempBus]          temp_b1_4_5_i;
wire signed [`CalcTempBus]          temp_b1_4_6_r;
wire signed [`CalcTempBus]          temp_b1_4_6_i;
wire signed [`CalcTempBus]          temp_b1_4_7_r;
wire signed [`CalcTempBus]          temp_b1_4_7_i;
wire signed [`CalcTempBus]          temp_b1_4_8_r;
wire signed [`CalcTempBus]          temp_b1_4_8_i;
wire signed [`CalcTempBus]          temp_b1_4_9_r;
wire signed [`CalcTempBus]          temp_b1_4_9_i;
wire signed [`CalcTempBus]          temp_b1_4_10_r;
wire signed [`CalcTempBus]          temp_b1_4_10_i;
wire signed [`CalcTempBus]          temp_b1_4_11_r;
wire signed [`CalcTempBus]          temp_b1_4_11_i;
wire signed [`CalcTempBus]          temp_b1_4_12_r;
wire signed [`CalcTempBus]          temp_b1_4_12_i;
wire signed [`CalcTempBus]          temp_b1_4_13_r;
wire signed [`CalcTempBus]          temp_b1_4_13_i;
wire signed [`CalcTempBus]          temp_b1_4_14_r;
wire signed [`CalcTempBus]          temp_b1_4_14_i;
wire signed [`CalcTempBus]          temp_b1_4_15_r;
wire signed [`CalcTempBus]          temp_b1_4_15_i;
wire signed [`CalcTempBus]          temp_b1_4_16_r;
wire signed [`CalcTempBus]          temp_b1_4_16_i;
wire signed [`CalcTempBus]          temp_b1_5_1_r;
wire signed [`CalcTempBus]          temp_b1_5_1_i;
wire signed [`CalcTempBus]          temp_b1_5_2_r;
wire signed [`CalcTempBus]          temp_b1_5_2_i;
wire signed [`CalcTempBus]          temp_b1_5_3_r;
wire signed [`CalcTempBus]          temp_b1_5_3_i;
wire signed [`CalcTempBus]          temp_b1_5_4_r;
wire signed [`CalcTempBus]          temp_b1_5_4_i;
wire signed [`CalcTempBus]          temp_b1_5_5_r;
wire signed [`CalcTempBus]          temp_b1_5_5_i;
wire signed [`CalcTempBus]          temp_b1_5_6_r;
wire signed [`CalcTempBus]          temp_b1_5_6_i;
wire signed [`CalcTempBus]          temp_b1_5_7_r;
wire signed [`CalcTempBus]          temp_b1_5_7_i;
wire signed [`CalcTempBus]          temp_b1_5_8_r;
wire signed [`CalcTempBus]          temp_b1_5_8_i;
wire signed [`CalcTempBus]          temp_b1_5_9_r;
wire signed [`CalcTempBus]          temp_b1_5_9_i;
wire signed [`CalcTempBus]          temp_b1_5_10_r;
wire signed [`CalcTempBus]          temp_b1_5_10_i;
wire signed [`CalcTempBus]          temp_b1_5_11_r;
wire signed [`CalcTempBus]          temp_b1_5_11_i;
wire signed [`CalcTempBus]          temp_b1_5_12_r;
wire signed [`CalcTempBus]          temp_b1_5_12_i;
wire signed [`CalcTempBus]          temp_b1_5_13_r;
wire signed [`CalcTempBus]          temp_b1_5_13_i;
wire signed [`CalcTempBus]          temp_b1_5_14_r;
wire signed [`CalcTempBus]          temp_b1_5_14_i;
wire signed [`CalcTempBus]          temp_b1_5_15_r;
wire signed [`CalcTempBus]          temp_b1_5_15_i;
wire signed [`CalcTempBus]          temp_b1_5_16_r;
wire signed [`CalcTempBus]          temp_b1_5_16_i;
wire signed [`CalcTempBus]          temp_b1_6_1_r;
wire signed [`CalcTempBus]          temp_b1_6_1_i;
wire signed [`CalcTempBus]          temp_b1_6_2_r;
wire signed [`CalcTempBus]          temp_b1_6_2_i;
wire signed [`CalcTempBus]          temp_b1_6_3_r;
wire signed [`CalcTempBus]          temp_b1_6_3_i;
wire signed [`CalcTempBus]          temp_b1_6_4_r;
wire signed [`CalcTempBus]          temp_b1_6_4_i;
wire signed [`CalcTempBus]          temp_b1_6_5_r;
wire signed [`CalcTempBus]          temp_b1_6_5_i;
wire signed [`CalcTempBus]          temp_b1_6_6_r;
wire signed [`CalcTempBus]          temp_b1_6_6_i;
wire signed [`CalcTempBus]          temp_b1_6_7_r;
wire signed [`CalcTempBus]          temp_b1_6_7_i;
wire signed [`CalcTempBus]          temp_b1_6_8_r;
wire signed [`CalcTempBus]          temp_b1_6_8_i;
wire signed [`CalcTempBus]          temp_b1_6_9_r;
wire signed [`CalcTempBus]          temp_b1_6_9_i;
wire signed [`CalcTempBus]          temp_b1_6_10_r;
wire signed [`CalcTempBus]          temp_b1_6_10_i;
wire signed [`CalcTempBus]          temp_b1_6_11_r;
wire signed [`CalcTempBus]          temp_b1_6_11_i;
wire signed [`CalcTempBus]          temp_b1_6_12_r;
wire signed [`CalcTempBus]          temp_b1_6_12_i;
wire signed [`CalcTempBus]          temp_b1_6_13_r;
wire signed [`CalcTempBus]          temp_b1_6_13_i;
wire signed [`CalcTempBus]          temp_b1_6_14_r;
wire signed [`CalcTempBus]          temp_b1_6_14_i;
wire signed [`CalcTempBus]          temp_b1_6_15_r;
wire signed [`CalcTempBus]          temp_b1_6_15_i;
wire signed [`CalcTempBus]          temp_b1_6_16_r;
wire signed [`CalcTempBus]          temp_b1_6_16_i;
wire signed [`CalcTempBus]          temp_b1_7_1_r;
wire signed [`CalcTempBus]          temp_b1_7_1_i;
wire signed [`CalcTempBus]          temp_b1_7_2_r;
wire signed [`CalcTempBus]          temp_b1_7_2_i;
wire signed [`CalcTempBus]          temp_b1_7_3_r;
wire signed [`CalcTempBus]          temp_b1_7_3_i;
wire signed [`CalcTempBus]          temp_b1_7_4_r;
wire signed [`CalcTempBus]          temp_b1_7_4_i;
wire signed [`CalcTempBus]          temp_b1_7_5_r;
wire signed [`CalcTempBus]          temp_b1_7_5_i;
wire signed [`CalcTempBus]          temp_b1_7_6_r;
wire signed [`CalcTempBus]          temp_b1_7_6_i;
wire signed [`CalcTempBus]          temp_b1_7_7_r;
wire signed [`CalcTempBus]          temp_b1_7_7_i;
wire signed [`CalcTempBus]          temp_b1_7_8_r;
wire signed [`CalcTempBus]          temp_b1_7_8_i;
wire signed [`CalcTempBus]          temp_b1_7_9_r;
wire signed [`CalcTempBus]          temp_b1_7_9_i;
wire signed [`CalcTempBus]          temp_b1_7_10_r;
wire signed [`CalcTempBus]          temp_b1_7_10_i;
wire signed [`CalcTempBus]          temp_b1_7_11_r;
wire signed [`CalcTempBus]          temp_b1_7_11_i;
wire signed [`CalcTempBus]          temp_b1_7_12_r;
wire signed [`CalcTempBus]          temp_b1_7_12_i;
wire signed [`CalcTempBus]          temp_b1_7_13_r;
wire signed [`CalcTempBus]          temp_b1_7_13_i;
wire signed [`CalcTempBus]          temp_b1_7_14_r;
wire signed [`CalcTempBus]          temp_b1_7_14_i;
wire signed [`CalcTempBus]          temp_b1_7_15_r;
wire signed [`CalcTempBus]          temp_b1_7_15_i;
wire signed [`CalcTempBus]          temp_b1_7_16_r;
wire signed [`CalcTempBus]          temp_b1_7_16_i;
wire signed [`CalcTempBus]          temp_b1_8_1_r;
wire signed [`CalcTempBus]          temp_b1_8_1_i;
wire signed [`CalcTempBus]          temp_b1_8_2_r;
wire signed [`CalcTempBus]          temp_b1_8_2_i;
wire signed [`CalcTempBus]          temp_b1_8_3_r;
wire signed [`CalcTempBus]          temp_b1_8_3_i;
wire signed [`CalcTempBus]          temp_b1_8_4_r;
wire signed [`CalcTempBus]          temp_b1_8_4_i;
wire signed [`CalcTempBus]          temp_b1_8_5_r;
wire signed [`CalcTempBus]          temp_b1_8_5_i;
wire signed [`CalcTempBus]          temp_b1_8_6_r;
wire signed [`CalcTempBus]          temp_b1_8_6_i;
wire signed [`CalcTempBus]          temp_b1_8_7_r;
wire signed [`CalcTempBus]          temp_b1_8_7_i;
wire signed [`CalcTempBus]          temp_b1_8_8_r;
wire signed [`CalcTempBus]          temp_b1_8_8_i;
wire signed [`CalcTempBus]          temp_b1_8_9_r;
wire signed [`CalcTempBus]          temp_b1_8_9_i;
wire signed [`CalcTempBus]          temp_b1_8_10_r;
wire signed [`CalcTempBus]          temp_b1_8_10_i;
wire signed [`CalcTempBus]          temp_b1_8_11_r;
wire signed [`CalcTempBus]          temp_b1_8_11_i;
wire signed [`CalcTempBus]          temp_b1_8_12_r;
wire signed [`CalcTempBus]          temp_b1_8_12_i;
wire signed [`CalcTempBus]          temp_b1_8_13_r;
wire signed [`CalcTempBus]          temp_b1_8_13_i;
wire signed [`CalcTempBus]          temp_b1_8_14_r;
wire signed [`CalcTempBus]          temp_b1_8_14_i;
wire signed [`CalcTempBus]          temp_b1_8_15_r;
wire signed [`CalcTempBus]          temp_b1_8_15_i;
wire signed [`CalcTempBus]          temp_b1_8_16_r;
wire signed [`CalcTempBus]          temp_b1_8_16_i;
wire signed [`CalcTempBus]          temp_b1_9_1_r;
wire signed [`CalcTempBus]          temp_b1_9_1_i;
wire signed [`CalcTempBus]          temp_b1_9_2_r;
wire signed [`CalcTempBus]          temp_b1_9_2_i;
wire signed [`CalcTempBus]          temp_b1_9_3_r;
wire signed [`CalcTempBus]          temp_b1_9_3_i;
wire signed [`CalcTempBus]          temp_b1_9_4_r;
wire signed [`CalcTempBus]          temp_b1_9_4_i;
wire signed [`CalcTempBus]          temp_b1_9_5_r;
wire signed [`CalcTempBus]          temp_b1_9_5_i;
wire signed [`CalcTempBus]          temp_b1_9_6_r;
wire signed [`CalcTempBus]          temp_b1_9_6_i;
wire signed [`CalcTempBus]          temp_b1_9_7_r;
wire signed [`CalcTempBus]          temp_b1_9_7_i;
wire signed [`CalcTempBus]          temp_b1_9_8_r;
wire signed [`CalcTempBus]          temp_b1_9_8_i;
wire signed [`CalcTempBus]          temp_b1_9_9_r;
wire signed [`CalcTempBus]          temp_b1_9_9_i;
wire signed [`CalcTempBus]          temp_b1_9_10_r;
wire signed [`CalcTempBus]          temp_b1_9_10_i;
wire signed [`CalcTempBus]          temp_b1_9_11_r;
wire signed [`CalcTempBus]          temp_b1_9_11_i;
wire signed [`CalcTempBus]          temp_b1_9_12_r;
wire signed [`CalcTempBus]          temp_b1_9_12_i;
wire signed [`CalcTempBus]          temp_b1_9_13_r;
wire signed [`CalcTempBus]          temp_b1_9_13_i;
wire signed [`CalcTempBus]          temp_b1_9_14_r;
wire signed [`CalcTempBus]          temp_b1_9_14_i;
wire signed [`CalcTempBus]          temp_b1_9_15_r;
wire signed [`CalcTempBus]          temp_b1_9_15_i;
wire signed [`CalcTempBus]          temp_b1_9_16_r;
wire signed [`CalcTempBus]          temp_b1_9_16_i;
wire signed [`CalcTempBus]          temp_b1_10_1_r;
wire signed [`CalcTempBus]          temp_b1_10_1_i;
wire signed [`CalcTempBus]          temp_b1_10_2_r;
wire signed [`CalcTempBus]          temp_b1_10_2_i;
wire signed [`CalcTempBus]          temp_b1_10_3_r;
wire signed [`CalcTempBus]          temp_b1_10_3_i;
wire signed [`CalcTempBus]          temp_b1_10_4_r;
wire signed [`CalcTempBus]          temp_b1_10_4_i;
wire signed [`CalcTempBus]          temp_b1_10_5_r;
wire signed [`CalcTempBus]          temp_b1_10_5_i;
wire signed [`CalcTempBus]          temp_b1_10_6_r;
wire signed [`CalcTempBus]          temp_b1_10_6_i;
wire signed [`CalcTempBus]          temp_b1_10_7_r;
wire signed [`CalcTempBus]          temp_b1_10_7_i;
wire signed [`CalcTempBus]          temp_b1_10_8_r;
wire signed [`CalcTempBus]          temp_b1_10_8_i;
wire signed [`CalcTempBus]          temp_b1_10_9_r;
wire signed [`CalcTempBus]          temp_b1_10_9_i;
wire signed [`CalcTempBus]          temp_b1_10_10_r;
wire signed [`CalcTempBus]          temp_b1_10_10_i;
wire signed [`CalcTempBus]          temp_b1_10_11_r;
wire signed [`CalcTempBus]          temp_b1_10_11_i;
wire signed [`CalcTempBus]          temp_b1_10_12_r;
wire signed [`CalcTempBus]          temp_b1_10_12_i;
wire signed [`CalcTempBus]          temp_b1_10_13_r;
wire signed [`CalcTempBus]          temp_b1_10_13_i;
wire signed [`CalcTempBus]          temp_b1_10_14_r;
wire signed [`CalcTempBus]          temp_b1_10_14_i;
wire signed [`CalcTempBus]          temp_b1_10_15_r;
wire signed [`CalcTempBus]          temp_b1_10_15_i;
wire signed [`CalcTempBus]          temp_b1_10_16_r;
wire signed [`CalcTempBus]          temp_b1_10_16_i;
wire signed [`CalcTempBus]          temp_b1_11_1_r;
wire signed [`CalcTempBus]          temp_b1_11_1_i;
wire signed [`CalcTempBus]          temp_b1_11_2_r;
wire signed [`CalcTempBus]          temp_b1_11_2_i;
wire signed [`CalcTempBus]          temp_b1_11_3_r;
wire signed [`CalcTempBus]          temp_b1_11_3_i;
wire signed [`CalcTempBus]          temp_b1_11_4_r;
wire signed [`CalcTempBus]          temp_b1_11_4_i;
wire signed [`CalcTempBus]          temp_b1_11_5_r;
wire signed [`CalcTempBus]          temp_b1_11_5_i;
wire signed [`CalcTempBus]          temp_b1_11_6_r;
wire signed [`CalcTempBus]          temp_b1_11_6_i;
wire signed [`CalcTempBus]          temp_b1_11_7_r;
wire signed [`CalcTempBus]          temp_b1_11_7_i;
wire signed [`CalcTempBus]          temp_b1_11_8_r;
wire signed [`CalcTempBus]          temp_b1_11_8_i;
wire signed [`CalcTempBus]          temp_b1_11_9_r;
wire signed [`CalcTempBus]          temp_b1_11_9_i;
wire signed [`CalcTempBus]          temp_b1_11_10_r;
wire signed [`CalcTempBus]          temp_b1_11_10_i;
wire signed [`CalcTempBus]          temp_b1_11_11_r;
wire signed [`CalcTempBus]          temp_b1_11_11_i;
wire signed [`CalcTempBus]          temp_b1_11_12_r;
wire signed [`CalcTempBus]          temp_b1_11_12_i;
wire signed [`CalcTempBus]          temp_b1_11_13_r;
wire signed [`CalcTempBus]          temp_b1_11_13_i;
wire signed [`CalcTempBus]          temp_b1_11_14_r;
wire signed [`CalcTempBus]          temp_b1_11_14_i;
wire signed [`CalcTempBus]          temp_b1_11_15_r;
wire signed [`CalcTempBus]          temp_b1_11_15_i;
wire signed [`CalcTempBus]          temp_b1_11_16_r;
wire signed [`CalcTempBus]          temp_b1_11_16_i;
wire signed [`CalcTempBus]          temp_b1_12_1_r;
wire signed [`CalcTempBus]          temp_b1_12_1_i;
wire signed [`CalcTempBus]          temp_b1_12_2_r;
wire signed [`CalcTempBus]          temp_b1_12_2_i;
wire signed [`CalcTempBus]          temp_b1_12_3_r;
wire signed [`CalcTempBus]          temp_b1_12_3_i;
wire signed [`CalcTempBus]          temp_b1_12_4_r;
wire signed [`CalcTempBus]          temp_b1_12_4_i;
wire signed [`CalcTempBus]          temp_b1_12_5_r;
wire signed [`CalcTempBus]          temp_b1_12_5_i;
wire signed [`CalcTempBus]          temp_b1_12_6_r;
wire signed [`CalcTempBus]          temp_b1_12_6_i;
wire signed [`CalcTempBus]          temp_b1_12_7_r;
wire signed [`CalcTempBus]          temp_b1_12_7_i;
wire signed [`CalcTempBus]          temp_b1_12_8_r;
wire signed [`CalcTempBus]          temp_b1_12_8_i;
wire signed [`CalcTempBus]          temp_b1_12_9_r;
wire signed [`CalcTempBus]          temp_b1_12_9_i;
wire signed [`CalcTempBus]          temp_b1_12_10_r;
wire signed [`CalcTempBus]          temp_b1_12_10_i;
wire signed [`CalcTempBus]          temp_b1_12_11_r;
wire signed [`CalcTempBus]          temp_b1_12_11_i;
wire signed [`CalcTempBus]          temp_b1_12_12_r;
wire signed [`CalcTempBus]          temp_b1_12_12_i;
wire signed [`CalcTempBus]          temp_b1_12_13_r;
wire signed [`CalcTempBus]          temp_b1_12_13_i;
wire signed [`CalcTempBus]          temp_b1_12_14_r;
wire signed [`CalcTempBus]          temp_b1_12_14_i;
wire signed [`CalcTempBus]          temp_b1_12_15_r;
wire signed [`CalcTempBus]          temp_b1_12_15_i;
wire signed [`CalcTempBus]          temp_b1_12_16_r;
wire signed [`CalcTempBus]          temp_b1_12_16_i;
wire signed [`CalcTempBus]          temp_b1_13_1_r;
wire signed [`CalcTempBus]          temp_b1_13_1_i;
wire signed [`CalcTempBus]          temp_b1_13_2_r;
wire signed [`CalcTempBus]          temp_b1_13_2_i;
wire signed [`CalcTempBus]          temp_b1_13_3_r;
wire signed [`CalcTempBus]          temp_b1_13_3_i;
wire signed [`CalcTempBus]          temp_b1_13_4_r;
wire signed [`CalcTempBus]          temp_b1_13_4_i;
wire signed [`CalcTempBus]          temp_b1_13_5_r;
wire signed [`CalcTempBus]          temp_b1_13_5_i;
wire signed [`CalcTempBus]          temp_b1_13_6_r;
wire signed [`CalcTempBus]          temp_b1_13_6_i;
wire signed [`CalcTempBus]          temp_b1_13_7_r;
wire signed [`CalcTempBus]          temp_b1_13_7_i;
wire signed [`CalcTempBus]          temp_b1_13_8_r;
wire signed [`CalcTempBus]          temp_b1_13_8_i;
wire signed [`CalcTempBus]          temp_b1_13_9_r;
wire signed [`CalcTempBus]          temp_b1_13_9_i;
wire signed [`CalcTempBus]          temp_b1_13_10_r;
wire signed [`CalcTempBus]          temp_b1_13_10_i;
wire signed [`CalcTempBus]          temp_b1_13_11_r;
wire signed [`CalcTempBus]          temp_b1_13_11_i;
wire signed [`CalcTempBus]          temp_b1_13_12_r;
wire signed [`CalcTempBus]          temp_b1_13_12_i;
wire signed [`CalcTempBus]          temp_b1_13_13_r;
wire signed [`CalcTempBus]          temp_b1_13_13_i;
wire signed [`CalcTempBus]          temp_b1_13_14_r;
wire signed [`CalcTempBus]          temp_b1_13_14_i;
wire signed [`CalcTempBus]          temp_b1_13_15_r;
wire signed [`CalcTempBus]          temp_b1_13_15_i;
wire signed [`CalcTempBus]          temp_b1_13_16_r;
wire signed [`CalcTempBus]          temp_b1_13_16_i;
wire signed [`CalcTempBus]          temp_b1_14_1_r;
wire signed [`CalcTempBus]          temp_b1_14_1_i;
wire signed [`CalcTempBus]          temp_b1_14_2_r;
wire signed [`CalcTempBus]          temp_b1_14_2_i;
wire signed [`CalcTempBus]          temp_b1_14_3_r;
wire signed [`CalcTempBus]          temp_b1_14_3_i;
wire signed [`CalcTempBus]          temp_b1_14_4_r;
wire signed [`CalcTempBus]          temp_b1_14_4_i;
wire signed [`CalcTempBus]          temp_b1_14_5_r;
wire signed [`CalcTempBus]          temp_b1_14_5_i;
wire signed [`CalcTempBus]          temp_b1_14_6_r;
wire signed [`CalcTempBus]          temp_b1_14_6_i;
wire signed [`CalcTempBus]          temp_b1_14_7_r;
wire signed [`CalcTempBus]          temp_b1_14_7_i;
wire signed [`CalcTempBus]          temp_b1_14_8_r;
wire signed [`CalcTempBus]          temp_b1_14_8_i;
wire signed [`CalcTempBus]          temp_b1_14_9_r;
wire signed [`CalcTempBus]          temp_b1_14_9_i;
wire signed [`CalcTempBus]          temp_b1_14_10_r;
wire signed [`CalcTempBus]          temp_b1_14_10_i;
wire signed [`CalcTempBus]          temp_b1_14_11_r;
wire signed [`CalcTempBus]          temp_b1_14_11_i;
wire signed [`CalcTempBus]          temp_b1_14_12_r;
wire signed [`CalcTempBus]          temp_b1_14_12_i;
wire signed [`CalcTempBus]          temp_b1_14_13_r;
wire signed [`CalcTempBus]          temp_b1_14_13_i;
wire signed [`CalcTempBus]          temp_b1_14_14_r;
wire signed [`CalcTempBus]          temp_b1_14_14_i;
wire signed [`CalcTempBus]          temp_b1_14_15_r;
wire signed [`CalcTempBus]          temp_b1_14_15_i;
wire signed [`CalcTempBus]          temp_b1_14_16_r;
wire signed [`CalcTempBus]          temp_b1_14_16_i;
wire signed [`CalcTempBus]          temp_b1_15_1_r;
wire signed [`CalcTempBus]          temp_b1_15_1_i;
wire signed [`CalcTempBus]          temp_b1_15_2_r;
wire signed [`CalcTempBus]          temp_b1_15_2_i;
wire signed [`CalcTempBus]          temp_b1_15_3_r;
wire signed [`CalcTempBus]          temp_b1_15_3_i;
wire signed [`CalcTempBus]          temp_b1_15_4_r;
wire signed [`CalcTempBus]          temp_b1_15_4_i;
wire signed [`CalcTempBus]          temp_b1_15_5_r;
wire signed [`CalcTempBus]          temp_b1_15_5_i;
wire signed [`CalcTempBus]          temp_b1_15_6_r;
wire signed [`CalcTempBus]          temp_b1_15_6_i;
wire signed [`CalcTempBus]          temp_b1_15_7_r;
wire signed [`CalcTempBus]          temp_b1_15_7_i;
wire signed [`CalcTempBus]          temp_b1_15_8_r;
wire signed [`CalcTempBus]          temp_b1_15_8_i;
wire signed [`CalcTempBus]          temp_b1_15_9_r;
wire signed [`CalcTempBus]          temp_b1_15_9_i;
wire signed [`CalcTempBus]          temp_b1_15_10_r;
wire signed [`CalcTempBus]          temp_b1_15_10_i;
wire signed [`CalcTempBus]          temp_b1_15_11_r;
wire signed [`CalcTempBus]          temp_b1_15_11_i;
wire signed [`CalcTempBus]          temp_b1_15_12_r;
wire signed [`CalcTempBus]          temp_b1_15_12_i;
wire signed [`CalcTempBus]          temp_b1_15_13_r;
wire signed [`CalcTempBus]          temp_b1_15_13_i;
wire signed [`CalcTempBus]          temp_b1_15_14_r;
wire signed [`CalcTempBus]          temp_b1_15_14_i;
wire signed [`CalcTempBus]          temp_b1_15_15_r;
wire signed [`CalcTempBus]          temp_b1_15_15_i;
wire signed [`CalcTempBus]          temp_b1_15_16_r;
wire signed [`CalcTempBus]          temp_b1_15_16_i;
wire signed [`CalcTempBus]          temp_b1_16_1_r;
wire signed [`CalcTempBus]          temp_b1_16_1_i;
wire signed [`CalcTempBus]          temp_b1_16_2_r;
wire signed [`CalcTempBus]          temp_b1_16_2_i;
wire signed [`CalcTempBus]          temp_b1_16_3_r;
wire signed [`CalcTempBus]          temp_b1_16_3_i;
wire signed [`CalcTempBus]          temp_b1_16_4_r;
wire signed [`CalcTempBus]          temp_b1_16_4_i;
wire signed [`CalcTempBus]          temp_b1_16_5_r;
wire signed [`CalcTempBus]          temp_b1_16_5_i;
wire signed [`CalcTempBus]          temp_b1_16_6_r;
wire signed [`CalcTempBus]          temp_b1_16_6_i;
wire signed [`CalcTempBus]          temp_b1_16_7_r;
wire signed [`CalcTempBus]          temp_b1_16_7_i;
wire signed [`CalcTempBus]          temp_b1_16_8_r;
wire signed [`CalcTempBus]          temp_b1_16_8_i;
wire signed [`CalcTempBus]          temp_b1_16_9_r;
wire signed [`CalcTempBus]          temp_b1_16_9_i;
wire signed [`CalcTempBus]          temp_b1_16_10_r;
wire signed [`CalcTempBus]          temp_b1_16_10_i;
wire signed [`CalcTempBus]          temp_b1_16_11_r;
wire signed [`CalcTempBus]          temp_b1_16_11_i;
wire signed [`CalcTempBus]          temp_b1_16_12_r;
wire signed [`CalcTempBus]          temp_b1_16_12_i;
wire signed [`CalcTempBus]          temp_b1_16_13_r;
wire signed [`CalcTempBus]          temp_b1_16_13_i;
wire signed [`CalcTempBus]          temp_b1_16_14_r;
wire signed [`CalcTempBus]          temp_b1_16_14_i;
wire signed [`CalcTempBus]          temp_b1_16_15_r;
wire signed [`CalcTempBus]          temp_b1_16_15_i;
wire signed [`CalcTempBus]          temp_b1_16_16_r;
wire signed [`CalcTempBus]          temp_b1_16_16_i;
wire signed [`CalcTempBus]          temp_b2_1_1_r;
wire signed [`CalcTempBus]          temp_b2_1_1_i;
wire signed [`CalcTempBus]          temp_b2_1_2_r;
wire signed [`CalcTempBus]          temp_b2_1_2_i;
wire signed [`CalcTempBus]          temp_b2_1_3_r;
wire signed [`CalcTempBus]          temp_b2_1_3_i;
wire signed [`CalcTempBus]          temp_b2_1_4_r;
wire signed [`CalcTempBus]          temp_b2_1_4_i;
wire signed [`CalcTempBus]          temp_b2_1_5_r;
wire signed [`CalcTempBus]          temp_b2_1_5_i;
wire signed [`CalcTempBus]          temp_b2_1_6_r;
wire signed [`CalcTempBus]          temp_b2_1_6_i;
wire signed [`CalcTempBus]          temp_b2_1_7_r;
wire signed [`CalcTempBus]          temp_b2_1_7_i;
wire signed [`CalcTempBus]          temp_b2_1_8_r;
wire signed [`CalcTempBus]          temp_b2_1_8_i;
wire signed [`CalcTempBus]          temp_b2_1_9_r;
wire signed [`CalcTempBus]          temp_b2_1_9_i;
wire signed [`CalcTempBus]          temp_b2_1_10_r;
wire signed [`CalcTempBus]          temp_b2_1_10_i;
wire signed [`CalcTempBus]          temp_b2_1_11_r;
wire signed [`CalcTempBus]          temp_b2_1_11_i;
wire signed [`CalcTempBus]          temp_b2_1_12_r;
wire signed [`CalcTempBus]          temp_b2_1_12_i;
wire signed [`CalcTempBus]          temp_b2_1_13_r;
wire signed [`CalcTempBus]          temp_b2_1_13_i;
wire signed [`CalcTempBus]          temp_b2_1_14_r;
wire signed [`CalcTempBus]          temp_b2_1_14_i;
wire signed [`CalcTempBus]          temp_b2_1_15_r;
wire signed [`CalcTempBus]          temp_b2_1_15_i;
wire signed [`CalcTempBus]          temp_b2_1_16_r;
wire signed [`CalcTempBus]          temp_b2_1_16_i;
wire signed [`CalcTempBus]          temp_b2_2_1_r;
wire signed [`CalcTempBus]          temp_b2_2_1_i;
wire signed [`CalcTempBus]          temp_b2_2_2_r;
wire signed [`CalcTempBus]          temp_b2_2_2_i;
wire signed [`CalcTempBus]          temp_b2_2_3_r;
wire signed [`CalcTempBus]          temp_b2_2_3_i;
wire signed [`CalcTempBus]          temp_b2_2_4_r;
wire signed [`CalcTempBus]          temp_b2_2_4_i;
wire signed [`CalcTempBus]          temp_b2_2_5_r;
wire signed [`CalcTempBus]          temp_b2_2_5_i;
wire signed [`CalcTempBus]          temp_b2_2_6_r;
wire signed [`CalcTempBus]          temp_b2_2_6_i;
wire signed [`CalcTempBus]          temp_b2_2_7_r;
wire signed [`CalcTempBus]          temp_b2_2_7_i;
wire signed [`CalcTempBus]          temp_b2_2_8_r;
wire signed [`CalcTempBus]          temp_b2_2_8_i;
wire signed [`CalcTempBus]          temp_b2_2_9_r;
wire signed [`CalcTempBus]          temp_b2_2_9_i;
wire signed [`CalcTempBus]          temp_b2_2_10_r;
wire signed [`CalcTempBus]          temp_b2_2_10_i;
wire signed [`CalcTempBus]          temp_b2_2_11_r;
wire signed [`CalcTempBus]          temp_b2_2_11_i;
wire signed [`CalcTempBus]          temp_b2_2_12_r;
wire signed [`CalcTempBus]          temp_b2_2_12_i;
wire signed [`CalcTempBus]          temp_b2_2_13_r;
wire signed [`CalcTempBus]          temp_b2_2_13_i;
wire signed [`CalcTempBus]          temp_b2_2_14_r;
wire signed [`CalcTempBus]          temp_b2_2_14_i;
wire signed [`CalcTempBus]          temp_b2_2_15_r;
wire signed [`CalcTempBus]          temp_b2_2_15_i;
wire signed [`CalcTempBus]          temp_b2_2_16_r;
wire signed [`CalcTempBus]          temp_b2_2_16_i;
wire signed [`CalcTempBus]          temp_b2_3_1_r;
wire signed [`CalcTempBus]          temp_b2_3_1_i;
wire signed [`CalcTempBus]          temp_b2_3_2_r;
wire signed [`CalcTempBus]          temp_b2_3_2_i;
wire signed [`CalcTempBus]          temp_b2_3_3_r;
wire signed [`CalcTempBus]          temp_b2_3_3_i;
wire signed [`CalcTempBus]          temp_b2_3_4_r;
wire signed [`CalcTempBus]          temp_b2_3_4_i;
wire signed [`CalcTempBus]          temp_b2_3_5_r;
wire signed [`CalcTempBus]          temp_b2_3_5_i;
wire signed [`CalcTempBus]          temp_b2_3_6_r;
wire signed [`CalcTempBus]          temp_b2_3_6_i;
wire signed [`CalcTempBus]          temp_b2_3_7_r;
wire signed [`CalcTempBus]          temp_b2_3_7_i;
wire signed [`CalcTempBus]          temp_b2_3_8_r;
wire signed [`CalcTempBus]          temp_b2_3_8_i;
wire signed [`CalcTempBus]          temp_b2_3_9_r;
wire signed [`CalcTempBus]          temp_b2_3_9_i;
wire signed [`CalcTempBus]          temp_b2_3_10_r;
wire signed [`CalcTempBus]          temp_b2_3_10_i;
wire signed [`CalcTempBus]          temp_b2_3_11_r;
wire signed [`CalcTempBus]          temp_b2_3_11_i;
wire signed [`CalcTempBus]          temp_b2_3_12_r;
wire signed [`CalcTempBus]          temp_b2_3_12_i;
wire signed [`CalcTempBus]          temp_b2_3_13_r;
wire signed [`CalcTempBus]          temp_b2_3_13_i;
wire signed [`CalcTempBus]          temp_b2_3_14_r;
wire signed [`CalcTempBus]          temp_b2_3_14_i;
wire signed [`CalcTempBus]          temp_b2_3_15_r;
wire signed [`CalcTempBus]          temp_b2_3_15_i;
wire signed [`CalcTempBus]          temp_b2_3_16_r;
wire signed [`CalcTempBus]          temp_b2_3_16_i;
wire signed [`CalcTempBus]          temp_b2_4_1_r;
wire signed [`CalcTempBus]          temp_b2_4_1_i;
wire signed [`CalcTempBus]          temp_b2_4_2_r;
wire signed [`CalcTempBus]          temp_b2_4_2_i;
wire signed [`CalcTempBus]          temp_b2_4_3_r;
wire signed [`CalcTempBus]          temp_b2_4_3_i;
wire signed [`CalcTempBus]          temp_b2_4_4_r;
wire signed [`CalcTempBus]          temp_b2_4_4_i;
wire signed [`CalcTempBus]          temp_b2_4_5_r;
wire signed [`CalcTempBus]          temp_b2_4_5_i;
wire signed [`CalcTempBus]          temp_b2_4_6_r;
wire signed [`CalcTempBus]          temp_b2_4_6_i;
wire signed [`CalcTempBus]          temp_b2_4_7_r;
wire signed [`CalcTempBus]          temp_b2_4_7_i;
wire signed [`CalcTempBus]          temp_b2_4_8_r;
wire signed [`CalcTempBus]          temp_b2_4_8_i;
wire signed [`CalcTempBus]          temp_b2_4_9_r;
wire signed [`CalcTempBus]          temp_b2_4_9_i;
wire signed [`CalcTempBus]          temp_b2_4_10_r;
wire signed [`CalcTempBus]          temp_b2_4_10_i;
wire signed [`CalcTempBus]          temp_b2_4_11_r;
wire signed [`CalcTempBus]          temp_b2_4_11_i;
wire signed [`CalcTempBus]          temp_b2_4_12_r;
wire signed [`CalcTempBus]          temp_b2_4_12_i;
wire signed [`CalcTempBus]          temp_b2_4_13_r;
wire signed [`CalcTempBus]          temp_b2_4_13_i;
wire signed [`CalcTempBus]          temp_b2_4_14_r;
wire signed [`CalcTempBus]          temp_b2_4_14_i;
wire signed [`CalcTempBus]          temp_b2_4_15_r;
wire signed [`CalcTempBus]          temp_b2_4_15_i;
wire signed [`CalcTempBus]          temp_b2_4_16_r;
wire signed [`CalcTempBus]          temp_b2_4_16_i;
wire signed [`CalcTempBus]          temp_b2_5_1_r;
wire signed [`CalcTempBus]          temp_b2_5_1_i;
wire signed [`CalcTempBus]          temp_b2_5_2_r;
wire signed [`CalcTempBus]          temp_b2_5_2_i;
wire signed [`CalcTempBus]          temp_b2_5_3_r;
wire signed [`CalcTempBus]          temp_b2_5_3_i;
wire signed [`CalcTempBus]          temp_b2_5_4_r;
wire signed [`CalcTempBus]          temp_b2_5_4_i;
wire signed [`CalcTempBus]          temp_b2_5_5_r;
wire signed [`CalcTempBus]          temp_b2_5_5_i;
wire signed [`CalcTempBus]          temp_b2_5_6_r;
wire signed [`CalcTempBus]          temp_b2_5_6_i;
wire signed [`CalcTempBus]          temp_b2_5_7_r;
wire signed [`CalcTempBus]          temp_b2_5_7_i;
wire signed [`CalcTempBus]          temp_b2_5_8_r;
wire signed [`CalcTempBus]          temp_b2_5_8_i;
wire signed [`CalcTempBus]          temp_b2_5_9_r;
wire signed [`CalcTempBus]          temp_b2_5_9_i;
wire signed [`CalcTempBus]          temp_b2_5_10_r;
wire signed [`CalcTempBus]          temp_b2_5_10_i;
wire signed [`CalcTempBus]          temp_b2_5_11_r;
wire signed [`CalcTempBus]          temp_b2_5_11_i;
wire signed [`CalcTempBus]          temp_b2_5_12_r;
wire signed [`CalcTempBus]          temp_b2_5_12_i;
wire signed [`CalcTempBus]          temp_b2_5_13_r;
wire signed [`CalcTempBus]          temp_b2_5_13_i;
wire signed [`CalcTempBus]          temp_b2_5_14_r;
wire signed [`CalcTempBus]          temp_b2_5_14_i;
wire signed [`CalcTempBus]          temp_b2_5_15_r;
wire signed [`CalcTempBus]          temp_b2_5_15_i;
wire signed [`CalcTempBus]          temp_b2_5_16_r;
wire signed [`CalcTempBus]          temp_b2_5_16_i;
wire signed [`CalcTempBus]          temp_b2_6_1_r;
wire signed [`CalcTempBus]          temp_b2_6_1_i;
wire signed [`CalcTempBus]          temp_b2_6_2_r;
wire signed [`CalcTempBus]          temp_b2_6_2_i;
wire signed [`CalcTempBus]          temp_b2_6_3_r;
wire signed [`CalcTempBus]          temp_b2_6_3_i;
wire signed [`CalcTempBus]          temp_b2_6_4_r;
wire signed [`CalcTempBus]          temp_b2_6_4_i;
wire signed [`CalcTempBus]          temp_b2_6_5_r;
wire signed [`CalcTempBus]          temp_b2_6_5_i;
wire signed [`CalcTempBus]          temp_b2_6_6_r;
wire signed [`CalcTempBus]          temp_b2_6_6_i;
wire signed [`CalcTempBus]          temp_b2_6_7_r;
wire signed [`CalcTempBus]          temp_b2_6_7_i;
wire signed [`CalcTempBus]          temp_b2_6_8_r;
wire signed [`CalcTempBus]          temp_b2_6_8_i;
wire signed [`CalcTempBus]          temp_b2_6_9_r;
wire signed [`CalcTempBus]          temp_b2_6_9_i;
wire signed [`CalcTempBus]          temp_b2_6_10_r;
wire signed [`CalcTempBus]          temp_b2_6_10_i;
wire signed [`CalcTempBus]          temp_b2_6_11_r;
wire signed [`CalcTempBus]          temp_b2_6_11_i;
wire signed [`CalcTempBus]          temp_b2_6_12_r;
wire signed [`CalcTempBus]          temp_b2_6_12_i;
wire signed [`CalcTempBus]          temp_b2_6_13_r;
wire signed [`CalcTempBus]          temp_b2_6_13_i;
wire signed [`CalcTempBus]          temp_b2_6_14_r;
wire signed [`CalcTempBus]          temp_b2_6_14_i;
wire signed [`CalcTempBus]          temp_b2_6_15_r;
wire signed [`CalcTempBus]          temp_b2_6_15_i;
wire signed [`CalcTempBus]          temp_b2_6_16_r;
wire signed [`CalcTempBus]          temp_b2_6_16_i;
wire signed [`CalcTempBus]          temp_b2_7_1_r;
wire signed [`CalcTempBus]          temp_b2_7_1_i;
wire signed [`CalcTempBus]          temp_b2_7_2_r;
wire signed [`CalcTempBus]          temp_b2_7_2_i;
wire signed [`CalcTempBus]          temp_b2_7_3_r;
wire signed [`CalcTempBus]          temp_b2_7_3_i;
wire signed [`CalcTempBus]          temp_b2_7_4_r;
wire signed [`CalcTempBus]          temp_b2_7_4_i;
wire signed [`CalcTempBus]          temp_b2_7_5_r;
wire signed [`CalcTempBus]          temp_b2_7_5_i;
wire signed [`CalcTempBus]          temp_b2_7_6_r;
wire signed [`CalcTempBus]          temp_b2_7_6_i;
wire signed [`CalcTempBus]          temp_b2_7_7_r;
wire signed [`CalcTempBus]          temp_b2_7_7_i;
wire signed [`CalcTempBus]          temp_b2_7_8_r;
wire signed [`CalcTempBus]          temp_b2_7_8_i;
wire signed [`CalcTempBus]          temp_b2_7_9_r;
wire signed [`CalcTempBus]          temp_b2_7_9_i;
wire signed [`CalcTempBus]          temp_b2_7_10_r;
wire signed [`CalcTempBus]          temp_b2_7_10_i;
wire signed [`CalcTempBus]          temp_b2_7_11_r;
wire signed [`CalcTempBus]          temp_b2_7_11_i;
wire signed [`CalcTempBus]          temp_b2_7_12_r;
wire signed [`CalcTempBus]          temp_b2_7_12_i;
wire signed [`CalcTempBus]          temp_b2_7_13_r;
wire signed [`CalcTempBus]          temp_b2_7_13_i;
wire signed [`CalcTempBus]          temp_b2_7_14_r;
wire signed [`CalcTempBus]          temp_b2_7_14_i;
wire signed [`CalcTempBus]          temp_b2_7_15_r;
wire signed [`CalcTempBus]          temp_b2_7_15_i;
wire signed [`CalcTempBus]          temp_b2_7_16_r;
wire signed [`CalcTempBus]          temp_b2_7_16_i;
wire signed [`CalcTempBus]          temp_b2_8_1_r;
wire signed [`CalcTempBus]          temp_b2_8_1_i;
wire signed [`CalcTempBus]          temp_b2_8_2_r;
wire signed [`CalcTempBus]          temp_b2_8_2_i;
wire signed [`CalcTempBus]          temp_b2_8_3_r;
wire signed [`CalcTempBus]          temp_b2_8_3_i;
wire signed [`CalcTempBus]          temp_b2_8_4_r;
wire signed [`CalcTempBus]          temp_b2_8_4_i;
wire signed [`CalcTempBus]          temp_b2_8_5_r;
wire signed [`CalcTempBus]          temp_b2_8_5_i;
wire signed [`CalcTempBus]          temp_b2_8_6_r;
wire signed [`CalcTempBus]          temp_b2_8_6_i;
wire signed [`CalcTempBus]          temp_b2_8_7_r;
wire signed [`CalcTempBus]          temp_b2_8_7_i;
wire signed [`CalcTempBus]          temp_b2_8_8_r;
wire signed [`CalcTempBus]          temp_b2_8_8_i;
wire signed [`CalcTempBus]          temp_b2_8_9_r;
wire signed [`CalcTempBus]          temp_b2_8_9_i;
wire signed [`CalcTempBus]          temp_b2_8_10_r;
wire signed [`CalcTempBus]          temp_b2_8_10_i;
wire signed [`CalcTempBus]          temp_b2_8_11_r;
wire signed [`CalcTempBus]          temp_b2_8_11_i;
wire signed [`CalcTempBus]          temp_b2_8_12_r;
wire signed [`CalcTempBus]          temp_b2_8_12_i;
wire signed [`CalcTempBus]          temp_b2_8_13_r;
wire signed [`CalcTempBus]          temp_b2_8_13_i;
wire signed [`CalcTempBus]          temp_b2_8_14_r;
wire signed [`CalcTempBus]          temp_b2_8_14_i;
wire signed [`CalcTempBus]          temp_b2_8_15_r;
wire signed [`CalcTempBus]          temp_b2_8_15_i;
wire signed [`CalcTempBus]          temp_b2_8_16_r;
wire signed [`CalcTempBus]          temp_b2_8_16_i;
wire signed [`CalcTempBus]          temp_b2_9_1_r;
wire signed [`CalcTempBus]          temp_b2_9_1_i;
wire signed [`CalcTempBus]          temp_b2_9_2_r;
wire signed [`CalcTempBus]          temp_b2_9_2_i;
wire signed [`CalcTempBus]          temp_b2_9_3_r;
wire signed [`CalcTempBus]          temp_b2_9_3_i;
wire signed [`CalcTempBus]          temp_b2_9_4_r;
wire signed [`CalcTempBus]          temp_b2_9_4_i;
wire signed [`CalcTempBus]          temp_b2_9_5_r;
wire signed [`CalcTempBus]          temp_b2_9_5_i;
wire signed [`CalcTempBus]          temp_b2_9_6_r;
wire signed [`CalcTempBus]          temp_b2_9_6_i;
wire signed [`CalcTempBus]          temp_b2_9_7_r;
wire signed [`CalcTempBus]          temp_b2_9_7_i;
wire signed [`CalcTempBus]          temp_b2_9_8_r;
wire signed [`CalcTempBus]          temp_b2_9_8_i;
wire signed [`CalcTempBus]          temp_b2_9_9_r;
wire signed [`CalcTempBus]          temp_b2_9_9_i;
wire signed [`CalcTempBus]          temp_b2_9_10_r;
wire signed [`CalcTempBus]          temp_b2_9_10_i;
wire signed [`CalcTempBus]          temp_b2_9_11_r;
wire signed [`CalcTempBus]          temp_b2_9_11_i;
wire signed [`CalcTempBus]          temp_b2_9_12_r;
wire signed [`CalcTempBus]          temp_b2_9_12_i;
wire signed [`CalcTempBus]          temp_b2_9_13_r;
wire signed [`CalcTempBus]          temp_b2_9_13_i;
wire signed [`CalcTempBus]          temp_b2_9_14_r;
wire signed [`CalcTempBus]          temp_b2_9_14_i;
wire signed [`CalcTempBus]          temp_b2_9_15_r;
wire signed [`CalcTempBus]          temp_b2_9_15_i;
wire signed [`CalcTempBus]          temp_b2_9_16_r;
wire signed [`CalcTempBus]          temp_b2_9_16_i;
wire signed [`CalcTempBus]          temp_b2_10_1_r;
wire signed [`CalcTempBus]          temp_b2_10_1_i;
wire signed [`CalcTempBus]          temp_b2_10_2_r;
wire signed [`CalcTempBus]          temp_b2_10_2_i;
wire signed [`CalcTempBus]          temp_b2_10_3_r;
wire signed [`CalcTempBus]          temp_b2_10_3_i;
wire signed [`CalcTempBus]          temp_b2_10_4_r;
wire signed [`CalcTempBus]          temp_b2_10_4_i;
wire signed [`CalcTempBus]          temp_b2_10_5_r;
wire signed [`CalcTempBus]          temp_b2_10_5_i;
wire signed [`CalcTempBus]          temp_b2_10_6_r;
wire signed [`CalcTempBus]          temp_b2_10_6_i;
wire signed [`CalcTempBus]          temp_b2_10_7_r;
wire signed [`CalcTempBus]          temp_b2_10_7_i;
wire signed [`CalcTempBus]          temp_b2_10_8_r;
wire signed [`CalcTempBus]          temp_b2_10_8_i;
wire signed [`CalcTempBus]          temp_b2_10_9_r;
wire signed [`CalcTempBus]          temp_b2_10_9_i;
wire signed [`CalcTempBus]          temp_b2_10_10_r;
wire signed [`CalcTempBus]          temp_b2_10_10_i;
wire signed [`CalcTempBus]          temp_b2_10_11_r;
wire signed [`CalcTempBus]          temp_b2_10_11_i;
wire signed [`CalcTempBus]          temp_b2_10_12_r;
wire signed [`CalcTempBus]          temp_b2_10_12_i;
wire signed [`CalcTempBus]          temp_b2_10_13_r;
wire signed [`CalcTempBus]          temp_b2_10_13_i;
wire signed [`CalcTempBus]          temp_b2_10_14_r;
wire signed [`CalcTempBus]          temp_b2_10_14_i;
wire signed [`CalcTempBus]          temp_b2_10_15_r;
wire signed [`CalcTempBus]          temp_b2_10_15_i;
wire signed [`CalcTempBus]          temp_b2_10_16_r;
wire signed [`CalcTempBus]          temp_b2_10_16_i;
wire signed [`CalcTempBus]          temp_b2_11_1_r;
wire signed [`CalcTempBus]          temp_b2_11_1_i;
wire signed [`CalcTempBus]          temp_b2_11_2_r;
wire signed [`CalcTempBus]          temp_b2_11_2_i;
wire signed [`CalcTempBus]          temp_b2_11_3_r;
wire signed [`CalcTempBus]          temp_b2_11_3_i;
wire signed [`CalcTempBus]          temp_b2_11_4_r;
wire signed [`CalcTempBus]          temp_b2_11_4_i;
wire signed [`CalcTempBus]          temp_b2_11_5_r;
wire signed [`CalcTempBus]          temp_b2_11_5_i;
wire signed [`CalcTempBus]          temp_b2_11_6_r;
wire signed [`CalcTempBus]          temp_b2_11_6_i;
wire signed [`CalcTempBus]          temp_b2_11_7_r;
wire signed [`CalcTempBus]          temp_b2_11_7_i;
wire signed [`CalcTempBus]          temp_b2_11_8_r;
wire signed [`CalcTempBus]          temp_b2_11_8_i;
wire signed [`CalcTempBus]          temp_b2_11_9_r;
wire signed [`CalcTempBus]          temp_b2_11_9_i;
wire signed [`CalcTempBus]          temp_b2_11_10_r;
wire signed [`CalcTempBus]          temp_b2_11_10_i;
wire signed [`CalcTempBus]          temp_b2_11_11_r;
wire signed [`CalcTempBus]          temp_b2_11_11_i;
wire signed [`CalcTempBus]          temp_b2_11_12_r;
wire signed [`CalcTempBus]          temp_b2_11_12_i;
wire signed [`CalcTempBus]          temp_b2_11_13_r;
wire signed [`CalcTempBus]          temp_b2_11_13_i;
wire signed [`CalcTempBus]          temp_b2_11_14_r;
wire signed [`CalcTempBus]          temp_b2_11_14_i;
wire signed [`CalcTempBus]          temp_b2_11_15_r;
wire signed [`CalcTempBus]          temp_b2_11_15_i;
wire signed [`CalcTempBus]          temp_b2_11_16_r;
wire signed [`CalcTempBus]          temp_b2_11_16_i;
wire signed [`CalcTempBus]          temp_b2_12_1_r;
wire signed [`CalcTempBus]          temp_b2_12_1_i;
wire signed [`CalcTempBus]          temp_b2_12_2_r;
wire signed [`CalcTempBus]          temp_b2_12_2_i;
wire signed [`CalcTempBus]          temp_b2_12_3_r;
wire signed [`CalcTempBus]          temp_b2_12_3_i;
wire signed [`CalcTempBus]          temp_b2_12_4_r;
wire signed [`CalcTempBus]          temp_b2_12_4_i;
wire signed [`CalcTempBus]          temp_b2_12_5_r;
wire signed [`CalcTempBus]          temp_b2_12_5_i;
wire signed [`CalcTempBus]          temp_b2_12_6_r;
wire signed [`CalcTempBus]          temp_b2_12_6_i;
wire signed [`CalcTempBus]          temp_b2_12_7_r;
wire signed [`CalcTempBus]          temp_b2_12_7_i;
wire signed [`CalcTempBus]          temp_b2_12_8_r;
wire signed [`CalcTempBus]          temp_b2_12_8_i;
wire signed [`CalcTempBus]          temp_b2_12_9_r;
wire signed [`CalcTempBus]          temp_b2_12_9_i;
wire signed [`CalcTempBus]          temp_b2_12_10_r;
wire signed [`CalcTempBus]          temp_b2_12_10_i;
wire signed [`CalcTempBus]          temp_b2_12_11_r;
wire signed [`CalcTempBus]          temp_b2_12_11_i;
wire signed [`CalcTempBus]          temp_b2_12_12_r;
wire signed [`CalcTempBus]          temp_b2_12_12_i;
wire signed [`CalcTempBus]          temp_b2_12_13_r;
wire signed [`CalcTempBus]          temp_b2_12_13_i;
wire signed [`CalcTempBus]          temp_b2_12_14_r;
wire signed [`CalcTempBus]          temp_b2_12_14_i;
wire signed [`CalcTempBus]          temp_b2_12_15_r;
wire signed [`CalcTempBus]          temp_b2_12_15_i;
wire signed [`CalcTempBus]          temp_b2_12_16_r;
wire signed [`CalcTempBus]          temp_b2_12_16_i;
wire signed [`CalcTempBus]          temp_b2_13_1_r;
wire signed [`CalcTempBus]          temp_b2_13_1_i;
wire signed [`CalcTempBus]          temp_b2_13_2_r;
wire signed [`CalcTempBus]          temp_b2_13_2_i;
wire signed [`CalcTempBus]          temp_b2_13_3_r;
wire signed [`CalcTempBus]          temp_b2_13_3_i;
wire signed [`CalcTempBus]          temp_b2_13_4_r;
wire signed [`CalcTempBus]          temp_b2_13_4_i;
wire signed [`CalcTempBus]          temp_b2_13_5_r;
wire signed [`CalcTempBus]          temp_b2_13_5_i;
wire signed [`CalcTempBus]          temp_b2_13_6_r;
wire signed [`CalcTempBus]          temp_b2_13_6_i;
wire signed [`CalcTempBus]          temp_b2_13_7_r;
wire signed [`CalcTempBus]          temp_b2_13_7_i;
wire signed [`CalcTempBus]          temp_b2_13_8_r;
wire signed [`CalcTempBus]          temp_b2_13_8_i;
wire signed [`CalcTempBus]          temp_b2_13_9_r;
wire signed [`CalcTempBus]          temp_b2_13_9_i;
wire signed [`CalcTempBus]          temp_b2_13_10_r;
wire signed [`CalcTempBus]          temp_b2_13_10_i;
wire signed [`CalcTempBus]          temp_b2_13_11_r;
wire signed [`CalcTempBus]          temp_b2_13_11_i;
wire signed [`CalcTempBus]          temp_b2_13_12_r;
wire signed [`CalcTempBus]          temp_b2_13_12_i;
wire signed [`CalcTempBus]          temp_b2_13_13_r;
wire signed [`CalcTempBus]          temp_b2_13_13_i;
wire signed [`CalcTempBus]          temp_b2_13_14_r;
wire signed [`CalcTempBus]          temp_b2_13_14_i;
wire signed [`CalcTempBus]          temp_b2_13_15_r;
wire signed [`CalcTempBus]          temp_b2_13_15_i;
wire signed [`CalcTempBus]          temp_b2_13_16_r;
wire signed [`CalcTempBus]          temp_b2_13_16_i;
wire signed [`CalcTempBus]          temp_b2_14_1_r;
wire signed [`CalcTempBus]          temp_b2_14_1_i;
wire signed [`CalcTempBus]          temp_b2_14_2_r;
wire signed [`CalcTempBus]          temp_b2_14_2_i;
wire signed [`CalcTempBus]          temp_b2_14_3_r;
wire signed [`CalcTempBus]          temp_b2_14_3_i;
wire signed [`CalcTempBus]          temp_b2_14_4_r;
wire signed [`CalcTempBus]          temp_b2_14_4_i;
wire signed [`CalcTempBus]          temp_b2_14_5_r;
wire signed [`CalcTempBus]          temp_b2_14_5_i;
wire signed [`CalcTempBus]          temp_b2_14_6_r;
wire signed [`CalcTempBus]          temp_b2_14_6_i;
wire signed [`CalcTempBus]          temp_b2_14_7_r;
wire signed [`CalcTempBus]          temp_b2_14_7_i;
wire signed [`CalcTempBus]          temp_b2_14_8_r;
wire signed [`CalcTempBus]          temp_b2_14_8_i;
wire signed [`CalcTempBus]          temp_b2_14_9_r;
wire signed [`CalcTempBus]          temp_b2_14_9_i;
wire signed [`CalcTempBus]          temp_b2_14_10_r;
wire signed [`CalcTempBus]          temp_b2_14_10_i;
wire signed [`CalcTempBus]          temp_b2_14_11_r;
wire signed [`CalcTempBus]          temp_b2_14_11_i;
wire signed [`CalcTempBus]          temp_b2_14_12_r;
wire signed [`CalcTempBus]          temp_b2_14_12_i;
wire signed [`CalcTempBus]          temp_b2_14_13_r;
wire signed [`CalcTempBus]          temp_b2_14_13_i;
wire signed [`CalcTempBus]          temp_b2_14_14_r;
wire signed [`CalcTempBus]          temp_b2_14_14_i;
wire signed [`CalcTempBus]          temp_b2_14_15_r;
wire signed [`CalcTempBus]          temp_b2_14_15_i;
wire signed [`CalcTempBus]          temp_b2_14_16_r;
wire signed [`CalcTempBus]          temp_b2_14_16_i;
wire signed [`CalcTempBus]          temp_b2_15_1_r;
wire signed [`CalcTempBus]          temp_b2_15_1_i;
wire signed [`CalcTempBus]          temp_b2_15_2_r;
wire signed [`CalcTempBus]          temp_b2_15_2_i;
wire signed [`CalcTempBus]          temp_b2_15_3_r;
wire signed [`CalcTempBus]          temp_b2_15_3_i;
wire signed [`CalcTempBus]          temp_b2_15_4_r;
wire signed [`CalcTempBus]          temp_b2_15_4_i;
wire signed [`CalcTempBus]          temp_b2_15_5_r;
wire signed [`CalcTempBus]          temp_b2_15_5_i;
wire signed [`CalcTempBus]          temp_b2_15_6_r;
wire signed [`CalcTempBus]          temp_b2_15_6_i;
wire signed [`CalcTempBus]          temp_b2_15_7_r;
wire signed [`CalcTempBus]          temp_b2_15_7_i;
wire signed [`CalcTempBus]          temp_b2_15_8_r;
wire signed [`CalcTempBus]          temp_b2_15_8_i;
wire signed [`CalcTempBus]          temp_b2_15_9_r;
wire signed [`CalcTempBus]          temp_b2_15_9_i;
wire signed [`CalcTempBus]          temp_b2_15_10_r;
wire signed [`CalcTempBus]          temp_b2_15_10_i;
wire signed [`CalcTempBus]          temp_b2_15_11_r;
wire signed [`CalcTempBus]          temp_b2_15_11_i;
wire signed [`CalcTempBus]          temp_b2_15_12_r;
wire signed [`CalcTempBus]          temp_b2_15_12_i;
wire signed [`CalcTempBus]          temp_b2_15_13_r;
wire signed [`CalcTempBus]          temp_b2_15_13_i;
wire signed [`CalcTempBus]          temp_b2_15_14_r;
wire signed [`CalcTempBus]          temp_b2_15_14_i;
wire signed [`CalcTempBus]          temp_b2_15_15_r;
wire signed [`CalcTempBus]          temp_b2_15_15_i;
wire signed [`CalcTempBus]          temp_b2_15_16_r;
wire signed [`CalcTempBus]          temp_b2_15_16_i;
wire signed [`CalcTempBus]          temp_b2_16_1_r;
wire signed [`CalcTempBus]          temp_b2_16_1_i;
wire signed [`CalcTempBus]          temp_b2_16_2_r;
wire signed [`CalcTempBus]          temp_b2_16_2_i;
wire signed [`CalcTempBus]          temp_b2_16_3_r;
wire signed [`CalcTempBus]          temp_b2_16_3_i;
wire signed [`CalcTempBus]          temp_b2_16_4_r;
wire signed [`CalcTempBus]          temp_b2_16_4_i;
wire signed [`CalcTempBus]          temp_b2_16_5_r;
wire signed [`CalcTempBus]          temp_b2_16_5_i;
wire signed [`CalcTempBus]          temp_b2_16_6_r;
wire signed [`CalcTempBus]          temp_b2_16_6_i;
wire signed [`CalcTempBus]          temp_b2_16_7_r;
wire signed [`CalcTempBus]          temp_b2_16_7_i;
wire signed [`CalcTempBus]          temp_b2_16_8_r;
wire signed [`CalcTempBus]          temp_b2_16_8_i;
wire signed [`CalcTempBus]          temp_b2_16_9_r;
wire signed [`CalcTempBus]          temp_b2_16_9_i;
wire signed [`CalcTempBus]          temp_b2_16_10_r;
wire signed [`CalcTempBus]          temp_b2_16_10_i;
wire signed [`CalcTempBus]          temp_b2_16_11_r;
wire signed [`CalcTempBus]          temp_b2_16_11_i;
wire signed [`CalcTempBus]          temp_b2_16_12_r;
wire signed [`CalcTempBus]          temp_b2_16_12_i;
wire signed [`CalcTempBus]          temp_b2_16_13_r;
wire signed [`CalcTempBus]          temp_b2_16_13_i;
wire signed [`CalcTempBus]          temp_b2_16_14_r;
wire signed [`CalcTempBus]          temp_b2_16_14_i;
wire signed [`CalcTempBus]          temp_b2_16_15_r;
wire signed [`CalcTempBus]          temp_b2_16_15_i;
wire signed [`CalcTempBus]          temp_b2_16_16_r;
wire signed [`CalcTempBus]          temp_b2_16_16_i;
wire signed [`CalcTempBus]          temp_b3_1_1_r;
wire signed [`CalcTempBus]          temp_b3_1_1_i;
wire signed [`CalcTempBus]          temp_b3_1_2_r;
wire signed [`CalcTempBus]          temp_b3_1_2_i;
wire signed [`CalcTempBus]          temp_b3_1_3_r;
wire signed [`CalcTempBus]          temp_b3_1_3_i;
wire signed [`CalcTempBus]          temp_b3_1_4_r;
wire signed [`CalcTempBus]          temp_b3_1_4_i;
wire signed [`CalcTempBus]          temp_b3_1_5_r;
wire signed [`CalcTempBus]          temp_b3_1_5_i;
wire signed [`CalcTempBus]          temp_b3_1_6_r;
wire signed [`CalcTempBus]          temp_b3_1_6_i;
wire signed [`CalcTempBus]          temp_b3_1_7_r;
wire signed [`CalcTempBus]          temp_b3_1_7_i;
wire signed [`CalcTempBus]          temp_b3_1_8_r;
wire signed [`CalcTempBus]          temp_b3_1_8_i;
wire signed [`CalcTempBus]          temp_b3_1_9_r;
wire signed [`CalcTempBus]          temp_b3_1_9_i;
wire signed [`CalcTempBus]          temp_b3_1_10_r;
wire signed [`CalcTempBus]          temp_b3_1_10_i;
wire signed [`CalcTempBus]          temp_b3_1_11_r;
wire signed [`CalcTempBus]          temp_b3_1_11_i;
wire signed [`CalcTempBus]          temp_b3_1_12_r;
wire signed [`CalcTempBus]          temp_b3_1_12_i;
wire signed [`CalcTempBus]          temp_b3_1_13_r;
wire signed [`CalcTempBus]          temp_b3_1_13_i;
wire signed [`CalcTempBus]          temp_b3_1_14_r;
wire signed [`CalcTempBus]          temp_b3_1_14_i;
wire signed [`CalcTempBus]          temp_b3_1_15_r;
wire signed [`CalcTempBus]          temp_b3_1_15_i;
wire signed [`CalcTempBus]          temp_b3_1_16_r;
wire signed [`CalcTempBus]          temp_b3_1_16_i;
wire signed [`CalcTempBus]          temp_b3_2_1_r;
wire signed [`CalcTempBus]          temp_b3_2_1_i;
wire signed [`CalcTempBus]          temp_b3_2_2_r;
wire signed [`CalcTempBus]          temp_b3_2_2_i;
wire signed [`CalcTempBus]          temp_b3_2_3_r;
wire signed [`CalcTempBus]          temp_b3_2_3_i;
wire signed [`CalcTempBus]          temp_b3_2_4_r;
wire signed [`CalcTempBus]          temp_b3_2_4_i;
wire signed [`CalcTempBus]          temp_b3_2_5_r;
wire signed [`CalcTempBus]          temp_b3_2_5_i;
wire signed [`CalcTempBus]          temp_b3_2_6_r;
wire signed [`CalcTempBus]          temp_b3_2_6_i;
wire signed [`CalcTempBus]          temp_b3_2_7_r;
wire signed [`CalcTempBus]          temp_b3_2_7_i;
wire signed [`CalcTempBus]          temp_b3_2_8_r;
wire signed [`CalcTempBus]          temp_b3_2_8_i;
wire signed [`CalcTempBus]          temp_b3_2_9_r;
wire signed [`CalcTempBus]          temp_b3_2_9_i;
wire signed [`CalcTempBus]          temp_b3_2_10_r;
wire signed [`CalcTempBus]          temp_b3_2_10_i;
wire signed [`CalcTempBus]          temp_b3_2_11_r;
wire signed [`CalcTempBus]          temp_b3_2_11_i;
wire signed [`CalcTempBus]          temp_b3_2_12_r;
wire signed [`CalcTempBus]          temp_b3_2_12_i;
wire signed [`CalcTempBus]          temp_b3_2_13_r;
wire signed [`CalcTempBus]          temp_b3_2_13_i;
wire signed [`CalcTempBus]          temp_b3_2_14_r;
wire signed [`CalcTempBus]          temp_b3_2_14_i;
wire signed [`CalcTempBus]          temp_b3_2_15_r;
wire signed [`CalcTempBus]          temp_b3_2_15_i;
wire signed [`CalcTempBus]          temp_b3_2_16_r;
wire signed [`CalcTempBus]          temp_b3_2_16_i;
wire signed [`CalcTempBus]          temp_b3_3_1_r;
wire signed [`CalcTempBus]          temp_b3_3_1_i;
wire signed [`CalcTempBus]          temp_b3_3_2_r;
wire signed [`CalcTempBus]          temp_b3_3_2_i;
wire signed [`CalcTempBus]          temp_b3_3_3_r;
wire signed [`CalcTempBus]          temp_b3_3_3_i;
wire signed [`CalcTempBus]          temp_b3_3_4_r;
wire signed [`CalcTempBus]          temp_b3_3_4_i;
wire signed [`CalcTempBus]          temp_b3_3_5_r;
wire signed [`CalcTempBus]          temp_b3_3_5_i;
wire signed [`CalcTempBus]          temp_b3_3_6_r;
wire signed [`CalcTempBus]          temp_b3_3_6_i;
wire signed [`CalcTempBus]          temp_b3_3_7_r;
wire signed [`CalcTempBus]          temp_b3_3_7_i;
wire signed [`CalcTempBus]          temp_b3_3_8_r;
wire signed [`CalcTempBus]          temp_b3_3_8_i;
wire signed [`CalcTempBus]          temp_b3_3_9_r;
wire signed [`CalcTempBus]          temp_b3_3_9_i;
wire signed [`CalcTempBus]          temp_b3_3_10_r;
wire signed [`CalcTempBus]          temp_b3_3_10_i;
wire signed [`CalcTempBus]          temp_b3_3_11_r;
wire signed [`CalcTempBus]          temp_b3_3_11_i;
wire signed [`CalcTempBus]          temp_b3_3_12_r;
wire signed [`CalcTempBus]          temp_b3_3_12_i;
wire signed [`CalcTempBus]          temp_b3_3_13_r;
wire signed [`CalcTempBus]          temp_b3_3_13_i;
wire signed [`CalcTempBus]          temp_b3_3_14_r;
wire signed [`CalcTempBus]          temp_b3_3_14_i;
wire signed [`CalcTempBus]          temp_b3_3_15_r;
wire signed [`CalcTempBus]          temp_b3_3_15_i;
wire signed [`CalcTempBus]          temp_b3_3_16_r;
wire signed [`CalcTempBus]          temp_b3_3_16_i;
wire signed [`CalcTempBus]          temp_b3_4_1_r;
wire signed [`CalcTempBus]          temp_b3_4_1_i;
wire signed [`CalcTempBus]          temp_b3_4_2_r;
wire signed [`CalcTempBus]          temp_b3_4_2_i;
wire signed [`CalcTempBus]          temp_b3_4_3_r;
wire signed [`CalcTempBus]          temp_b3_4_3_i;
wire signed [`CalcTempBus]          temp_b3_4_4_r;
wire signed [`CalcTempBus]          temp_b3_4_4_i;
wire signed [`CalcTempBus]          temp_b3_4_5_r;
wire signed [`CalcTempBus]          temp_b3_4_5_i;
wire signed [`CalcTempBus]          temp_b3_4_6_r;
wire signed [`CalcTempBus]          temp_b3_4_6_i;
wire signed [`CalcTempBus]          temp_b3_4_7_r;
wire signed [`CalcTempBus]          temp_b3_4_7_i;
wire signed [`CalcTempBus]          temp_b3_4_8_r;
wire signed [`CalcTempBus]          temp_b3_4_8_i;
wire signed [`CalcTempBus]          temp_b3_4_9_r;
wire signed [`CalcTempBus]          temp_b3_4_9_i;
wire signed [`CalcTempBus]          temp_b3_4_10_r;
wire signed [`CalcTempBus]          temp_b3_4_10_i;
wire signed [`CalcTempBus]          temp_b3_4_11_r;
wire signed [`CalcTempBus]          temp_b3_4_11_i;
wire signed [`CalcTempBus]          temp_b3_4_12_r;
wire signed [`CalcTempBus]          temp_b3_4_12_i;
wire signed [`CalcTempBus]          temp_b3_4_13_r;
wire signed [`CalcTempBus]          temp_b3_4_13_i;
wire signed [`CalcTempBus]          temp_b3_4_14_r;
wire signed [`CalcTempBus]          temp_b3_4_14_i;
wire signed [`CalcTempBus]          temp_b3_4_15_r;
wire signed [`CalcTempBus]          temp_b3_4_15_i;
wire signed [`CalcTempBus]          temp_b3_4_16_r;
wire signed [`CalcTempBus]          temp_b3_4_16_i;
wire signed [`CalcTempBus]          temp_b3_5_1_r;
wire signed [`CalcTempBus]          temp_b3_5_1_i;
wire signed [`CalcTempBus]          temp_b3_5_2_r;
wire signed [`CalcTempBus]          temp_b3_5_2_i;
wire signed [`CalcTempBus]          temp_b3_5_3_r;
wire signed [`CalcTempBus]          temp_b3_5_3_i;
wire signed [`CalcTempBus]          temp_b3_5_4_r;
wire signed [`CalcTempBus]          temp_b3_5_4_i;
wire signed [`CalcTempBus]          temp_b3_5_5_r;
wire signed [`CalcTempBus]          temp_b3_5_5_i;
wire signed [`CalcTempBus]          temp_b3_5_6_r;
wire signed [`CalcTempBus]          temp_b3_5_6_i;
wire signed [`CalcTempBus]          temp_b3_5_7_r;
wire signed [`CalcTempBus]          temp_b3_5_7_i;
wire signed [`CalcTempBus]          temp_b3_5_8_r;
wire signed [`CalcTempBus]          temp_b3_5_8_i;
wire signed [`CalcTempBus]          temp_b3_5_9_r;
wire signed [`CalcTempBus]          temp_b3_5_9_i;
wire signed [`CalcTempBus]          temp_b3_5_10_r;
wire signed [`CalcTempBus]          temp_b3_5_10_i;
wire signed [`CalcTempBus]          temp_b3_5_11_r;
wire signed [`CalcTempBus]          temp_b3_5_11_i;
wire signed [`CalcTempBus]          temp_b3_5_12_r;
wire signed [`CalcTempBus]          temp_b3_5_12_i;
wire signed [`CalcTempBus]          temp_b3_5_13_r;
wire signed [`CalcTempBus]          temp_b3_5_13_i;
wire signed [`CalcTempBus]          temp_b3_5_14_r;
wire signed [`CalcTempBus]          temp_b3_5_14_i;
wire signed [`CalcTempBus]          temp_b3_5_15_r;
wire signed [`CalcTempBus]          temp_b3_5_15_i;
wire signed [`CalcTempBus]          temp_b3_5_16_r;
wire signed [`CalcTempBus]          temp_b3_5_16_i;
wire signed [`CalcTempBus]          temp_b3_6_1_r;
wire signed [`CalcTempBus]          temp_b3_6_1_i;
wire signed [`CalcTempBus]          temp_b3_6_2_r;
wire signed [`CalcTempBus]          temp_b3_6_2_i;
wire signed [`CalcTempBus]          temp_b3_6_3_r;
wire signed [`CalcTempBus]          temp_b3_6_3_i;
wire signed [`CalcTempBus]          temp_b3_6_4_r;
wire signed [`CalcTempBus]          temp_b3_6_4_i;
wire signed [`CalcTempBus]          temp_b3_6_5_r;
wire signed [`CalcTempBus]          temp_b3_6_5_i;
wire signed [`CalcTempBus]          temp_b3_6_6_r;
wire signed [`CalcTempBus]          temp_b3_6_6_i;
wire signed [`CalcTempBus]          temp_b3_6_7_r;
wire signed [`CalcTempBus]          temp_b3_6_7_i;
wire signed [`CalcTempBus]          temp_b3_6_8_r;
wire signed [`CalcTempBus]          temp_b3_6_8_i;
wire signed [`CalcTempBus]          temp_b3_6_9_r;
wire signed [`CalcTempBus]          temp_b3_6_9_i;
wire signed [`CalcTempBus]          temp_b3_6_10_r;
wire signed [`CalcTempBus]          temp_b3_6_10_i;
wire signed [`CalcTempBus]          temp_b3_6_11_r;
wire signed [`CalcTempBus]          temp_b3_6_11_i;
wire signed [`CalcTempBus]          temp_b3_6_12_r;
wire signed [`CalcTempBus]          temp_b3_6_12_i;
wire signed [`CalcTempBus]          temp_b3_6_13_r;
wire signed [`CalcTempBus]          temp_b3_6_13_i;
wire signed [`CalcTempBus]          temp_b3_6_14_r;
wire signed [`CalcTempBus]          temp_b3_6_14_i;
wire signed [`CalcTempBus]          temp_b3_6_15_r;
wire signed [`CalcTempBus]          temp_b3_6_15_i;
wire signed [`CalcTempBus]          temp_b3_6_16_r;
wire signed [`CalcTempBus]          temp_b3_6_16_i;
wire signed [`CalcTempBus]          temp_b3_7_1_r;
wire signed [`CalcTempBus]          temp_b3_7_1_i;
wire signed [`CalcTempBus]          temp_b3_7_2_r;
wire signed [`CalcTempBus]          temp_b3_7_2_i;
wire signed [`CalcTempBus]          temp_b3_7_3_r;
wire signed [`CalcTempBus]          temp_b3_7_3_i;
wire signed [`CalcTempBus]          temp_b3_7_4_r;
wire signed [`CalcTempBus]          temp_b3_7_4_i;
wire signed [`CalcTempBus]          temp_b3_7_5_r;
wire signed [`CalcTempBus]          temp_b3_7_5_i;
wire signed [`CalcTempBus]          temp_b3_7_6_r;
wire signed [`CalcTempBus]          temp_b3_7_6_i;
wire signed [`CalcTempBus]          temp_b3_7_7_r;
wire signed [`CalcTempBus]          temp_b3_7_7_i;
wire signed [`CalcTempBus]          temp_b3_7_8_r;
wire signed [`CalcTempBus]          temp_b3_7_8_i;
wire signed [`CalcTempBus]          temp_b3_7_9_r;
wire signed [`CalcTempBus]          temp_b3_7_9_i;
wire signed [`CalcTempBus]          temp_b3_7_10_r;
wire signed [`CalcTempBus]          temp_b3_7_10_i;
wire signed [`CalcTempBus]          temp_b3_7_11_r;
wire signed [`CalcTempBus]          temp_b3_7_11_i;
wire signed [`CalcTempBus]          temp_b3_7_12_r;
wire signed [`CalcTempBus]          temp_b3_7_12_i;
wire signed [`CalcTempBus]          temp_b3_7_13_r;
wire signed [`CalcTempBus]          temp_b3_7_13_i;
wire signed [`CalcTempBus]          temp_b3_7_14_r;
wire signed [`CalcTempBus]          temp_b3_7_14_i;
wire signed [`CalcTempBus]          temp_b3_7_15_r;
wire signed [`CalcTempBus]          temp_b3_7_15_i;
wire signed [`CalcTempBus]          temp_b3_7_16_r;
wire signed [`CalcTempBus]          temp_b3_7_16_i;
wire signed [`CalcTempBus]          temp_b3_8_1_r;
wire signed [`CalcTempBus]          temp_b3_8_1_i;
wire signed [`CalcTempBus]          temp_b3_8_2_r;
wire signed [`CalcTempBus]          temp_b3_8_2_i;
wire signed [`CalcTempBus]          temp_b3_8_3_r;
wire signed [`CalcTempBus]          temp_b3_8_3_i;
wire signed [`CalcTempBus]          temp_b3_8_4_r;
wire signed [`CalcTempBus]          temp_b3_8_4_i;
wire signed [`CalcTempBus]          temp_b3_8_5_r;
wire signed [`CalcTempBus]          temp_b3_8_5_i;
wire signed [`CalcTempBus]          temp_b3_8_6_r;
wire signed [`CalcTempBus]          temp_b3_8_6_i;
wire signed [`CalcTempBus]          temp_b3_8_7_r;
wire signed [`CalcTempBus]          temp_b3_8_7_i;
wire signed [`CalcTempBus]          temp_b3_8_8_r;
wire signed [`CalcTempBus]          temp_b3_8_8_i;
wire signed [`CalcTempBus]          temp_b3_8_9_r;
wire signed [`CalcTempBus]          temp_b3_8_9_i;
wire signed [`CalcTempBus]          temp_b3_8_10_r;
wire signed [`CalcTempBus]          temp_b3_8_10_i;
wire signed [`CalcTempBus]          temp_b3_8_11_r;
wire signed [`CalcTempBus]          temp_b3_8_11_i;
wire signed [`CalcTempBus]          temp_b3_8_12_r;
wire signed [`CalcTempBus]          temp_b3_8_12_i;
wire signed [`CalcTempBus]          temp_b3_8_13_r;
wire signed [`CalcTempBus]          temp_b3_8_13_i;
wire signed [`CalcTempBus]          temp_b3_8_14_r;
wire signed [`CalcTempBus]          temp_b3_8_14_i;
wire signed [`CalcTempBus]          temp_b3_8_15_r;
wire signed [`CalcTempBus]          temp_b3_8_15_i;
wire signed [`CalcTempBus]          temp_b3_8_16_r;
wire signed [`CalcTempBus]          temp_b3_8_16_i;
wire signed [`CalcTempBus]          temp_b3_9_1_r;
wire signed [`CalcTempBus]          temp_b3_9_1_i;
wire signed [`CalcTempBus]          temp_b3_9_2_r;
wire signed [`CalcTempBus]          temp_b3_9_2_i;
wire signed [`CalcTempBus]          temp_b3_9_3_r;
wire signed [`CalcTempBus]          temp_b3_9_3_i;
wire signed [`CalcTempBus]          temp_b3_9_4_r;
wire signed [`CalcTempBus]          temp_b3_9_4_i;
wire signed [`CalcTempBus]          temp_b3_9_5_r;
wire signed [`CalcTempBus]          temp_b3_9_5_i;
wire signed [`CalcTempBus]          temp_b3_9_6_r;
wire signed [`CalcTempBus]          temp_b3_9_6_i;
wire signed [`CalcTempBus]          temp_b3_9_7_r;
wire signed [`CalcTempBus]          temp_b3_9_7_i;
wire signed [`CalcTempBus]          temp_b3_9_8_r;
wire signed [`CalcTempBus]          temp_b3_9_8_i;
wire signed [`CalcTempBus]          temp_b3_9_9_r;
wire signed [`CalcTempBus]          temp_b3_9_9_i;
wire signed [`CalcTempBus]          temp_b3_9_10_r;
wire signed [`CalcTempBus]          temp_b3_9_10_i;
wire signed [`CalcTempBus]          temp_b3_9_11_r;
wire signed [`CalcTempBus]          temp_b3_9_11_i;
wire signed [`CalcTempBus]          temp_b3_9_12_r;
wire signed [`CalcTempBus]          temp_b3_9_12_i;
wire signed [`CalcTempBus]          temp_b3_9_13_r;
wire signed [`CalcTempBus]          temp_b3_9_13_i;
wire signed [`CalcTempBus]          temp_b3_9_14_r;
wire signed [`CalcTempBus]          temp_b3_9_14_i;
wire signed [`CalcTempBus]          temp_b3_9_15_r;
wire signed [`CalcTempBus]          temp_b3_9_15_i;
wire signed [`CalcTempBus]          temp_b3_9_16_r;
wire signed [`CalcTempBus]          temp_b3_9_16_i;
wire signed [`CalcTempBus]          temp_b3_10_1_r;
wire signed [`CalcTempBus]          temp_b3_10_1_i;
wire signed [`CalcTempBus]          temp_b3_10_2_r;
wire signed [`CalcTempBus]          temp_b3_10_2_i;
wire signed [`CalcTempBus]          temp_b3_10_3_r;
wire signed [`CalcTempBus]          temp_b3_10_3_i;
wire signed [`CalcTempBus]          temp_b3_10_4_r;
wire signed [`CalcTempBus]          temp_b3_10_4_i;
wire signed [`CalcTempBus]          temp_b3_10_5_r;
wire signed [`CalcTempBus]          temp_b3_10_5_i;
wire signed [`CalcTempBus]          temp_b3_10_6_r;
wire signed [`CalcTempBus]          temp_b3_10_6_i;
wire signed [`CalcTempBus]          temp_b3_10_7_r;
wire signed [`CalcTempBus]          temp_b3_10_7_i;
wire signed [`CalcTempBus]          temp_b3_10_8_r;
wire signed [`CalcTempBus]          temp_b3_10_8_i;
wire signed [`CalcTempBus]          temp_b3_10_9_r;
wire signed [`CalcTempBus]          temp_b3_10_9_i;
wire signed [`CalcTempBus]          temp_b3_10_10_r;
wire signed [`CalcTempBus]          temp_b3_10_10_i;
wire signed [`CalcTempBus]          temp_b3_10_11_r;
wire signed [`CalcTempBus]          temp_b3_10_11_i;
wire signed [`CalcTempBus]          temp_b3_10_12_r;
wire signed [`CalcTempBus]          temp_b3_10_12_i;
wire signed [`CalcTempBus]          temp_b3_10_13_r;
wire signed [`CalcTempBus]          temp_b3_10_13_i;
wire signed [`CalcTempBus]          temp_b3_10_14_r;
wire signed [`CalcTempBus]          temp_b3_10_14_i;
wire signed [`CalcTempBus]          temp_b3_10_15_r;
wire signed [`CalcTempBus]          temp_b3_10_15_i;
wire signed [`CalcTempBus]          temp_b3_10_16_r;
wire signed [`CalcTempBus]          temp_b3_10_16_i;
wire signed [`CalcTempBus]          temp_b3_11_1_r;
wire signed [`CalcTempBus]          temp_b3_11_1_i;
wire signed [`CalcTempBus]          temp_b3_11_2_r;
wire signed [`CalcTempBus]          temp_b3_11_2_i;
wire signed [`CalcTempBus]          temp_b3_11_3_r;
wire signed [`CalcTempBus]          temp_b3_11_3_i;
wire signed [`CalcTempBus]          temp_b3_11_4_r;
wire signed [`CalcTempBus]          temp_b3_11_4_i;
wire signed [`CalcTempBus]          temp_b3_11_5_r;
wire signed [`CalcTempBus]          temp_b3_11_5_i;
wire signed [`CalcTempBus]          temp_b3_11_6_r;
wire signed [`CalcTempBus]          temp_b3_11_6_i;
wire signed [`CalcTempBus]          temp_b3_11_7_r;
wire signed [`CalcTempBus]          temp_b3_11_7_i;
wire signed [`CalcTempBus]          temp_b3_11_8_r;
wire signed [`CalcTempBus]          temp_b3_11_8_i;
wire signed [`CalcTempBus]          temp_b3_11_9_r;
wire signed [`CalcTempBus]          temp_b3_11_9_i;
wire signed [`CalcTempBus]          temp_b3_11_10_r;
wire signed [`CalcTempBus]          temp_b3_11_10_i;
wire signed [`CalcTempBus]          temp_b3_11_11_r;
wire signed [`CalcTempBus]          temp_b3_11_11_i;
wire signed [`CalcTempBus]          temp_b3_11_12_r;
wire signed [`CalcTempBus]          temp_b3_11_12_i;
wire signed [`CalcTempBus]          temp_b3_11_13_r;
wire signed [`CalcTempBus]          temp_b3_11_13_i;
wire signed [`CalcTempBus]          temp_b3_11_14_r;
wire signed [`CalcTempBus]          temp_b3_11_14_i;
wire signed [`CalcTempBus]          temp_b3_11_15_r;
wire signed [`CalcTempBus]          temp_b3_11_15_i;
wire signed [`CalcTempBus]          temp_b3_11_16_r;
wire signed [`CalcTempBus]          temp_b3_11_16_i;
wire signed [`CalcTempBus]          temp_b3_12_1_r;
wire signed [`CalcTempBus]          temp_b3_12_1_i;
wire signed [`CalcTempBus]          temp_b3_12_2_r;
wire signed [`CalcTempBus]          temp_b3_12_2_i;
wire signed [`CalcTempBus]          temp_b3_12_3_r;
wire signed [`CalcTempBus]          temp_b3_12_3_i;
wire signed [`CalcTempBus]          temp_b3_12_4_r;
wire signed [`CalcTempBus]          temp_b3_12_4_i;
wire signed [`CalcTempBus]          temp_b3_12_5_r;
wire signed [`CalcTempBus]          temp_b3_12_5_i;
wire signed [`CalcTempBus]          temp_b3_12_6_r;
wire signed [`CalcTempBus]          temp_b3_12_6_i;
wire signed [`CalcTempBus]          temp_b3_12_7_r;
wire signed [`CalcTempBus]          temp_b3_12_7_i;
wire signed [`CalcTempBus]          temp_b3_12_8_r;
wire signed [`CalcTempBus]          temp_b3_12_8_i;
wire signed [`CalcTempBus]          temp_b3_12_9_r;
wire signed [`CalcTempBus]          temp_b3_12_9_i;
wire signed [`CalcTempBus]          temp_b3_12_10_r;
wire signed [`CalcTempBus]          temp_b3_12_10_i;
wire signed [`CalcTempBus]          temp_b3_12_11_r;
wire signed [`CalcTempBus]          temp_b3_12_11_i;
wire signed [`CalcTempBus]          temp_b3_12_12_r;
wire signed [`CalcTempBus]          temp_b3_12_12_i;
wire signed [`CalcTempBus]          temp_b3_12_13_r;
wire signed [`CalcTempBus]          temp_b3_12_13_i;
wire signed [`CalcTempBus]          temp_b3_12_14_r;
wire signed [`CalcTempBus]          temp_b3_12_14_i;
wire signed [`CalcTempBus]          temp_b3_12_15_r;
wire signed [`CalcTempBus]          temp_b3_12_15_i;
wire signed [`CalcTempBus]          temp_b3_12_16_r;
wire signed [`CalcTempBus]          temp_b3_12_16_i;
wire signed [`CalcTempBus]          temp_b3_13_1_r;
wire signed [`CalcTempBus]          temp_b3_13_1_i;
wire signed [`CalcTempBus]          temp_b3_13_2_r;
wire signed [`CalcTempBus]          temp_b3_13_2_i;
wire signed [`CalcTempBus]          temp_b3_13_3_r;
wire signed [`CalcTempBus]          temp_b3_13_3_i;
wire signed [`CalcTempBus]          temp_b3_13_4_r;
wire signed [`CalcTempBus]          temp_b3_13_4_i;
wire signed [`CalcTempBus]          temp_b3_13_5_r;
wire signed [`CalcTempBus]          temp_b3_13_5_i;
wire signed [`CalcTempBus]          temp_b3_13_6_r;
wire signed [`CalcTempBus]          temp_b3_13_6_i;
wire signed [`CalcTempBus]          temp_b3_13_7_r;
wire signed [`CalcTempBus]          temp_b3_13_7_i;
wire signed [`CalcTempBus]          temp_b3_13_8_r;
wire signed [`CalcTempBus]          temp_b3_13_8_i;
wire signed [`CalcTempBus]          temp_b3_13_9_r;
wire signed [`CalcTempBus]          temp_b3_13_9_i;
wire signed [`CalcTempBus]          temp_b3_13_10_r;
wire signed [`CalcTempBus]          temp_b3_13_10_i;
wire signed [`CalcTempBus]          temp_b3_13_11_r;
wire signed [`CalcTempBus]          temp_b3_13_11_i;
wire signed [`CalcTempBus]          temp_b3_13_12_r;
wire signed [`CalcTempBus]          temp_b3_13_12_i;
wire signed [`CalcTempBus]          temp_b3_13_13_r;
wire signed [`CalcTempBus]          temp_b3_13_13_i;
wire signed [`CalcTempBus]          temp_b3_13_14_r;
wire signed [`CalcTempBus]          temp_b3_13_14_i;
wire signed [`CalcTempBus]          temp_b3_13_15_r;
wire signed [`CalcTempBus]          temp_b3_13_15_i;
wire signed [`CalcTempBus]          temp_b3_13_16_r;
wire signed [`CalcTempBus]          temp_b3_13_16_i;
wire signed [`CalcTempBus]          temp_b3_14_1_r;
wire signed [`CalcTempBus]          temp_b3_14_1_i;
wire signed [`CalcTempBus]          temp_b3_14_2_r;
wire signed [`CalcTempBus]          temp_b3_14_2_i;
wire signed [`CalcTempBus]          temp_b3_14_3_r;
wire signed [`CalcTempBus]          temp_b3_14_3_i;
wire signed [`CalcTempBus]          temp_b3_14_4_r;
wire signed [`CalcTempBus]          temp_b3_14_4_i;
wire signed [`CalcTempBus]          temp_b3_14_5_r;
wire signed [`CalcTempBus]          temp_b3_14_5_i;
wire signed [`CalcTempBus]          temp_b3_14_6_r;
wire signed [`CalcTempBus]          temp_b3_14_6_i;
wire signed [`CalcTempBus]          temp_b3_14_7_r;
wire signed [`CalcTempBus]          temp_b3_14_7_i;
wire signed [`CalcTempBus]          temp_b3_14_8_r;
wire signed [`CalcTempBus]          temp_b3_14_8_i;
wire signed [`CalcTempBus]          temp_b3_14_9_r;
wire signed [`CalcTempBus]          temp_b3_14_9_i;
wire signed [`CalcTempBus]          temp_b3_14_10_r;
wire signed [`CalcTempBus]          temp_b3_14_10_i;
wire signed [`CalcTempBus]          temp_b3_14_11_r;
wire signed [`CalcTempBus]          temp_b3_14_11_i;
wire signed [`CalcTempBus]          temp_b3_14_12_r;
wire signed [`CalcTempBus]          temp_b3_14_12_i;
wire signed [`CalcTempBus]          temp_b3_14_13_r;
wire signed [`CalcTempBus]          temp_b3_14_13_i;
wire signed [`CalcTempBus]          temp_b3_14_14_r;
wire signed [`CalcTempBus]          temp_b3_14_14_i;
wire signed [`CalcTempBus]          temp_b3_14_15_r;
wire signed [`CalcTempBus]          temp_b3_14_15_i;
wire signed [`CalcTempBus]          temp_b3_14_16_r;
wire signed [`CalcTempBus]          temp_b3_14_16_i;
wire signed [`CalcTempBus]          temp_b3_15_1_r;
wire signed [`CalcTempBus]          temp_b3_15_1_i;
wire signed [`CalcTempBus]          temp_b3_15_2_r;
wire signed [`CalcTempBus]          temp_b3_15_2_i;
wire signed [`CalcTempBus]          temp_b3_15_3_r;
wire signed [`CalcTempBus]          temp_b3_15_3_i;
wire signed [`CalcTempBus]          temp_b3_15_4_r;
wire signed [`CalcTempBus]          temp_b3_15_4_i;
wire signed [`CalcTempBus]          temp_b3_15_5_r;
wire signed [`CalcTempBus]          temp_b3_15_5_i;
wire signed [`CalcTempBus]          temp_b3_15_6_r;
wire signed [`CalcTempBus]          temp_b3_15_6_i;
wire signed [`CalcTempBus]          temp_b3_15_7_r;
wire signed [`CalcTempBus]          temp_b3_15_7_i;
wire signed [`CalcTempBus]          temp_b3_15_8_r;
wire signed [`CalcTempBus]          temp_b3_15_8_i;
wire signed [`CalcTempBus]          temp_b3_15_9_r;
wire signed [`CalcTempBus]          temp_b3_15_9_i;
wire signed [`CalcTempBus]          temp_b3_15_10_r;
wire signed [`CalcTempBus]          temp_b3_15_10_i;
wire signed [`CalcTempBus]          temp_b3_15_11_r;
wire signed [`CalcTempBus]          temp_b3_15_11_i;
wire signed [`CalcTempBus]          temp_b3_15_12_r;
wire signed [`CalcTempBus]          temp_b3_15_12_i;
wire signed [`CalcTempBus]          temp_b3_15_13_r;
wire signed [`CalcTempBus]          temp_b3_15_13_i;
wire signed [`CalcTempBus]          temp_b3_15_14_r;
wire signed [`CalcTempBus]          temp_b3_15_14_i;
wire signed [`CalcTempBus]          temp_b3_15_15_r;
wire signed [`CalcTempBus]          temp_b3_15_15_i;
wire signed [`CalcTempBus]          temp_b3_15_16_r;
wire signed [`CalcTempBus]          temp_b3_15_16_i;
wire signed [`CalcTempBus]          temp_b3_16_1_r;
wire signed [`CalcTempBus]          temp_b3_16_1_i;
wire signed [`CalcTempBus]          temp_b3_16_2_r;
wire signed [`CalcTempBus]          temp_b3_16_2_i;
wire signed [`CalcTempBus]          temp_b3_16_3_r;
wire signed [`CalcTempBus]          temp_b3_16_3_i;
wire signed [`CalcTempBus]          temp_b3_16_4_r;
wire signed [`CalcTempBus]          temp_b3_16_4_i;
wire signed [`CalcTempBus]          temp_b3_16_5_r;
wire signed [`CalcTempBus]          temp_b3_16_5_i;
wire signed [`CalcTempBus]          temp_b3_16_6_r;
wire signed [`CalcTempBus]          temp_b3_16_6_i;
wire signed [`CalcTempBus]          temp_b3_16_7_r;
wire signed [`CalcTempBus]          temp_b3_16_7_i;
wire signed [`CalcTempBus]          temp_b3_16_8_r;
wire signed [`CalcTempBus]          temp_b3_16_8_i;
wire signed [`CalcTempBus]          temp_b3_16_9_r;
wire signed [`CalcTempBus]          temp_b3_16_9_i;
wire signed [`CalcTempBus]          temp_b3_16_10_r;
wire signed [`CalcTempBus]          temp_b3_16_10_i;
wire signed [`CalcTempBus]          temp_b3_16_11_r;
wire signed [`CalcTempBus]          temp_b3_16_11_i;
wire signed [`CalcTempBus]          temp_b3_16_12_r;
wire signed [`CalcTempBus]          temp_b3_16_12_i;
wire signed [`CalcTempBus]          temp_b3_16_13_r;
wire signed [`CalcTempBus]          temp_b3_16_13_i;
wire signed [`CalcTempBus]          temp_b3_16_14_r;
wire signed [`CalcTempBus]          temp_b3_16_14_i;
wire signed [`CalcTempBus]          temp_b3_16_15_r;
wire signed [`CalcTempBus]          temp_b3_16_15_i;
wire signed [`CalcTempBus]          temp_b3_16_16_r;
wire signed [`CalcTempBus]          temp_b3_16_16_i;
wire signed [`CalcTempBus]          temp_b4_1_1_r;
wire signed [`CalcTempBus]          temp_b4_1_1_i;
wire signed [`CalcTempBus]          temp_b4_1_2_r;
wire signed [`CalcTempBus]          temp_b4_1_2_i;
wire signed [`CalcTempBus]          temp_b4_1_3_r;
wire signed [`CalcTempBus]          temp_b4_1_3_i;
wire signed [`CalcTempBus]          temp_b4_1_4_r;
wire signed [`CalcTempBus]          temp_b4_1_4_i;
wire signed [`CalcTempBus]          temp_b4_1_5_r;
wire signed [`CalcTempBus]          temp_b4_1_5_i;
wire signed [`CalcTempBus]          temp_b4_1_6_r;
wire signed [`CalcTempBus]          temp_b4_1_6_i;
wire signed [`CalcTempBus]          temp_b4_1_7_r;
wire signed [`CalcTempBus]          temp_b4_1_7_i;
wire signed [`CalcTempBus]          temp_b4_1_8_r;
wire signed [`CalcTempBus]          temp_b4_1_8_i;
wire signed [`CalcTempBus]          temp_b4_1_9_r;
wire signed [`CalcTempBus]          temp_b4_1_9_i;
wire signed [`CalcTempBus]          temp_b4_1_10_r;
wire signed [`CalcTempBus]          temp_b4_1_10_i;
wire signed [`CalcTempBus]          temp_b4_1_11_r;
wire signed [`CalcTempBus]          temp_b4_1_11_i;
wire signed [`CalcTempBus]          temp_b4_1_12_r;
wire signed [`CalcTempBus]          temp_b4_1_12_i;
wire signed [`CalcTempBus]          temp_b4_1_13_r;
wire signed [`CalcTempBus]          temp_b4_1_13_i;
wire signed [`CalcTempBus]          temp_b4_1_14_r;
wire signed [`CalcTempBus]          temp_b4_1_14_i;
wire signed [`CalcTempBus]          temp_b4_1_15_r;
wire signed [`CalcTempBus]          temp_b4_1_15_i;
wire signed [`CalcTempBus]          temp_b4_1_16_r;
wire signed [`CalcTempBus]          temp_b4_1_16_i;
wire signed [`CalcTempBus]          temp_b4_2_1_r;
wire signed [`CalcTempBus]          temp_b4_2_1_i;
wire signed [`CalcTempBus]          temp_b4_2_2_r;
wire signed [`CalcTempBus]          temp_b4_2_2_i;
wire signed [`CalcTempBus]          temp_b4_2_3_r;
wire signed [`CalcTempBus]          temp_b4_2_3_i;
wire signed [`CalcTempBus]          temp_b4_2_4_r;
wire signed [`CalcTempBus]          temp_b4_2_4_i;
wire signed [`CalcTempBus]          temp_b4_2_5_r;
wire signed [`CalcTempBus]          temp_b4_2_5_i;
wire signed [`CalcTempBus]          temp_b4_2_6_r;
wire signed [`CalcTempBus]          temp_b4_2_6_i;
wire signed [`CalcTempBus]          temp_b4_2_7_r;
wire signed [`CalcTempBus]          temp_b4_2_7_i;
wire signed [`CalcTempBus]          temp_b4_2_8_r;
wire signed [`CalcTempBus]          temp_b4_2_8_i;
wire signed [`CalcTempBus]          temp_b4_2_9_r;
wire signed [`CalcTempBus]          temp_b4_2_9_i;
wire signed [`CalcTempBus]          temp_b4_2_10_r;
wire signed [`CalcTempBus]          temp_b4_2_10_i;
wire signed [`CalcTempBus]          temp_b4_2_11_r;
wire signed [`CalcTempBus]          temp_b4_2_11_i;
wire signed [`CalcTempBus]          temp_b4_2_12_r;
wire signed [`CalcTempBus]          temp_b4_2_12_i;
wire signed [`CalcTempBus]          temp_b4_2_13_r;
wire signed [`CalcTempBus]          temp_b4_2_13_i;
wire signed [`CalcTempBus]          temp_b4_2_14_r;
wire signed [`CalcTempBus]          temp_b4_2_14_i;
wire signed [`CalcTempBus]          temp_b4_2_15_r;
wire signed [`CalcTempBus]          temp_b4_2_15_i;
wire signed [`CalcTempBus]          temp_b4_2_16_r;
wire signed [`CalcTempBus]          temp_b4_2_16_i;
wire signed [`CalcTempBus]          temp_b4_3_1_r;
wire signed [`CalcTempBus]          temp_b4_3_1_i;
wire signed [`CalcTempBus]          temp_b4_3_2_r;
wire signed [`CalcTempBus]          temp_b4_3_2_i;
wire signed [`CalcTempBus]          temp_b4_3_3_r;
wire signed [`CalcTempBus]          temp_b4_3_3_i;
wire signed [`CalcTempBus]          temp_b4_3_4_r;
wire signed [`CalcTempBus]          temp_b4_3_4_i;
wire signed [`CalcTempBus]          temp_b4_3_5_r;
wire signed [`CalcTempBus]          temp_b4_3_5_i;
wire signed [`CalcTempBus]          temp_b4_3_6_r;
wire signed [`CalcTempBus]          temp_b4_3_6_i;
wire signed [`CalcTempBus]          temp_b4_3_7_r;
wire signed [`CalcTempBus]          temp_b4_3_7_i;
wire signed [`CalcTempBus]          temp_b4_3_8_r;
wire signed [`CalcTempBus]          temp_b4_3_8_i;
wire signed [`CalcTempBus]          temp_b4_3_9_r;
wire signed [`CalcTempBus]          temp_b4_3_9_i;
wire signed [`CalcTempBus]          temp_b4_3_10_r;
wire signed [`CalcTempBus]          temp_b4_3_10_i;
wire signed [`CalcTempBus]          temp_b4_3_11_r;
wire signed [`CalcTempBus]          temp_b4_3_11_i;
wire signed [`CalcTempBus]          temp_b4_3_12_r;
wire signed [`CalcTempBus]          temp_b4_3_12_i;
wire signed [`CalcTempBus]          temp_b4_3_13_r;
wire signed [`CalcTempBus]          temp_b4_3_13_i;
wire signed [`CalcTempBus]          temp_b4_3_14_r;
wire signed [`CalcTempBus]          temp_b4_3_14_i;
wire signed [`CalcTempBus]          temp_b4_3_15_r;
wire signed [`CalcTempBus]          temp_b4_3_15_i;
wire signed [`CalcTempBus]          temp_b4_3_16_r;
wire signed [`CalcTempBus]          temp_b4_3_16_i;
wire signed [`CalcTempBus]          temp_b4_4_1_r;
wire signed [`CalcTempBus]          temp_b4_4_1_i;
wire signed [`CalcTempBus]          temp_b4_4_2_r;
wire signed [`CalcTempBus]          temp_b4_4_2_i;
wire signed [`CalcTempBus]          temp_b4_4_3_r;
wire signed [`CalcTempBus]          temp_b4_4_3_i;
wire signed [`CalcTempBus]          temp_b4_4_4_r;
wire signed [`CalcTempBus]          temp_b4_4_4_i;
wire signed [`CalcTempBus]          temp_b4_4_5_r;
wire signed [`CalcTempBus]          temp_b4_4_5_i;
wire signed [`CalcTempBus]          temp_b4_4_6_r;
wire signed [`CalcTempBus]          temp_b4_4_6_i;
wire signed [`CalcTempBus]          temp_b4_4_7_r;
wire signed [`CalcTempBus]          temp_b4_4_7_i;
wire signed [`CalcTempBus]          temp_b4_4_8_r;
wire signed [`CalcTempBus]          temp_b4_4_8_i;
wire signed [`CalcTempBus]          temp_b4_4_9_r;
wire signed [`CalcTempBus]          temp_b4_4_9_i;
wire signed [`CalcTempBus]          temp_b4_4_10_r;
wire signed [`CalcTempBus]          temp_b4_4_10_i;
wire signed [`CalcTempBus]          temp_b4_4_11_r;
wire signed [`CalcTempBus]          temp_b4_4_11_i;
wire signed [`CalcTempBus]          temp_b4_4_12_r;
wire signed [`CalcTempBus]          temp_b4_4_12_i;
wire signed [`CalcTempBus]          temp_b4_4_13_r;
wire signed [`CalcTempBus]          temp_b4_4_13_i;
wire signed [`CalcTempBus]          temp_b4_4_14_r;
wire signed [`CalcTempBus]          temp_b4_4_14_i;
wire signed [`CalcTempBus]          temp_b4_4_15_r;
wire signed [`CalcTempBus]          temp_b4_4_15_i;
wire signed [`CalcTempBus]          temp_b4_4_16_r;
wire signed [`CalcTempBus]          temp_b4_4_16_i;
wire signed [`CalcTempBus]          temp_b4_5_1_r;
wire signed [`CalcTempBus]          temp_b4_5_1_i;
wire signed [`CalcTempBus]          temp_b4_5_2_r;
wire signed [`CalcTempBus]          temp_b4_5_2_i;
wire signed [`CalcTempBus]          temp_b4_5_3_r;
wire signed [`CalcTempBus]          temp_b4_5_3_i;
wire signed [`CalcTempBus]          temp_b4_5_4_r;
wire signed [`CalcTempBus]          temp_b4_5_4_i;
wire signed [`CalcTempBus]          temp_b4_5_5_r;
wire signed [`CalcTempBus]          temp_b4_5_5_i;
wire signed [`CalcTempBus]          temp_b4_5_6_r;
wire signed [`CalcTempBus]          temp_b4_5_6_i;
wire signed [`CalcTempBus]          temp_b4_5_7_r;
wire signed [`CalcTempBus]          temp_b4_5_7_i;
wire signed [`CalcTempBus]          temp_b4_5_8_r;
wire signed [`CalcTempBus]          temp_b4_5_8_i;
wire signed [`CalcTempBus]          temp_b4_5_9_r;
wire signed [`CalcTempBus]          temp_b4_5_9_i;
wire signed [`CalcTempBus]          temp_b4_5_10_r;
wire signed [`CalcTempBus]          temp_b4_5_10_i;
wire signed [`CalcTempBus]          temp_b4_5_11_r;
wire signed [`CalcTempBus]          temp_b4_5_11_i;
wire signed [`CalcTempBus]          temp_b4_5_12_r;
wire signed [`CalcTempBus]          temp_b4_5_12_i;
wire signed [`CalcTempBus]          temp_b4_5_13_r;
wire signed [`CalcTempBus]          temp_b4_5_13_i;
wire signed [`CalcTempBus]          temp_b4_5_14_r;
wire signed [`CalcTempBus]          temp_b4_5_14_i;
wire signed [`CalcTempBus]          temp_b4_5_15_r;
wire signed [`CalcTempBus]          temp_b4_5_15_i;
wire signed [`CalcTempBus]          temp_b4_5_16_r;
wire signed [`CalcTempBus]          temp_b4_5_16_i;
wire signed [`CalcTempBus]          temp_b4_6_1_r;
wire signed [`CalcTempBus]          temp_b4_6_1_i;
wire signed [`CalcTempBus]          temp_b4_6_2_r;
wire signed [`CalcTempBus]          temp_b4_6_2_i;
wire signed [`CalcTempBus]          temp_b4_6_3_r;
wire signed [`CalcTempBus]          temp_b4_6_3_i;
wire signed [`CalcTempBus]          temp_b4_6_4_r;
wire signed [`CalcTempBus]          temp_b4_6_4_i;
wire signed [`CalcTempBus]          temp_b4_6_5_r;
wire signed [`CalcTempBus]          temp_b4_6_5_i;
wire signed [`CalcTempBus]          temp_b4_6_6_r;
wire signed [`CalcTempBus]          temp_b4_6_6_i;
wire signed [`CalcTempBus]          temp_b4_6_7_r;
wire signed [`CalcTempBus]          temp_b4_6_7_i;
wire signed [`CalcTempBus]          temp_b4_6_8_r;
wire signed [`CalcTempBus]          temp_b4_6_8_i;
wire signed [`CalcTempBus]          temp_b4_6_9_r;
wire signed [`CalcTempBus]          temp_b4_6_9_i;
wire signed [`CalcTempBus]          temp_b4_6_10_r;
wire signed [`CalcTempBus]          temp_b4_6_10_i;
wire signed [`CalcTempBus]          temp_b4_6_11_r;
wire signed [`CalcTempBus]          temp_b4_6_11_i;
wire signed [`CalcTempBus]          temp_b4_6_12_r;
wire signed [`CalcTempBus]          temp_b4_6_12_i;
wire signed [`CalcTempBus]          temp_b4_6_13_r;
wire signed [`CalcTempBus]          temp_b4_6_13_i;
wire signed [`CalcTempBus]          temp_b4_6_14_r;
wire signed [`CalcTempBus]          temp_b4_6_14_i;
wire signed [`CalcTempBus]          temp_b4_6_15_r;
wire signed [`CalcTempBus]          temp_b4_6_15_i;
wire signed [`CalcTempBus]          temp_b4_6_16_r;
wire signed [`CalcTempBus]          temp_b4_6_16_i;
wire signed [`CalcTempBus]          temp_b4_7_1_r;
wire signed [`CalcTempBus]          temp_b4_7_1_i;
wire signed [`CalcTempBus]          temp_b4_7_2_r;
wire signed [`CalcTempBus]          temp_b4_7_2_i;
wire signed [`CalcTempBus]          temp_b4_7_3_r;
wire signed [`CalcTempBus]          temp_b4_7_3_i;
wire signed [`CalcTempBus]          temp_b4_7_4_r;
wire signed [`CalcTempBus]          temp_b4_7_4_i;
wire signed [`CalcTempBus]          temp_b4_7_5_r;
wire signed [`CalcTempBus]          temp_b4_7_5_i;
wire signed [`CalcTempBus]          temp_b4_7_6_r;
wire signed [`CalcTempBus]          temp_b4_7_6_i;
wire signed [`CalcTempBus]          temp_b4_7_7_r;
wire signed [`CalcTempBus]          temp_b4_7_7_i;
wire signed [`CalcTempBus]          temp_b4_7_8_r;
wire signed [`CalcTempBus]          temp_b4_7_8_i;
wire signed [`CalcTempBus]          temp_b4_7_9_r;
wire signed [`CalcTempBus]          temp_b4_7_9_i;
wire signed [`CalcTempBus]          temp_b4_7_10_r;
wire signed [`CalcTempBus]          temp_b4_7_10_i;
wire signed [`CalcTempBus]          temp_b4_7_11_r;
wire signed [`CalcTempBus]          temp_b4_7_11_i;
wire signed [`CalcTempBus]          temp_b4_7_12_r;
wire signed [`CalcTempBus]          temp_b4_7_12_i;
wire signed [`CalcTempBus]          temp_b4_7_13_r;
wire signed [`CalcTempBus]          temp_b4_7_13_i;
wire signed [`CalcTempBus]          temp_b4_7_14_r;
wire signed [`CalcTempBus]          temp_b4_7_14_i;
wire signed [`CalcTempBus]          temp_b4_7_15_r;
wire signed [`CalcTempBus]          temp_b4_7_15_i;
wire signed [`CalcTempBus]          temp_b4_7_16_r;
wire signed [`CalcTempBus]          temp_b4_7_16_i;
wire signed [`CalcTempBus]          temp_b4_8_1_r;
wire signed [`CalcTempBus]          temp_b4_8_1_i;
wire signed [`CalcTempBus]          temp_b4_8_2_r;
wire signed [`CalcTempBus]          temp_b4_8_2_i;
wire signed [`CalcTempBus]          temp_b4_8_3_r;
wire signed [`CalcTempBus]          temp_b4_8_3_i;
wire signed [`CalcTempBus]          temp_b4_8_4_r;
wire signed [`CalcTempBus]          temp_b4_8_4_i;
wire signed [`CalcTempBus]          temp_b4_8_5_r;
wire signed [`CalcTempBus]          temp_b4_8_5_i;
wire signed [`CalcTempBus]          temp_b4_8_6_r;
wire signed [`CalcTempBus]          temp_b4_8_6_i;
wire signed [`CalcTempBus]          temp_b4_8_7_r;
wire signed [`CalcTempBus]          temp_b4_8_7_i;
wire signed [`CalcTempBus]          temp_b4_8_8_r;
wire signed [`CalcTempBus]          temp_b4_8_8_i;
wire signed [`CalcTempBus]          temp_b4_8_9_r;
wire signed [`CalcTempBus]          temp_b4_8_9_i;
wire signed [`CalcTempBus]          temp_b4_8_10_r;
wire signed [`CalcTempBus]          temp_b4_8_10_i;
wire signed [`CalcTempBus]          temp_b4_8_11_r;
wire signed [`CalcTempBus]          temp_b4_8_11_i;
wire signed [`CalcTempBus]          temp_b4_8_12_r;
wire signed [`CalcTempBus]          temp_b4_8_12_i;
wire signed [`CalcTempBus]          temp_b4_8_13_r;
wire signed [`CalcTempBus]          temp_b4_8_13_i;
wire signed [`CalcTempBus]          temp_b4_8_14_r;
wire signed [`CalcTempBus]          temp_b4_8_14_i;
wire signed [`CalcTempBus]          temp_b4_8_15_r;
wire signed [`CalcTempBus]          temp_b4_8_15_i;
wire signed [`CalcTempBus]          temp_b4_8_16_r;
wire signed [`CalcTempBus]          temp_b4_8_16_i;
wire signed [`CalcTempBus]          temp_b4_9_1_r;
wire signed [`CalcTempBus]          temp_b4_9_1_i;
wire signed [`CalcTempBus]          temp_b4_9_2_r;
wire signed [`CalcTempBus]          temp_b4_9_2_i;
wire signed [`CalcTempBus]          temp_b4_9_3_r;
wire signed [`CalcTempBus]          temp_b4_9_3_i;
wire signed [`CalcTempBus]          temp_b4_9_4_r;
wire signed [`CalcTempBus]          temp_b4_9_4_i;
wire signed [`CalcTempBus]          temp_b4_9_5_r;
wire signed [`CalcTempBus]          temp_b4_9_5_i;
wire signed [`CalcTempBus]          temp_b4_9_6_r;
wire signed [`CalcTempBus]          temp_b4_9_6_i;
wire signed [`CalcTempBus]          temp_b4_9_7_r;
wire signed [`CalcTempBus]          temp_b4_9_7_i;
wire signed [`CalcTempBus]          temp_b4_9_8_r;
wire signed [`CalcTempBus]          temp_b4_9_8_i;
wire signed [`CalcTempBus]          temp_b4_9_9_r;
wire signed [`CalcTempBus]          temp_b4_9_9_i;
wire signed [`CalcTempBus]          temp_b4_9_10_r;
wire signed [`CalcTempBus]          temp_b4_9_10_i;
wire signed [`CalcTempBus]          temp_b4_9_11_r;
wire signed [`CalcTempBus]          temp_b4_9_11_i;
wire signed [`CalcTempBus]          temp_b4_9_12_r;
wire signed [`CalcTempBus]          temp_b4_9_12_i;
wire signed [`CalcTempBus]          temp_b4_9_13_r;
wire signed [`CalcTempBus]          temp_b4_9_13_i;
wire signed [`CalcTempBus]          temp_b4_9_14_r;
wire signed [`CalcTempBus]          temp_b4_9_14_i;
wire signed [`CalcTempBus]          temp_b4_9_15_r;
wire signed [`CalcTempBus]          temp_b4_9_15_i;
wire signed [`CalcTempBus]          temp_b4_9_16_r;
wire signed [`CalcTempBus]          temp_b4_9_16_i;
wire signed [`CalcTempBus]          temp_b4_10_1_r;
wire signed [`CalcTempBus]          temp_b4_10_1_i;
wire signed [`CalcTempBus]          temp_b4_10_2_r;
wire signed [`CalcTempBus]          temp_b4_10_2_i;
wire signed [`CalcTempBus]          temp_b4_10_3_r;
wire signed [`CalcTempBus]          temp_b4_10_3_i;
wire signed [`CalcTempBus]          temp_b4_10_4_r;
wire signed [`CalcTempBus]          temp_b4_10_4_i;
wire signed [`CalcTempBus]          temp_b4_10_5_r;
wire signed [`CalcTempBus]          temp_b4_10_5_i;
wire signed [`CalcTempBus]          temp_b4_10_6_r;
wire signed [`CalcTempBus]          temp_b4_10_6_i;
wire signed [`CalcTempBus]          temp_b4_10_7_r;
wire signed [`CalcTempBus]          temp_b4_10_7_i;
wire signed [`CalcTempBus]          temp_b4_10_8_r;
wire signed [`CalcTempBus]          temp_b4_10_8_i;
wire signed [`CalcTempBus]          temp_b4_10_9_r;
wire signed [`CalcTempBus]          temp_b4_10_9_i;
wire signed [`CalcTempBus]          temp_b4_10_10_r;
wire signed [`CalcTempBus]          temp_b4_10_10_i;
wire signed [`CalcTempBus]          temp_b4_10_11_r;
wire signed [`CalcTempBus]          temp_b4_10_11_i;
wire signed [`CalcTempBus]          temp_b4_10_12_r;
wire signed [`CalcTempBus]          temp_b4_10_12_i;
wire signed [`CalcTempBus]          temp_b4_10_13_r;
wire signed [`CalcTempBus]          temp_b4_10_13_i;
wire signed [`CalcTempBus]          temp_b4_10_14_r;
wire signed [`CalcTempBus]          temp_b4_10_14_i;
wire signed [`CalcTempBus]          temp_b4_10_15_r;
wire signed [`CalcTempBus]          temp_b4_10_15_i;
wire signed [`CalcTempBus]          temp_b4_10_16_r;
wire signed [`CalcTempBus]          temp_b4_10_16_i;
wire signed [`CalcTempBus]          temp_b4_11_1_r;
wire signed [`CalcTempBus]          temp_b4_11_1_i;
wire signed [`CalcTempBus]          temp_b4_11_2_r;
wire signed [`CalcTempBus]          temp_b4_11_2_i;
wire signed [`CalcTempBus]          temp_b4_11_3_r;
wire signed [`CalcTempBus]          temp_b4_11_3_i;
wire signed [`CalcTempBus]          temp_b4_11_4_r;
wire signed [`CalcTempBus]          temp_b4_11_4_i;
wire signed [`CalcTempBus]          temp_b4_11_5_r;
wire signed [`CalcTempBus]          temp_b4_11_5_i;
wire signed [`CalcTempBus]          temp_b4_11_6_r;
wire signed [`CalcTempBus]          temp_b4_11_6_i;
wire signed [`CalcTempBus]          temp_b4_11_7_r;
wire signed [`CalcTempBus]          temp_b4_11_7_i;
wire signed [`CalcTempBus]          temp_b4_11_8_r;
wire signed [`CalcTempBus]          temp_b4_11_8_i;
wire signed [`CalcTempBus]          temp_b4_11_9_r;
wire signed [`CalcTempBus]          temp_b4_11_9_i;
wire signed [`CalcTempBus]          temp_b4_11_10_r;
wire signed [`CalcTempBus]          temp_b4_11_10_i;
wire signed [`CalcTempBus]          temp_b4_11_11_r;
wire signed [`CalcTempBus]          temp_b4_11_11_i;
wire signed [`CalcTempBus]          temp_b4_11_12_r;
wire signed [`CalcTempBus]          temp_b4_11_12_i;
wire signed [`CalcTempBus]          temp_b4_11_13_r;
wire signed [`CalcTempBus]          temp_b4_11_13_i;
wire signed [`CalcTempBus]          temp_b4_11_14_r;
wire signed [`CalcTempBus]          temp_b4_11_14_i;
wire signed [`CalcTempBus]          temp_b4_11_15_r;
wire signed [`CalcTempBus]          temp_b4_11_15_i;
wire signed [`CalcTempBus]          temp_b4_11_16_r;
wire signed [`CalcTempBus]          temp_b4_11_16_i;
wire signed [`CalcTempBus]          temp_b4_12_1_r;
wire signed [`CalcTempBus]          temp_b4_12_1_i;
wire signed [`CalcTempBus]          temp_b4_12_2_r;
wire signed [`CalcTempBus]          temp_b4_12_2_i;
wire signed [`CalcTempBus]          temp_b4_12_3_r;
wire signed [`CalcTempBus]          temp_b4_12_3_i;
wire signed [`CalcTempBus]          temp_b4_12_4_r;
wire signed [`CalcTempBus]          temp_b4_12_4_i;
wire signed [`CalcTempBus]          temp_b4_12_5_r;
wire signed [`CalcTempBus]          temp_b4_12_5_i;
wire signed [`CalcTempBus]          temp_b4_12_6_r;
wire signed [`CalcTempBus]          temp_b4_12_6_i;
wire signed [`CalcTempBus]          temp_b4_12_7_r;
wire signed [`CalcTempBus]          temp_b4_12_7_i;
wire signed [`CalcTempBus]          temp_b4_12_8_r;
wire signed [`CalcTempBus]          temp_b4_12_8_i;
wire signed [`CalcTempBus]          temp_b4_12_9_r;
wire signed [`CalcTempBus]          temp_b4_12_9_i;
wire signed [`CalcTempBus]          temp_b4_12_10_r;
wire signed [`CalcTempBus]          temp_b4_12_10_i;
wire signed [`CalcTempBus]          temp_b4_12_11_r;
wire signed [`CalcTempBus]          temp_b4_12_11_i;
wire signed [`CalcTempBus]          temp_b4_12_12_r;
wire signed [`CalcTempBus]          temp_b4_12_12_i;
wire signed [`CalcTempBus]          temp_b4_12_13_r;
wire signed [`CalcTempBus]          temp_b4_12_13_i;
wire signed [`CalcTempBus]          temp_b4_12_14_r;
wire signed [`CalcTempBus]          temp_b4_12_14_i;
wire signed [`CalcTempBus]          temp_b4_12_15_r;
wire signed [`CalcTempBus]          temp_b4_12_15_i;
wire signed [`CalcTempBus]          temp_b4_12_16_r;
wire signed [`CalcTempBus]          temp_b4_12_16_i;
wire signed [`CalcTempBus]          temp_b4_13_1_r;
wire signed [`CalcTempBus]          temp_b4_13_1_i;
wire signed [`CalcTempBus]          temp_b4_13_2_r;
wire signed [`CalcTempBus]          temp_b4_13_2_i;
wire signed [`CalcTempBus]          temp_b4_13_3_r;
wire signed [`CalcTempBus]          temp_b4_13_3_i;
wire signed [`CalcTempBus]          temp_b4_13_4_r;
wire signed [`CalcTempBus]          temp_b4_13_4_i;
wire signed [`CalcTempBus]          temp_b4_13_5_r;
wire signed [`CalcTempBus]          temp_b4_13_5_i;
wire signed [`CalcTempBus]          temp_b4_13_6_r;
wire signed [`CalcTempBus]          temp_b4_13_6_i;
wire signed [`CalcTempBus]          temp_b4_13_7_r;
wire signed [`CalcTempBus]          temp_b4_13_7_i;
wire signed [`CalcTempBus]          temp_b4_13_8_r;
wire signed [`CalcTempBus]          temp_b4_13_8_i;
wire signed [`CalcTempBus]          temp_b4_13_9_r;
wire signed [`CalcTempBus]          temp_b4_13_9_i;
wire signed [`CalcTempBus]          temp_b4_13_10_r;
wire signed [`CalcTempBus]          temp_b4_13_10_i;
wire signed [`CalcTempBus]          temp_b4_13_11_r;
wire signed [`CalcTempBus]          temp_b4_13_11_i;
wire signed [`CalcTempBus]          temp_b4_13_12_r;
wire signed [`CalcTempBus]          temp_b4_13_12_i;
wire signed [`CalcTempBus]          temp_b4_13_13_r;
wire signed [`CalcTempBus]          temp_b4_13_13_i;
wire signed [`CalcTempBus]          temp_b4_13_14_r;
wire signed [`CalcTempBus]          temp_b4_13_14_i;
wire signed [`CalcTempBus]          temp_b4_13_15_r;
wire signed [`CalcTempBus]          temp_b4_13_15_i;
wire signed [`CalcTempBus]          temp_b4_13_16_r;
wire signed [`CalcTempBus]          temp_b4_13_16_i;
wire signed [`CalcTempBus]          temp_b4_14_1_r;
wire signed [`CalcTempBus]          temp_b4_14_1_i;
wire signed [`CalcTempBus]          temp_b4_14_2_r;
wire signed [`CalcTempBus]          temp_b4_14_2_i;
wire signed [`CalcTempBus]          temp_b4_14_3_r;
wire signed [`CalcTempBus]          temp_b4_14_3_i;
wire signed [`CalcTempBus]          temp_b4_14_4_r;
wire signed [`CalcTempBus]          temp_b4_14_4_i;
wire signed [`CalcTempBus]          temp_b4_14_5_r;
wire signed [`CalcTempBus]          temp_b4_14_5_i;
wire signed [`CalcTempBus]          temp_b4_14_6_r;
wire signed [`CalcTempBus]          temp_b4_14_6_i;
wire signed [`CalcTempBus]          temp_b4_14_7_r;
wire signed [`CalcTempBus]          temp_b4_14_7_i;
wire signed [`CalcTempBus]          temp_b4_14_8_r;
wire signed [`CalcTempBus]          temp_b4_14_8_i;
wire signed [`CalcTempBus]          temp_b4_14_9_r;
wire signed [`CalcTempBus]          temp_b4_14_9_i;
wire signed [`CalcTempBus]          temp_b4_14_10_r;
wire signed [`CalcTempBus]          temp_b4_14_10_i;
wire signed [`CalcTempBus]          temp_b4_14_11_r;
wire signed [`CalcTempBus]          temp_b4_14_11_i;
wire signed [`CalcTempBus]          temp_b4_14_12_r;
wire signed [`CalcTempBus]          temp_b4_14_12_i;
wire signed [`CalcTempBus]          temp_b4_14_13_r;
wire signed [`CalcTempBus]          temp_b4_14_13_i;
wire signed [`CalcTempBus]          temp_b4_14_14_r;
wire signed [`CalcTempBus]          temp_b4_14_14_i;
wire signed [`CalcTempBus]          temp_b4_14_15_r;
wire signed [`CalcTempBus]          temp_b4_14_15_i;
wire signed [`CalcTempBus]          temp_b4_14_16_r;
wire signed [`CalcTempBus]          temp_b4_14_16_i;
wire signed [`CalcTempBus]          temp_b4_15_1_r;
wire signed [`CalcTempBus]          temp_b4_15_1_i;
wire signed [`CalcTempBus]          temp_b4_15_2_r;
wire signed [`CalcTempBus]          temp_b4_15_2_i;
wire signed [`CalcTempBus]          temp_b4_15_3_r;
wire signed [`CalcTempBus]          temp_b4_15_3_i;
wire signed [`CalcTempBus]          temp_b4_15_4_r;
wire signed [`CalcTempBus]          temp_b4_15_4_i;
wire signed [`CalcTempBus]          temp_b4_15_5_r;
wire signed [`CalcTempBus]          temp_b4_15_5_i;
wire signed [`CalcTempBus]          temp_b4_15_6_r;
wire signed [`CalcTempBus]          temp_b4_15_6_i;
wire signed [`CalcTempBus]          temp_b4_15_7_r;
wire signed [`CalcTempBus]          temp_b4_15_7_i;
wire signed [`CalcTempBus]          temp_b4_15_8_r;
wire signed [`CalcTempBus]          temp_b4_15_8_i;
wire signed [`CalcTempBus]          temp_b4_15_9_r;
wire signed [`CalcTempBus]          temp_b4_15_9_i;
wire signed [`CalcTempBus]          temp_b4_15_10_r;
wire signed [`CalcTempBus]          temp_b4_15_10_i;
wire signed [`CalcTempBus]          temp_b4_15_11_r;
wire signed [`CalcTempBus]          temp_b4_15_11_i;
wire signed [`CalcTempBus]          temp_b4_15_12_r;
wire signed [`CalcTempBus]          temp_b4_15_12_i;
wire signed [`CalcTempBus]          temp_b4_15_13_r;
wire signed [`CalcTempBus]          temp_b4_15_13_i;
wire signed [`CalcTempBus]          temp_b4_15_14_r;
wire signed [`CalcTempBus]          temp_b4_15_14_i;
wire signed [`CalcTempBus]          temp_b4_15_15_r;
wire signed [`CalcTempBus]          temp_b4_15_15_i;
wire signed [`CalcTempBus]          temp_b4_15_16_r;
wire signed [`CalcTempBus]          temp_b4_15_16_i;
wire signed [`CalcTempBus]          temp_b4_16_1_r;
wire signed [`CalcTempBus]          temp_b4_16_1_i;
wire signed [`CalcTempBus]          temp_b4_16_2_r;
wire signed [`CalcTempBus]          temp_b4_16_2_i;
wire signed [`CalcTempBus]          temp_b4_16_3_r;
wire signed [`CalcTempBus]          temp_b4_16_3_i;
wire signed [`CalcTempBus]          temp_b4_16_4_r;
wire signed [`CalcTempBus]          temp_b4_16_4_i;
wire signed [`CalcTempBus]          temp_b4_16_5_r;
wire signed [`CalcTempBus]          temp_b4_16_5_i;
wire signed [`CalcTempBus]          temp_b4_16_6_r;
wire signed [`CalcTempBus]          temp_b4_16_6_i;
wire signed [`CalcTempBus]          temp_b4_16_7_r;
wire signed [`CalcTempBus]          temp_b4_16_7_i;
wire signed [`CalcTempBus]          temp_b4_16_8_r;
wire signed [`CalcTempBus]          temp_b4_16_8_i;
wire signed [`CalcTempBus]          temp_b4_16_9_r;
wire signed [`CalcTempBus]          temp_b4_16_9_i;
wire signed [`CalcTempBus]          temp_b4_16_10_r;
wire signed [`CalcTempBus]          temp_b4_16_10_i;
wire signed [`CalcTempBus]          temp_b4_16_11_r;
wire signed [`CalcTempBus]          temp_b4_16_11_i;
wire signed [`CalcTempBus]          temp_b4_16_12_r;
wire signed [`CalcTempBus]          temp_b4_16_12_i;
wire signed [`CalcTempBus]          temp_b4_16_13_r;
wire signed [`CalcTempBus]          temp_b4_16_13_i;
wire signed [`CalcTempBus]          temp_b4_16_14_r;
wire signed [`CalcTempBus]          temp_b4_16_14_i;
wire signed [`CalcTempBus]          temp_b4_16_15_r;
wire signed [`CalcTempBus]          temp_b4_16_15_i;
wire signed [`CalcTempBus]          temp_b4_16_16_r;
wire signed [`CalcTempBus]          temp_b4_16_16_i;

/******************port map******************/
MULT MULT1 (clk,in_1_1_r,in_1_1_i,in_1_2_r,in_1_2_i,in_2_1_r,in_2_1_i,in_2_2_r,in_2_2_i,temp_m1_1_1_r,temp_m1_1_1_i,temp_m1_1_2_r,temp_m1_1_2_i,temp_m1_2_1_r,temp_m1_2_1_i,temp_m1_2_2_r,temp_m1_2_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly1 (clk,temp_m1_1_1_r,temp_m1_1_1_i,temp_m1_1_2_r,temp_m1_1_2_i,temp_m1_2_1_r,temp_m1_2_1_i,temp_m1_2_2_r,temp_m1_2_2_i,temp_b1_1_1_r,temp_b1_1_1_i,temp_b1_1_2_r,temp_b1_1_2_i,temp_b1_2_1_r,temp_b1_2_1_i,temp_b1_2_2_r,temp_b1_2_2_i);
MULT MULT2 (clk,in_1_3_r,in_1_3_i,in_1_4_r,in_1_4_i,in_2_3_r,in_2_3_i,in_2_4_r,in_2_4_i,temp_m1_1_3_r,temp_m1_1_3_i,temp_m1_1_4_r,temp_m1_1_4_i,temp_m1_2_3_r,temp_m1_2_3_i,temp_m1_2_4_r,temp_m1_2_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly2 (clk,temp_m1_1_3_r,temp_m1_1_3_i,temp_m1_1_4_r,temp_m1_1_4_i,temp_m1_2_3_r,temp_m1_2_3_i,temp_m1_2_4_r,temp_m1_2_4_i,temp_b1_1_3_r,temp_b1_1_3_i,temp_b1_1_4_r,temp_b1_1_4_i,temp_b1_2_3_r,temp_b1_2_3_i,temp_b1_2_4_r,temp_b1_2_4_i);
MULT MULT3 (clk,in_1_5_r,in_1_5_i,in_1_6_r,in_1_6_i,in_2_5_r,in_2_5_i,in_2_6_r,in_2_6_i,temp_m1_1_5_r,temp_m1_1_5_i,temp_m1_1_6_r,temp_m1_1_6_i,temp_m1_2_5_r,temp_m1_2_5_i,temp_m1_2_6_r,temp_m1_2_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly3 (clk,temp_m1_1_5_r,temp_m1_1_5_i,temp_m1_1_6_r,temp_m1_1_6_i,temp_m1_2_5_r,temp_m1_2_5_i,temp_m1_2_6_r,temp_m1_2_6_i,temp_b1_1_5_r,temp_b1_1_5_i,temp_b1_1_6_r,temp_b1_1_6_i,temp_b1_2_5_r,temp_b1_2_5_i,temp_b1_2_6_r,temp_b1_2_6_i);
MULT MULT4 (clk,in_1_7_r,in_1_7_i,in_1_8_r,in_1_8_i,in_2_7_r,in_2_7_i,in_2_8_r,in_2_8_i,temp_m1_1_7_r,temp_m1_1_7_i,temp_m1_1_8_r,temp_m1_1_8_i,temp_m1_2_7_r,temp_m1_2_7_i,temp_m1_2_8_r,temp_m1_2_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly4 (clk,temp_m1_1_7_r,temp_m1_1_7_i,temp_m1_1_8_r,temp_m1_1_8_i,temp_m1_2_7_r,temp_m1_2_7_i,temp_m1_2_8_r,temp_m1_2_8_i,temp_b1_1_7_r,temp_b1_1_7_i,temp_b1_1_8_r,temp_b1_1_8_i,temp_b1_2_7_r,temp_b1_2_7_i,temp_b1_2_8_r,temp_b1_2_8_i);
MULT MULT5 (clk,in_1_9_r,in_1_9_i,in_1_10_r,in_1_10_i,in_2_9_r,in_2_9_i,in_2_10_r,in_2_10_i,temp_m1_1_9_r,temp_m1_1_9_i,temp_m1_1_10_r,temp_m1_1_10_i,temp_m1_2_9_r,temp_m1_2_9_i,temp_m1_2_10_r,temp_m1_2_10_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly5 (clk,temp_m1_1_9_r,temp_m1_1_9_i,temp_m1_1_10_r,temp_m1_1_10_i,temp_m1_2_9_r,temp_m1_2_9_i,temp_m1_2_10_r,temp_m1_2_10_i,temp_b1_1_9_r,temp_b1_1_9_i,temp_b1_1_10_r,temp_b1_1_10_i,temp_b1_2_9_r,temp_b1_2_9_i,temp_b1_2_10_r,temp_b1_2_10_i);
MULT MULT6 (clk,in_1_11_r,in_1_11_i,in_1_12_r,in_1_12_i,in_2_11_r,in_2_11_i,in_2_12_r,in_2_12_i,temp_m1_1_11_r,temp_m1_1_11_i,temp_m1_1_12_r,temp_m1_1_12_i,temp_m1_2_11_r,temp_m1_2_11_i,temp_m1_2_12_r,temp_m1_2_12_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly6 (clk,temp_m1_1_11_r,temp_m1_1_11_i,temp_m1_1_12_r,temp_m1_1_12_i,temp_m1_2_11_r,temp_m1_2_11_i,temp_m1_2_12_r,temp_m1_2_12_i,temp_b1_1_11_r,temp_b1_1_11_i,temp_b1_1_12_r,temp_b1_1_12_i,temp_b1_2_11_r,temp_b1_2_11_i,temp_b1_2_12_r,temp_b1_2_12_i);
MULT MULT7 (clk,in_1_13_r,in_1_13_i,in_1_14_r,in_1_14_i,in_2_13_r,in_2_13_i,in_2_14_r,in_2_14_i,temp_m1_1_13_r,temp_m1_1_13_i,temp_m1_1_14_r,temp_m1_1_14_i,temp_m1_2_13_r,temp_m1_2_13_i,temp_m1_2_14_r,temp_m1_2_14_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly7 (clk,temp_m1_1_13_r,temp_m1_1_13_i,temp_m1_1_14_r,temp_m1_1_14_i,temp_m1_2_13_r,temp_m1_2_13_i,temp_m1_2_14_r,temp_m1_2_14_i,temp_b1_1_13_r,temp_b1_1_13_i,temp_b1_1_14_r,temp_b1_1_14_i,temp_b1_2_13_r,temp_b1_2_13_i,temp_b1_2_14_r,temp_b1_2_14_i);
MULT MULT8 (clk,in_1_15_r,in_1_15_i,in_1_16_r,in_1_16_i,in_2_15_r,in_2_15_i,in_2_16_r,in_2_16_i,temp_m1_1_15_r,temp_m1_1_15_i,temp_m1_1_16_r,temp_m1_1_16_i,temp_m1_2_15_r,temp_m1_2_15_i,temp_m1_2_16_r,temp_m1_2_16_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly8 (clk,temp_m1_1_15_r,temp_m1_1_15_i,temp_m1_1_16_r,temp_m1_1_16_i,temp_m1_2_15_r,temp_m1_2_15_i,temp_m1_2_16_r,temp_m1_2_16_i,temp_b1_1_15_r,temp_b1_1_15_i,temp_b1_1_16_r,temp_b1_1_16_i,temp_b1_2_15_r,temp_b1_2_15_i,temp_b1_2_16_r,temp_b1_2_16_i);
MULT MULT9 (clk,in_3_1_r,in_3_1_i,in_3_2_r,in_3_2_i,in_4_1_r,in_4_1_i,in_4_2_r,in_4_2_i,temp_m1_3_1_r,temp_m1_3_1_i,temp_m1_3_2_r,temp_m1_3_2_i,temp_m1_4_1_r,temp_m1_4_1_i,temp_m1_4_2_r,temp_m1_4_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly9 (clk,temp_m1_3_1_r,temp_m1_3_1_i,temp_m1_3_2_r,temp_m1_3_2_i,temp_m1_4_1_r,temp_m1_4_1_i,temp_m1_4_2_r,temp_m1_4_2_i,temp_b1_3_1_r,temp_b1_3_1_i,temp_b1_3_2_r,temp_b1_3_2_i,temp_b1_4_1_r,temp_b1_4_1_i,temp_b1_4_2_r,temp_b1_4_2_i);
MULT MULT10 (clk,in_3_3_r,in_3_3_i,in_3_4_r,in_3_4_i,in_4_3_r,in_4_3_i,in_4_4_r,in_4_4_i,temp_m1_3_3_r,temp_m1_3_3_i,temp_m1_3_4_r,temp_m1_3_4_i,temp_m1_4_3_r,temp_m1_4_3_i,temp_m1_4_4_r,temp_m1_4_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly10 (clk,temp_m1_3_3_r,temp_m1_3_3_i,temp_m1_3_4_r,temp_m1_3_4_i,temp_m1_4_3_r,temp_m1_4_3_i,temp_m1_4_4_r,temp_m1_4_4_i,temp_b1_3_3_r,temp_b1_3_3_i,temp_b1_3_4_r,temp_b1_3_4_i,temp_b1_4_3_r,temp_b1_4_3_i,temp_b1_4_4_r,temp_b1_4_4_i);
MULT MULT11 (clk,in_3_5_r,in_3_5_i,in_3_6_r,in_3_6_i,in_4_5_r,in_4_5_i,in_4_6_r,in_4_6_i,temp_m1_3_5_r,temp_m1_3_5_i,temp_m1_3_6_r,temp_m1_3_6_i,temp_m1_4_5_r,temp_m1_4_5_i,temp_m1_4_6_r,temp_m1_4_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly11 (clk,temp_m1_3_5_r,temp_m1_3_5_i,temp_m1_3_6_r,temp_m1_3_6_i,temp_m1_4_5_r,temp_m1_4_5_i,temp_m1_4_6_r,temp_m1_4_6_i,temp_b1_3_5_r,temp_b1_3_5_i,temp_b1_3_6_r,temp_b1_3_6_i,temp_b1_4_5_r,temp_b1_4_5_i,temp_b1_4_6_r,temp_b1_4_6_i);
MULT MULT12 (clk,in_3_7_r,in_3_7_i,in_3_8_r,in_3_8_i,in_4_7_r,in_4_7_i,in_4_8_r,in_4_8_i,temp_m1_3_7_r,temp_m1_3_7_i,temp_m1_3_8_r,temp_m1_3_8_i,temp_m1_4_7_r,temp_m1_4_7_i,temp_m1_4_8_r,temp_m1_4_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly12 (clk,temp_m1_3_7_r,temp_m1_3_7_i,temp_m1_3_8_r,temp_m1_3_8_i,temp_m1_4_7_r,temp_m1_4_7_i,temp_m1_4_8_r,temp_m1_4_8_i,temp_b1_3_7_r,temp_b1_3_7_i,temp_b1_3_8_r,temp_b1_3_8_i,temp_b1_4_7_r,temp_b1_4_7_i,temp_b1_4_8_r,temp_b1_4_8_i);
MULT MULT13 (clk,in_3_9_r,in_3_9_i,in_3_10_r,in_3_10_i,in_4_9_r,in_4_9_i,in_4_10_r,in_4_10_i,temp_m1_3_9_r,temp_m1_3_9_i,temp_m1_3_10_r,temp_m1_3_10_i,temp_m1_4_9_r,temp_m1_4_9_i,temp_m1_4_10_r,temp_m1_4_10_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly13 (clk,temp_m1_3_9_r,temp_m1_3_9_i,temp_m1_3_10_r,temp_m1_3_10_i,temp_m1_4_9_r,temp_m1_4_9_i,temp_m1_4_10_r,temp_m1_4_10_i,temp_b1_3_9_r,temp_b1_3_9_i,temp_b1_3_10_r,temp_b1_3_10_i,temp_b1_4_9_r,temp_b1_4_9_i,temp_b1_4_10_r,temp_b1_4_10_i);
MULT MULT14 (clk,in_3_11_r,in_3_11_i,in_3_12_r,in_3_12_i,in_4_11_r,in_4_11_i,in_4_12_r,in_4_12_i,temp_m1_3_11_r,temp_m1_3_11_i,temp_m1_3_12_r,temp_m1_3_12_i,temp_m1_4_11_r,temp_m1_4_11_i,temp_m1_4_12_r,temp_m1_4_12_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly14 (clk,temp_m1_3_11_r,temp_m1_3_11_i,temp_m1_3_12_r,temp_m1_3_12_i,temp_m1_4_11_r,temp_m1_4_11_i,temp_m1_4_12_r,temp_m1_4_12_i,temp_b1_3_11_r,temp_b1_3_11_i,temp_b1_3_12_r,temp_b1_3_12_i,temp_b1_4_11_r,temp_b1_4_11_i,temp_b1_4_12_r,temp_b1_4_12_i);
MULT MULT15 (clk,in_3_13_r,in_3_13_i,in_3_14_r,in_3_14_i,in_4_13_r,in_4_13_i,in_4_14_r,in_4_14_i,temp_m1_3_13_r,temp_m1_3_13_i,temp_m1_3_14_r,temp_m1_3_14_i,temp_m1_4_13_r,temp_m1_4_13_i,temp_m1_4_14_r,temp_m1_4_14_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly15 (clk,temp_m1_3_13_r,temp_m1_3_13_i,temp_m1_3_14_r,temp_m1_3_14_i,temp_m1_4_13_r,temp_m1_4_13_i,temp_m1_4_14_r,temp_m1_4_14_i,temp_b1_3_13_r,temp_b1_3_13_i,temp_b1_3_14_r,temp_b1_3_14_i,temp_b1_4_13_r,temp_b1_4_13_i,temp_b1_4_14_r,temp_b1_4_14_i);
MULT MULT16 (clk,in_3_15_r,in_3_15_i,in_3_16_r,in_3_16_i,in_4_15_r,in_4_15_i,in_4_16_r,in_4_16_i,temp_m1_3_15_r,temp_m1_3_15_i,temp_m1_3_16_r,temp_m1_3_16_i,temp_m1_4_15_r,temp_m1_4_15_i,temp_m1_4_16_r,temp_m1_4_16_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly16 (clk,temp_m1_3_15_r,temp_m1_3_15_i,temp_m1_3_16_r,temp_m1_3_16_i,temp_m1_4_15_r,temp_m1_4_15_i,temp_m1_4_16_r,temp_m1_4_16_i,temp_b1_3_15_r,temp_b1_3_15_i,temp_b1_3_16_r,temp_b1_3_16_i,temp_b1_4_15_r,temp_b1_4_15_i,temp_b1_4_16_r,temp_b1_4_16_i);
MULT MULT17 (clk,in_5_1_r,in_5_1_i,in_5_2_r,in_5_2_i,in_6_1_r,in_6_1_i,in_6_2_r,in_6_2_i,temp_m1_5_1_r,temp_m1_5_1_i,temp_m1_5_2_r,temp_m1_5_2_i,temp_m1_6_1_r,temp_m1_6_1_i,temp_m1_6_2_r,temp_m1_6_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly17 (clk,temp_m1_5_1_r,temp_m1_5_1_i,temp_m1_5_2_r,temp_m1_5_2_i,temp_m1_6_1_r,temp_m1_6_1_i,temp_m1_6_2_r,temp_m1_6_2_i,temp_b1_5_1_r,temp_b1_5_1_i,temp_b1_5_2_r,temp_b1_5_2_i,temp_b1_6_1_r,temp_b1_6_1_i,temp_b1_6_2_r,temp_b1_6_2_i);
MULT MULT18 (clk,in_5_3_r,in_5_3_i,in_5_4_r,in_5_4_i,in_6_3_r,in_6_3_i,in_6_4_r,in_6_4_i,temp_m1_5_3_r,temp_m1_5_3_i,temp_m1_5_4_r,temp_m1_5_4_i,temp_m1_6_3_r,temp_m1_6_3_i,temp_m1_6_4_r,temp_m1_6_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly18 (clk,temp_m1_5_3_r,temp_m1_5_3_i,temp_m1_5_4_r,temp_m1_5_4_i,temp_m1_6_3_r,temp_m1_6_3_i,temp_m1_6_4_r,temp_m1_6_4_i,temp_b1_5_3_r,temp_b1_5_3_i,temp_b1_5_4_r,temp_b1_5_4_i,temp_b1_6_3_r,temp_b1_6_3_i,temp_b1_6_4_r,temp_b1_6_4_i);
MULT MULT19 (clk,in_5_5_r,in_5_5_i,in_5_6_r,in_5_6_i,in_6_5_r,in_6_5_i,in_6_6_r,in_6_6_i,temp_m1_5_5_r,temp_m1_5_5_i,temp_m1_5_6_r,temp_m1_5_6_i,temp_m1_6_5_r,temp_m1_6_5_i,temp_m1_6_6_r,temp_m1_6_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly19 (clk,temp_m1_5_5_r,temp_m1_5_5_i,temp_m1_5_6_r,temp_m1_5_6_i,temp_m1_6_5_r,temp_m1_6_5_i,temp_m1_6_6_r,temp_m1_6_6_i,temp_b1_5_5_r,temp_b1_5_5_i,temp_b1_5_6_r,temp_b1_5_6_i,temp_b1_6_5_r,temp_b1_6_5_i,temp_b1_6_6_r,temp_b1_6_6_i);
MULT MULT20 (clk,in_5_7_r,in_5_7_i,in_5_8_r,in_5_8_i,in_6_7_r,in_6_7_i,in_6_8_r,in_6_8_i,temp_m1_5_7_r,temp_m1_5_7_i,temp_m1_5_8_r,temp_m1_5_8_i,temp_m1_6_7_r,temp_m1_6_7_i,temp_m1_6_8_r,temp_m1_6_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly20 (clk,temp_m1_5_7_r,temp_m1_5_7_i,temp_m1_5_8_r,temp_m1_5_8_i,temp_m1_6_7_r,temp_m1_6_7_i,temp_m1_6_8_r,temp_m1_6_8_i,temp_b1_5_7_r,temp_b1_5_7_i,temp_b1_5_8_r,temp_b1_5_8_i,temp_b1_6_7_r,temp_b1_6_7_i,temp_b1_6_8_r,temp_b1_6_8_i);
MULT MULT21 (clk,in_5_9_r,in_5_9_i,in_5_10_r,in_5_10_i,in_6_9_r,in_6_9_i,in_6_10_r,in_6_10_i,temp_m1_5_9_r,temp_m1_5_9_i,temp_m1_5_10_r,temp_m1_5_10_i,temp_m1_6_9_r,temp_m1_6_9_i,temp_m1_6_10_r,temp_m1_6_10_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly21 (clk,temp_m1_5_9_r,temp_m1_5_9_i,temp_m1_5_10_r,temp_m1_5_10_i,temp_m1_6_9_r,temp_m1_6_9_i,temp_m1_6_10_r,temp_m1_6_10_i,temp_b1_5_9_r,temp_b1_5_9_i,temp_b1_5_10_r,temp_b1_5_10_i,temp_b1_6_9_r,temp_b1_6_9_i,temp_b1_6_10_r,temp_b1_6_10_i);
MULT MULT22 (clk,in_5_11_r,in_5_11_i,in_5_12_r,in_5_12_i,in_6_11_r,in_6_11_i,in_6_12_r,in_6_12_i,temp_m1_5_11_r,temp_m1_5_11_i,temp_m1_5_12_r,temp_m1_5_12_i,temp_m1_6_11_r,temp_m1_6_11_i,temp_m1_6_12_r,temp_m1_6_12_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly22 (clk,temp_m1_5_11_r,temp_m1_5_11_i,temp_m1_5_12_r,temp_m1_5_12_i,temp_m1_6_11_r,temp_m1_6_11_i,temp_m1_6_12_r,temp_m1_6_12_i,temp_b1_5_11_r,temp_b1_5_11_i,temp_b1_5_12_r,temp_b1_5_12_i,temp_b1_6_11_r,temp_b1_6_11_i,temp_b1_6_12_r,temp_b1_6_12_i);
MULT MULT23 (clk,in_5_13_r,in_5_13_i,in_5_14_r,in_5_14_i,in_6_13_r,in_6_13_i,in_6_14_r,in_6_14_i,temp_m1_5_13_r,temp_m1_5_13_i,temp_m1_5_14_r,temp_m1_5_14_i,temp_m1_6_13_r,temp_m1_6_13_i,temp_m1_6_14_r,temp_m1_6_14_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly23 (clk,temp_m1_5_13_r,temp_m1_5_13_i,temp_m1_5_14_r,temp_m1_5_14_i,temp_m1_6_13_r,temp_m1_6_13_i,temp_m1_6_14_r,temp_m1_6_14_i,temp_b1_5_13_r,temp_b1_5_13_i,temp_b1_5_14_r,temp_b1_5_14_i,temp_b1_6_13_r,temp_b1_6_13_i,temp_b1_6_14_r,temp_b1_6_14_i);
MULT MULT24 (clk,in_5_15_r,in_5_15_i,in_5_16_r,in_5_16_i,in_6_15_r,in_6_15_i,in_6_16_r,in_6_16_i,temp_m1_5_15_r,temp_m1_5_15_i,temp_m1_5_16_r,temp_m1_5_16_i,temp_m1_6_15_r,temp_m1_6_15_i,temp_m1_6_16_r,temp_m1_6_16_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly24 (clk,temp_m1_5_15_r,temp_m1_5_15_i,temp_m1_5_16_r,temp_m1_5_16_i,temp_m1_6_15_r,temp_m1_6_15_i,temp_m1_6_16_r,temp_m1_6_16_i,temp_b1_5_15_r,temp_b1_5_15_i,temp_b1_5_16_r,temp_b1_5_16_i,temp_b1_6_15_r,temp_b1_6_15_i,temp_b1_6_16_r,temp_b1_6_16_i);
MULT MULT25 (clk,in_7_1_r,in_7_1_i,in_7_2_r,in_7_2_i,in_8_1_r,in_8_1_i,in_8_2_r,in_8_2_i,temp_m1_7_1_r,temp_m1_7_1_i,temp_m1_7_2_r,temp_m1_7_2_i,temp_m1_8_1_r,temp_m1_8_1_i,temp_m1_8_2_r,temp_m1_8_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly25 (clk,temp_m1_7_1_r,temp_m1_7_1_i,temp_m1_7_2_r,temp_m1_7_2_i,temp_m1_8_1_r,temp_m1_8_1_i,temp_m1_8_2_r,temp_m1_8_2_i,temp_b1_7_1_r,temp_b1_7_1_i,temp_b1_7_2_r,temp_b1_7_2_i,temp_b1_8_1_r,temp_b1_8_1_i,temp_b1_8_2_r,temp_b1_8_2_i);
MULT MULT26 (clk,in_7_3_r,in_7_3_i,in_7_4_r,in_7_4_i,in_8_3_r,in_8_3_i,in_8_4_r,in_8_4_i,temp_m1_7_3_r,temp_m1_7_3_i,temp_m1_7_4_r,temp_m1_7_4_i,temp_m1_8_3_r,temp_m1_8_3_i,temp_m1_8_4_r,temp_m1_8_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly26 (clk,temp_m1_7_3_r,temp_m1_7_3_i,temp_m1_7_4_r,temp_m1_7_4_i,temp_m1_8_3_r,temp_m1_8_3_i,temp_m1_8_4_r,temp_m1_8_4_i,temp_b1_7_3_r,temp_b1_7_3_i,temp_b1_7_4_r,temp_b1_7_4_i,temp_b1_8_3_r,temp_b1_8_3_i,temp_b1_8_4_r,temp_b1_8_4_i);
MULT MULT27 (clk,in_7_5_r,in_7_5_i,in_7_6_r,in_7_6_i,in_8_5_r,in_8_5_i,in_8_6_r,in_8_6_i,temp_m1_7_5_r,temp_m1_7_5_i,temp_m1_7_6_r,temp_m1_7_6_i,temp_m1_8_5_r,temp_m1_8_5_i,temp_m1_8_6_r,temp_m1_8_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly27 (clk,temp_m1_7_5_r,temp_m1_7_5_i,temp_m1_7_6_r,temp_m1_7_6_i,temp_m1_8_5_r,temp_m1_8_5_i,temp_m1_8_6_r,temp_m1_8_6_i,temp_b1_7_5_r,temp_b1_7_5_i,temp_b1_7_6_r,temp_b1_7_6_i,temp_b1_8_5_r,temp_b1_8_5_i,temp_b1_8_6_r,temp_b1_8_6_i);
MULT MULT28 (clk,in_7_7_r,in_7_7_i,in_7_8_r,in_7_8_i,in_8_7_r,in_8_7_i,in_8_8_r,in_8_8_i,temp_m1_7_7_r,temp_m1_7_7_i,temp_m1_7_8_r,temp_m1_7_8_i,temp_m1_8_7_r,temp_m1_8_7_i,temp_m1_8_8_r,temp_m1_8_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly28 (clk,temp_m1_7_7_r,temp_m1_7_7_i,temp_m1_7_8_r,temp_m1_7_8_i,temp_m1_8_7_r,temp_m1_8_7_i,temp_m1_8_8_r,temp_m1_8_8_i,temp_b1_7_7_r,temp_b1_7_7_i,temp_b1_7_8_r,temp_b1_7_8_i,temp_b1_8_7_r,temp_b1_8_7_i,temp_b1_8_8_r,temp_b1_8_8_i);
MULT MULT29 (clk,in_7_9_r,in_7_9_i,in_7_10_r,in_7_10_i,in_8_9_r,in_8_9_i,in_8_10_r,in_8_10_i,temp_m1_7_9_r,temp_m1_7_9_i,temp_m1_7_10_r,temp_m1_7_10_i,temp_m1_8_9_r,temp_m1_8_9_i,temp_m1_8_10_r,temp_m1_8_10_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly29 (clk,temp_m1_7_9_r,temp_m1_7_9_i,temp_m1_7_10_r,temp_m1_7_10_i,temp_m1_8_9_r,temp_m1_8_9_i,temp_m1_8_10_r,temp_m1_8_10_i,temp_b1_7_9_r,temp_b1_7_9_i,temp_b1_7_10_r,temp_b1_7_10_i,temp_b1_8_9_r,temp_b1_8_9_i,temp_b1_8_10_r,temp_b1_8_10_i);
MULT MULT30 (clk,in_7_11_r,in_7_11_i,in_7_12_r,in_7_12_i,in_8_11_r,in_8_11_i,in_8_12_r,in_8_12_i,temp_m1_7_11_r,temp_m1_7_11_i,temp_m1_7_12_r,temp_m1_7_12_i,temp_m1_8_11_r,temp_m1_8_11_i,temp_m1_8_12_r,temp_m1_8_12_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly30 (clk,temp_m1_7_11_r,temp_m1_7_11_i,temp_m1_7_12_r,temp_m1_7_12_i,temp_m1_8_11_r,temp_m1_8_11_i,temp_m1_8_12_r,temp_m1_8_12_i,temp_b1_7_11_r,temp_b1_7_11_i,temp_b1_7_12_r,temp_b1_7_12_i,temp_b1_8_11_r,temp_b1_8_11_i,temp_b1_8_12_r,temp_b1_8_12_i);
MULT MULT31 (clk,in_7_13_r,in_7_13_i,in_7_14_r,in_7_14_i,in_8_13_r,in_8_13_i,in_8_14_r,in_8_14_i,temp_m1_7_13_r,temp_m1_7_13_i,temp_m1_7_14_r,temp_m1_7_14_i,temp_m1_8_13_r,temp_m1_8_13_i,temp_m1_8_14_r,temp_m1_8_14_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly31 (clk,temp_m1_7_13_r,temp_m1_7_13_i,temp_m1_7_14_r,temp_m1_7_14_i,temp_m1_8_13_r,temp_m1_8_13_i,temp_m1_8_14_r,temp_m1_8_14_i,temp_b1_7_13_r,temp_b1_7_13_i,temp_b1_7_14_r,temp_b1_7_14_i,temp_b1_8_13_r,temp_b1_8_13_i,temp_b1_8_14_r,temp_b1_8_14_i);
MULT MULT32 (clk,in_7_15_r,in_7_15_i,in_7_16_r,in_7_16_i,in_8_15_r,in_8_15_i,in_8_16_r,in_8_16_i,temp_m1_7_15_r,temp_m1_7_15_i,temp_m1_7_16_r,temp_m1_7_16_i,temp_m1_8_15_r,temp_m1_8_15_i,temp_m1_8_16_r,temp_m1_8_16_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly32 (clk,temp_m1_7_15_r,temp_m1_7_15_i,temp_m1_7_16_r,temp_m1_7_16_i,temp_m1_8_15_r,temp_m1_8_15_i,temp_m1_8_16_r,temp_m1_8_16_i,temp_b1_7_15_r,temp_b1_7_15_i,temp_b1_7_16_r,temp_b1_7_16_i,temp_b1_8_15_r,temp_b1_8_15_i,temp_b1_8_16_r,temp_b1_8_16_i);
MULT MULT33 (clk,in_9_1_r,in_9_1_i,in_9_2_r,in_9_2_i,in_10_1_r,in_10_1_i,in_10_2_r,in_10_2_i,temp_m1_9_1_r,temp_m1_9_1_i,temp_m1_9_2_r,temp_m1_9_2_i,temp_m1_10_1_r,temp_m1_10_1_i,temp_m1_10_2_r,temp_m1_10_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly33 (clk,temp_m1_9_1_r,temp_m1_9_1_i,temp_m1_9_2_r,temp_m1_9_2_i,temp_m1_10_1_r,temp_m1_10_1_i,temp_m1_10_2_r,temp_m1_10_2_i,temp_b1_9_1_r,temp_b1_9_1_i,temp_b1_9_2_r,temp_b1_9_2_i,temp_b1_10_1_r,temp_b1_10_1_i,temp_b1_10_2_r,temp_b1_10_2_i);
MULT MULT34 (clk,in_9_3_r,in_9_3_i,in_9_4_r,in_9_4_i,in_10_3_r,in_10_3_i,in_10_4_r,in_10_4_i,temp_m1_9_3_r,temp_m1_9_3_i,temp_m1_9_4_r,temp_m1_9_4_i,temp_m1_10_3_r,temp_m1_10_3_i,temp_m1_10_4_r,temp_m1_10_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly34 (clk,temp_m1_9_3_r,temp_m1_9_3_i,temp_m1_9_4_r,temp_m1_9_4_i,temp_m1_10_3_r,temp_m1_10_3_i,temp_m1_10_4_r,temp_m1_10_4_i,temp_b1_9_3_r,temp_b1_9_3_i,temp_b1_9_4_r,temp_b1_9_4_i,temp_b1_10_3_r,temp_b1_10_3_i,temp_b1_10_4_r,temp_b1_10_4_i);
MULT MULT35 (clk,in_9_5_r,in_9_5_i,in_9_6_r,in_9_6_i,in_10_5_r,in_10_5_i,in_10_6_r,in_10_6_i,temp_m1_9_5_r,temp_m1_9_5_i,temp_m1_9_6_r,temp_m1_9_6_i,temp_m1_10_5_r,temp_m1_10_5_i,temp_m1_10_6_r,temp_m1_10_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly35 (clk,temp_m1_9_5_r,temp_m1_9_5_i,temp_m1_9_6_r,temp_m1_9_6_i,temp_m1_10_5_r,temp_m1_10_5_i,temp_m1_10_6_r,temp_m1_10_6_i,temp_b1_9_5_r,temp_b1_9_5_i,temp_b1_9_6_r,temp_b1_9_6_i,temp_b1_10_5_r,temp_b1_10_5_i,temp_b1_10_6_r,temp_b1_10_6_i);
MULT MULT36 (clk,in_9_7_r,in_9_7_i,in_9_8_r,in_9_8_i,in_10_7_r,in_10_7_i,in_10_8_r,in_10_8_i,temp_m1_9_7_r,temp_m1_9_7_i,temp_m1_9_8_r,temp_m1_9_8_i,temp_m1_10_7_r,temp_m1_10_7_i,temp_m1_10_8_r,temp_m1_10_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly36 (clk,temp_m1_9_7_r,temp_m1_9_7_i,temp_m1_9_8_r,temp_m1_9_8_i,temp_m1_10_7_r,temp_m1_10_7_i,temp_m1_10_8_r,temp_m1_10_8_i,temp_b1_9_7_r,temp_b1_9_7_i,temp_b1_9_8_r,temp_b1_9_8_i,temp_b1_10_7_r,temp_b1_10_7_i,temp_b1_10_8_r,temp_b1_10_8_i);
MULT MULT37 (clk,in_9_9_r,in_9_9_i,in_9_10_r,in_9_10_i,in_10_9_r,in_10_9_i,in_10_10_r,in_10_10_i,temp_m1_9_9_r,temp_m1_9_9_i,temp_m1_9_10_r,temp_m1_9_10_i,temp_m1_10_9_r,temp_m1_10_9_i,temp_m1_10_10_r,temp_m1_10_10_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly37 (clk,temp_m1_9_9_r,temp_m1_9_9_i,temp_m1_9_10_r,temp_m1_9_10_i,temp_m1_10_9_r,temp_m1_10_9_i,temp_m1_10_10_r,temp_m1_10_10_i,temp_b1_9_9_r,temp_b1_9_9_i,temp_b1_9_10_r,temp_b1_9_10_i,temp_b1_10_9_r,temp_b1_10_9_i,temp_b1_10_10_r,temp_b1_10_10_i);
MULT MULT38 (clk,in_9_11_r,in_9_11_i,in_9_12_r,in_9_12_i,in_10_11_r,in_10_11_i,in_10_12_r,in_10_12_i,temp_m1_9_11_r,temp_m1_9_11_i,temp_m1_9_12_r,temp_m1_9_12_i,temp_m1_10_11_r,temp_m1_10_11_i,temp_m1_10_12_r,temp_m1_10_12_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly38 (clk,temp_m1_9_11_r,temp_m1_9_11_i,temp_m1_9_12_r,temp_m1_9_12_i,temp_m1_10_11_r,temp_m1_10_11_i,temp_m1_10_12_r,temp_m1_10_12_i,temp_b1_9_11_r,temp_b1_9_11_i,temp_b1_9_12_r,temp_b1_9_12_i,temp_b1_10_11_r,temp_b1_10_11_i,temp_b1_10_12_r,temp_b1_10_12_i);
MULT MULT39 (clk,in_9_13_r,in_9_13_i,in_9_14_r,in_9_14_i,in_10_13_r,in_10_13_i,in_10_14_r,in_10_14_i,temp_m1_9_13_r,temp_m1_9_13_i,temp_m1_9_14_r,temp_m1_9_14_i,temp_m1_10_13_r,temp_m1_10_13_i,temp_m1_10_14_r,temp_m1_10_14_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly39 (clk,temp_m1_9_13_r,temp_m1_9_13_i,temp_m1_9_14_r,temp_m1_9_14_i,temp_m1_10_13_r,temp_m1_10_13_i,temp_m1_10_14_r,temp_m1_10_14_i,temp_b1_9_13_r,temp_b1_9_13_i,temp_b1_9_14_r,temp_b1_9_14_i,temp_b1_10_13_r,temp_b1_10_13_i,temp_b1_10_14_r,temp_b1_10_14_i);
MULT MULT40 (clk,in_9_15_r,in_9_15_i,in_9_16_r,in_9_16_i,in_10_15_r,in_10_15_i,in_10_16_r,in_10_16_i,temp_m1_9_15_r,temp_m1_9_15_i,temp_m1_9_16_r,temp_m1_9_16_i,temp_m1_10_15_r,temp_m1_10_15_i,temp_m1_10_16_r,temp_m1_10_16_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly40 (clk,temp_m1_9_15_r,temp_m1_9_15_i,temp_m1_9_16_r,temp_m1_9_16_i,temp_m1_10_15_r,temp_m1_10_15_i,temp_m1_10_16_r,temp_m1_10_16_i,temp_b1_9_15_r,temp_b1_9_15_i,temp_b1_9_16_r,temp_b1_9_16_i,temp_b1_10_15_r,temp_b1_10_15_i,temp_b1_10_16_r,temp_b1_10_16_i);
MULT MULT41 (clk,in_11_1_r,in_11_1_i,in_11_2_r,in_11_2_i,in_12_1_r,in_12_1_i,in_12_2_r,in_12_2_i,temp_m1_11_1_r,temp_m1_11_1_i,temp_m1_11_2_r,temp_m1_11_2_i,temp_m1_12_1_r,temp_m1_12_1_i,temp_m1_12_2_r,temp_m1_12_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly41 (clk,temp_m1_11_1_r,temp_m1_11_1_i,temp_m1_11_2_r,temp_m1_11_2_i,temp_m1_12_1_r,temp_m1_12_1_i,temp_m1_12_2_r,temp_m1_12_2_i,temp_b1_11_1_r,temp_b1_11_1_i,temp_b1_11_2_r,temp_b1_11_2_i,temp_b1_12_1_r,temp_b1_12_1_i,temp_b1_12_2_r,temp_b1_12_2_i);
MULT MULT42 (clk,in_11_3_r,in_11_3_i,in_11_4_r,in_11_4_i,in_12_3_r,in_12_3_i,in_12_4_r,in_12_4_i,temp_m1_11_3_r,temp_m1_11_3_i,temp_m1_11_4_r,temp_m1_11_4_i,temp_m1_12_3_r,temp_m1_12_3_i,temp_m1_12_4_r,temp_m1_12_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly42 (clk,temp_m1_11_3_r,temp_m1_11_3_i,temp_m1_11_4_r,temp_m1_11_4_i,temp_m1_12_3_r,temp_m1_12_3_i,temp_m1_12_4_r,temp_m1_12_4_i,temp_b1_11_3_r,temp_b1_11_3_i,temp_b1_11_4_r,temp_b1_11_4_i,temp_b1_12_3_r,temp_b1_12_3_i,temp_b1_12_4_r,temp_b1_12_4_i);
MULT MULT43 (clk,in_11_5_r,in_11_5_i,in_11_6_r,in_11_6_i,in_12_5_r,in_12_5_i,in_12_6_r,in_12_6_i,temp_m1_11_5_r,temp_m1_11_5_i,temp_m1_11_6_r,temp_m1_11_6_i,temp_m1_12_5_r,temp_m1_12_5_i,temp_m1_12_6_r,temp_m1_12_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly43 (clk,temp_m1_11_5_r,temp_m1_11_5_i,temp_m1_11_6_r,temp_m1_11_6_i,temp_m1_12_5_r,temp_m1_12_5_i,temp_m1_12_6_r,temp_m1_12_6_i,temp_b1_11_5_r,temp_b1_11_5_i,temp_b1_11_6_r,temp_b1_11_6_i,temp_b1_12_5_r,temp_b1_12_5_i,temp_b1_12_6_r,temp_b1_12_6_i);
MULT MULT44 (clk,in_11_7_r,in_11_7_i,in_11_8_r,in_11_8_i,in_12_7_r,in_12_7_i,in_12_8_r,in_12_8_i,temp_m1_11_7_r,temp_m1_11_7_i,temp_m1_11_8_r,temp_m1_11_8_i,temp_m1_12_7_r,temp_m1_12_7_i,temp_m1_12_8_r,temp_m1_12_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly44 (clk,temp_m1_11_7_r,temp_m1_11_7_i,temp_m1_11_8_r,temp_m1_11_8_i,temp_m1_12_7_r,temp_m1_12_7_i,temp_m1_12_8_r,temp_m1_12_8_i,temp_b1_11_7_r,temp_b1_11_7_i,temp_b1_11_8_r,temp_b1_11_8_i,temp_b1_12_7_r,temp_b1_12_7_i,temp_b1_12_8_r,temp_b1_12_8_i);
MULT MULT45 (clk,in_11_9_r,in_11_9_i,in_11_10_r,in_11_10_i,in_12_9_r,in_12_9_i,in_12_10_r,in_12_10_i,temp_m1_11_9_r,temp_m1_11_9_i,temp_m1_11_10_r,temp_m1_11_10_i,temp_m1_12_9_r,temp_m1_12_9_i,temp_m1_12_10_r,temp_m1_12_10_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly45 (clk,temp_m1_11_9_r,temp_m1_11_9_i,temp_m1_11_10_r,temp_m1_11_10_i,temp_m1_12_9_r,temp_m1_12_9_i,temp_m1_12_10_r,temp_m1_12_10_i,temp_b1_11_9_r,temp_b1_11_9_i,temp_b1_11_10_r,temp_b1_11_10_i,temp_b1_12_9_r,temp_b1_12_9_i,temp_b1_12_10_r,temp_b1_12_10_i);
MULT MULT46 (clk,in_11_11_r,in_11_11_i,in_11_12_r,in_11_12_i,in_12_11_r,in_12_11_i,in_12_12_r,in_12_12_i,temp_m1_11_11_r,temp_m1_11_11_i,temp_m1_11_12_r,temp_m1_11_12_i,temp_m1_12_11_r,temp_m1_12_11_i,temp_m1_12_12_r,temp_m1_12_12_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly46 (clk,temp_m1_11_11_r,temp_m1_11_11_i,temp_m1_11_12_r,temp_m1_11_12_i,temp_m1_12_11_r,temp_m1_12_11_i,temp_m1_12_12_r,temp_m1_12_12_i,temp_b1_11_11_r,temp_b1_11_11_i,temp_b1_11_12_r,temp_b1_11_12_i,temp_b1_12_11_r,temp_b1_12_11_i,temp_b1_12_12_r,temp_b1_12_12_i);
MULT MULT47 (clk,in_11_13_r,in_11_13_i,in_11_14_r,in_11_14_i,in_12_13_r,in_12_13_i,in_12_14_r,in_12_14_i,temp_m1_11_13_r,temp_m1_11_13_i,temp_m1_11_14_r,temp_m1_11_14_i,temp_m1_12_13_r,temp_m1_12_13_i,temp_m1_12_14_r,temp_m1_12_14_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly47 (clk,temp_m1_11_13_r,temp_m1_11_13_i,temp_m1_11_14_r,temp_m1_11_14_i,temp_m1_12_13_r,temp_m1_12_13_i,temp_m1_12_14_r,temp_m1_12_14_i,temp_b1_11_13_r,temp_b1_11_13_i,temp_b1_11_14_r,temp_b1_11_14_i,temp_b1_12_13_r,temp_b1_12_13_i,temp_b1_12_14_r,temp_b1_12_14_i);
MULT MULT48 (clk,in_11_15_r,in_11_15_i,in_11_16_r,in_11_16_i,in_12_15_r,in_12_15_i,in_12_16_r,in_12_16_i,temp_m1_11_15_r,temp_m1_11_15_i,temp_m1_11_16_r,temp_m1_11_16_i,temp_m1_12_15_r,temp_m1_12_15_i,temp_m1_12_16_r,temp_m1_12_16_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly48 (clk,temp_m1_11_15_r,temp_m1_11_15_i,temp_m1_11_16_r,temp_m1_11_16_i,temp_m1_12_15_r,temp_m1_12_15_i,temp_m1_12_16_r,temp_m1_12_16_i,temp_b1_11_15_r,temp_b1_11_15_i,temp_b1_11_16_r,temp_b1_11_16_i,temp_b1_12_15_r,temp_b1_12_15_i,temp_b1_12_16_r,temp_b1_12_16_i);
MULT MULT49 (clk,in_13_1_r,in_13_1_i,in_13_2_r,in_13_2_i,in_14_1_r,in_14_1_i,in_14_2_r,in_14_2_i,temp_m1_13_1_r,temp_m1_13_1_i,temp_m1_13_2_r,temp_m1_13_2_i,temp_m1_14_1_r,temp_m1_14_1_i,temp_m1_14_2_r,temp_m1_14_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly49 (clk,temp_m1_13_1_r,temp_m1_13_1_i,temp_m1_13_2_r,temp_m1_13_2_i,temp_m1_14_1_r,temp_m1_14_1_i,temp_m1_14_2_r,temp_m1_14_2_i,temp_b1_13_1_r,temp_b1_13_1_i,temp_b1_13_2_r,temp_b1_13_2_i,temp_b1_14_1_r,temp_b1_14_1_i,temp_b1_14_2_r,temp_b1_14_2_i);
MULT MULT50 (clk,in_13_3_r,in_13_3_i,in_13_4_r,in_13_4_i,in_14_3_r,in_14_3_i,in_14_4_r,in_14_4_i,temp_m1_13_3_r,temp_m1_13_3_i,temp_m1_13_4_r,temp_m1_13_4_i,temp_m1_14_3_r,temp_m1_14_3_i,temp_m1_14_4_r,temp_m1_14_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly50 (clk,temp_m1_13_3_r,temp_m1_13_3_i,temp_m1_13_4_r,temp_m1_13_4_i,temp_m1_14_3_r,temp_m1_14_3_i,temp_m1_14_4_r,temp_m1_14_4_i,temp_b1_13_3_r,temp_b1_13_3_i,temp_b1_13_4_r,temp_b1_13_4_i,temp_b1_14_3_r,temp_b1_14_3_i,temp_b1_14_4_r,temp_b1_14_4_i);
MULT MULT51 (clk,in_13_5_r,in_13_5_i,in_13_6_r,in_13_6_i,in_14_5_r,in_14_5_i,in_14_6_r,in_14_6_i,temp_m1_13_5_r,temp_m1_13_5_i,temp_m1_13_6_r,temp_m1_13_6_i,temp_m1_14_5_r,temp_m1_14_5_i,temp_m1_14_6_r,temp_m1_14_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly51 (clk,temp_m1_13_5_r,temp_m1_13_5_i,temp_m1_13_6_r,temp_m1_13_6_i,temp_m1_14_5_r,temp_m1_14_5_i,temp_m1_14_6_r,temp_m1_14_6_i,temp_b1_13_5_r,temp_b1_13_5_i,temp_b1_13_6_r,temp_b1_13_6_i,temp_b1_14_5_r,temp_b1_14_5_i,temp_b1_14_6_r,temp_b1_14_6_i);
MULT MULT52 (clk,in_13_7_r,in_13_7_i,in_13_8_r,in_13_8_i,in_14_7_r,in_14_7_i,in_14_8_r,in_14_8_i,temp_m1_13_7_r,temp_m1_13_7_i,temp_m1_13_8_r,temp_m1_13_8_i,temp_m1_14_7_r,temp_m1_14_7_i,temp_m1_14_8_r,temp_m1_14_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly52 (clk,temp_m1_13_7_r,temp_m1_13_7_i,temp_m1_13_8_r,temp_m1_13_8_i,temp_m1_14_7_r,temp_m1_14_7_i,temp_m1_14_8_r,temp_m1_14_8_i,temp_b1_13_7_r,temp_b1_13_7_i,temp_b1_13_8_r,temp_b1_13_8_i,temp_b1_14_7_r,temp_b1_14_7_i,temp_b1_14_8_r,temp_b1_14_8_i);
MULT MULT53 (clk,in_13_9_r,in_13_9_i,in_13_10_r,in_13_10_i,in_14_9_r,in_14_9_i,in_14_10_r,in_14_10_i,temp_m1_13_9_r,temp_m1_13_9_i,temp_m1_13_10_r,temp_m1_13_10_i,temp_m1_14_9_r,temp_m1_14_9_i,temp_m1_14_10_r,temp_m1_14_10_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly53 (clk,temp_m1_13_9_r,temp_m1_13_9_i,temp_m1_13_10_r,temp_m1_13_10_i,temp_m1_14_9_r,temp_m1_14_9_i,temp_m1_14_10_r,temp_m1_14_10_i,temp_b1_13_9_r,temp_b1_13_9_i,temp_b1_13_10_r,temp_b1_13_10_i,temp_b1_14_9_r,temp_b1_14_9_i,temp_b1_14_10_r,temp_b1_14_10_i);
MULT MULT54 (clk,in_13_11_r,in_13_11_i,in_13_12_r,in_13_12_i,in_14_11_r,in_14_11_i,in_14_12_r,in_14_12_i,temp_m1_13_11_r,temp_m1_13_11_i,temp_m1_13_12_r,temp_m1_13_12_i,temp_m1_14_11_r,temp_m1_14_11_i,temp_m1_14_12_r,temp_m1_14_12_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly54 (clk,temp_m1_13_11_r,temp_m1_13_11_i,temp_m1_13_12_r,temp_m1_13_12_i,temp_m1_14_11_r,temp_m1_14_11_i,temp_m1_14_12_r,temp_m1_14_12_i,temp_b1_13_11_r,temp_b1_13_11_i,temp_b1_13_12_r,temp_b1_13_12_i,temp_b1_14_11_r,temp_b1_14_11_i,temp_b1_14_12_r,temp_b1_14_12_i);
MULT MULT55 (clk,in_13_13_r,in_13_13_i,in_13_14_r,in_13_14_i,in_14_13_r,in_14_13_i,in_14_14_r,in_14_14_i,temp_m1_13_13_r,temp_m1_13_13_i,temp_m1_13_14_r,temp_m1_13_14_i,temp_m1_14_13_r,temp_m1_14_13_i,temp_m1_14_14_r,temp_m1_14_14_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly55 (clk,temp_m1_13_13_r,temp_m1_13_13_i,temp_m1_13_14_r,temp_m1_13_14_i,temp_m1_14_13_r,temp_m1_14_13_i,temp_m1_14_14_r,temp_m1_14_14_i,temp_b1_13_13_r,temp_b1_13_13_i,temp_b1_13_14_r,temp_b1_13_14_i,temp_b1_14_13_r,temp_b1_14_13_i,temp_b1_14_14_r,temp_b1_14_14_i);
MULT MULT56 (clk,in_13_15_r,in_13_15_i,in_13_16_r,in_13_16_i,in_14_15_r,in_14_15_i,in_14_16_r,in_14_16_i,temp_m1_13_15_r,temp_m1_13_15_i,temp_m1_13_16_r,temp_m1_13_16_i,temp_m1_14_15_r,temp_m1_14_15_i,temp_m1_14_16_r,temp_m1_14_16_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly56 (clk,temp_m1_13_15_r,temp_m1_13_15_i,temp_m1_13_16_r,temp_m1_13_16_i,temp_m1_14_15_r,temp_m1_14_15_i,temp_m1_14_16_r,temp_m1_14_16_i,temp_b1_13_15_r,temp_b1_13_15_i,temp_b1_13_16_r,temp_b1_13_16_i,temp_b1_14_15_r,temp_b1_14_15_i,temp_b1_14_16_r,temp_b1_14_16_i);
MULT MULT57 (clk,in_15_1_r,in_15_1_i,in_15_2_r,in_15_2_i,in_16_1_r,in_16_1_i,in_16_2_r,in_16_2_i,temp_m1_15_1_r,temp_m1_15_1_i,temp_m1_15_2_r,temp_m1_15_2_i,temp_m1_16_1_r,temp_m1_16_1_i,temp_m1_16_2_r,temp_m1_16_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly57 (clk,temp_m1_15_1_r,temp_m1_15_1_i,temp_m1_15_2_r,temp_m1_15_2_i,temp_m1_16_1_r,temp_m1_16_1_i,temp_m1_16_2_r,temp_m1_16_2_i,temp_b1_15_1_r,temp_b1_15_1_i,temp_b1_15_2_r,temp_b1_15_2_i,temp_b1_16_1_r,temp_b1_16_1_i,temp_b1_16_2_r,temp_b1_16_2_i);
MULT MULT58 (clk,in_15_3_r,in_15_3_i,in_15_4_r,in_15_4_i,in_16_3_r,in_16_3_i,in_16_4_r,in_16_4_i,temp_m1_15_3_r,temp_m1_15_3_i,temp_m1_15_4_r,temp_m1_15_4_i,temp_m1_16_3_r,temp_m1_16_3_i,temp_m1_16_4_r,temp_m1_16_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly58 (clk,temp_m1_15_3_r,temp_m1_15_3_i,temp_m1_15_4_r,temp_m1_15_4_i,temp_m1_16_3_r,temp_m1_16_3_i,temp_m1_16_4_r,temp_m1_16_4_i,temp_b1_15_3_r,temp_b1_15_3_i,temp_b1_15_4_r,temp_b1_15_4_i,temp_b1_16_3_r,temp_b1_16_3_i,temp_b1_16_4_r,temp_b1_16_4_i);
MULT MULT59 (clk,in_15_5_r,in_15_5_i,in_15_6_r,in_15_6_i,in_16_5_r,in_16_5_i,in_16_6_r,in_16_6_i,temp_m1_15_5_r,temp_m1_15_5_i,temp_m1_15_6_r,temp_m1_15_6_i,temp_m1_16_5_r,temp_m1_16_5_i,temp_m1_16_6_r,temp_m1_16_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly59 (clk,temp_m1_15_5_r,temp_m1_15_5_i,temp_m1_15_6_r,temp_m1_15_6_i,temp_m1_16_5_r,temp_m1_16_5_i,temp_m1_16_6_r,temp_m1_16_6_i,temp_b1_15_5_r,temp_b1_15_5_i,temp_b1_15_6_r,temp_b1_15_6_i,temp_b1_16_5_r,temp_b1_16_5_i,temp_b1_16_6_r,temp_b1_16_6_i);
MULT MULT60 (clk,in_15_7_r,in_15_7_i,in_15_8_r,in_15_8_i,in_16_7_r,in_16_7_i,in_16_8_r,in_16_8_i,temp_m1_15_7_r,temp_m1_15_7_i,temp_m1_15_8_r,temp_m1_15_8_i,temp_m1_16_7_r,temp_m1_16_7_i,temp_m1_16_8_r,temp_m1_16_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly60 (clk,temp_m1_15_7_r,temp_m1_15_7_i,temp_m1_15_8_r,temp_m1_15_8_i,temp_m1_16_7_r,temp_m1_16_7_i,temp_m1_16_8_r,temp_m1_16_8_i,temp_b1_15_7_r,temp_b1_15_7_i,temp_b1_15_8_r,temp_b1_15_8_i,temp_b1_16_7_r,temp_b1_16_7_i,temp_b1_16_8_r,temp_b1_16_8_i);
MULT MULT61 (clk,in_15_9_r,in_15_9_i,in_15_10_r,in_15_10_i,in_16_9_r,in_16_9_i,in_16_10_r,in_16_10_i,temp_m1_15_9_r,temp_m1_15_9_i,temp_m1_15_10_r,temp_m1_15_10_i,temp_m1_16_9_r,temp_m1_16_9_i,temp_m1_16_10_r,temp_m1_16_10_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly61 (clk,temp_m1_15_9_r,temp_m1_15_9_i,temp_m1_15_10_r,temp_m1_15_10_i,temp_m1_16_9_r,temp_m1_16_9_i,temp_m1_16_10_r,temp_m1_16_10_i,temp_b1_15_9_r,temp_b1_15_9_i,temp_b1_15_10_r,temp_b1_15_10_i,temp_b1_16_9_r,temp_b1_16_9_i,temp_b1_16_10_r,temp_b1_16_10_i);
MULT MULT62 (clk,in_15_11_r,in_15_11_i,in_15_12_r,in_15_12_i,in_16_11_r,in_16_11_i,in_16_12_r,in_16_12_i,temp_m1_15_11_r,temp_m1_15_11_i,temp_m1_15_12_r,temp_m1_15_12_i,temp_m1_16_11_r,temp_m1_16_11_i,temp_m1_16_12_r,temp_m1_16_12_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly62 (clk,temp_m1_15_11_r,temp_m1_15_11_i,temp_m1_15_12_r,temp_m1_15_12_i,temp_m1_16_11_r,temp_m1_16_11_i,temp_m1_16_12_r,temp_m1_16_12_i,temp_b1_15_11_r,temp_b1_15_11_i,temp_b1_15_12_r,temp_b1_15_12_i,temp_b1_16_11_r,temp_b1_16_11_i,temp_b1_16_12_r,temp_b1_16_12_i);
MULT MULT63 (clk,in_15_13_r,in_15_13_i,in_15_14_r,in_15_14_i,in_16_13_r,in_16_13_i,in_16_14_r,in_16_14_i,temp_m1_15_13_r,temp_m1_15_13_i,temp_m1_15_14_r,temp_m1_15_14_i,temp_m1_16_13_r,temp_m1_16_13_i,temp_m1_16_14_r,temp_m1_16_14_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly63 (clk,temp_m1_15_13_r,temp_m1_15_13_i,temp_m1_15_14_r,temp_m1_15_14_i,temp_m1_16_13_r,temp_m1_16_13_i,temp_m1_16_14_r,temp_m1_16_14_i,temp_b1_15_13_r,temp_b1_15_13_i,temp_b1_15_14_r,temp_b1_15_14_i,temp_b1_16_13_r,temp_b1_16_13_i,temp_b1_16_14_r,temp_b1_16_14_i);
MULT MULT64 (clk,in_15_15_r,in_15_15_i,in_15_16_r,in_15_16_i,in_16_15_r,in_16_15_i,in_16_16_r,in_16_16_i,temp_m1_15_15_r,temp_m1_15_15_i,temp_m1_15_16_r,temp_m1_15_16_i,temp_m1_16_15_r,temp_m1_16_15_i,temp_m1_16_16_r,temp_m1_16_16_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly64 (clk,temp_m1_15_15_r,temp_m1_15_15_i,temp_m1_15_16_r,temp_m1_15_16_i,temp_m1_16_15_r,temp_m1_16_15_i,temp_m1_16_16_r,temp_m1_16_16_i,temp_b1_15_15_r,temp_b1_15_15_i,temp_b1_15_16_r,temp_b1_15_16_i,temp_b1_16_15_r,temp_b1_16_15_i,temp_b1_16_16_r,temp_b1_16_16_i);
MULT MULT65 (clk,temp_b1_1_1_r,temp_b1_1_1_i,temp_b1_1_3_r,temp_b1_1_3_i,temp_b1_3_1_r,temp_b1_3_1_i,temp_b1_3_3_r,temp_b1_3_3_i,temp_m2_1_1_r,temp_m2_1_1_i,temp_m2_1_3_r,temp_m2_1_3_i,temp_m2_3_1_r,temp_m2_3_1_i,temp_m2_3_3_r,temp_m2_3_3_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly65 (clk,temp_m2_1_1_r,temp_m2_1_1_i,temp_m2_1_3_r,temp_m2_1_3_i,temp_m2_3_1_r,temp_m2_3_1_i,temp_m2_3_3_r,temp_m2_3_3_i,temp_b2_1_1_r,temp_b2_1_1_i,temp_b2_1_3_r,temp_b2_1_3_i,temp_b2_3_1_r,temp_b2_3_1_i,temp_b2_3_3_r,temp_b2_3_3_i);
MULT MULT66 (clk,temp_b1_1_2_r,temp_b1_1_2_i,temp_b1_1_4_r,temp_b1_1_4_i,temp_b1_3_2_r,temp_b1_3_2_i,temp_b1_3_4_r,temp_b1_3_4_i,temp_m2_1_2_r,temp_m2_1_2_i,temp_m2_1_4_r,temp_m2_1_4_i,temp_m2_3_2_r,temp_m2_3_2_i,temp_m2_3_4_r,temp_m2_3_4_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly66 (clk,temp_m2_1_2_r,temp_m2_1_2_i,temp_m2_1_4_r,temp_m2_1_4_i,temp_m2_3_2_r,temp_m2_3_2_i,temp_m2_3_4_r,temp_m2_3_4_i,temp_b2_1_2_r,temp_b2_1_2_i,temp_b2_1_4_r,temp_b2_1_4_i,temp_b2_3_2_r,temp_b2_3_2_i,temp_b2_3_4_r,temp_b2_3_4_i);
MULT MULT67 (clk,temp_b1_2_1_r,temp_b1_2_1_i,temp_b1_2_3_r,temp_b1_2_3_i,temp_b1_4_1_r,temp_b1_4_1_i,temp_b1_4_3_r,temp_b1_4_3_i,temp_m2_2_1_r,temp_m2_2_1_i,temp_m2_2_3_r,temp_m2_2_3_i,temp_m2_4_1_r,temp_m2_4_1_i,temp_m2_4_3_r,temp_m2_4_3_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly67 (clk,temp_m2_2_1_r,temp_m2_2_1_i,temp_m2_2_3_r,temp_m2_2_3_i,temp_m2_4_1_r,temp_m2_4_1_i,temp_m2_4_3_r,temp_m2_4_3_i,temp_b2_2_1_r,temp_b2_2_1_i,temp_b2_2_3_r,temp_b2_2_3_i,temp_b2_4_1_r,temp_b2_4_1_i,temp_b2_4_3_r,temp_b2_4_3_i);
MULT MULT68 (clk,temp_b1_2_2_r,temp_b1_2_2_i,temp_b1_2_4_r,temp_b1_2_4_i,temp_b1_4_2_r,temp_b1_4_2_i,temp_b1_4_4_r,temp_b1_4_4_i,temp_m2_2_2_r,temp_m2_2_2_i,temp_m2_2_4_r,temp_m2_2_4_i,temp_m2_4_2_r,temp_m2_4_2_i,temp_m2_4_4_r,temp_m2_4_4_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly68 (clk,temp_m2_2_2_r,temp_m2_2_2_i,temp_m2_2_4_r,temp_m2_2_4_i,temp_m2_4_2_r,temp_m2_4_2_i,temp_m2_4_4_r,temp_m2_4_4_i,temp_b2_2_2_r,temp_b2_2_2_i,temp_b2_2_4_r,temp_b2_2_4_i,temp_b2_4_2_r,temp_b2_4_2_i,temp_b2_4_4_r,temp_b2_4_4_i);
MULT MULT69 (clk,temp_b1_1_5_r,temp_b1_1_5_i,temp_b1_1_7_r,temp_b1_1_7_i,temp_b1_3_5_r,temp_b1_3_5_i,temp_b1_3_7_r,temp_b1_3_7_i,temp_m2_1_5_r,temp_m2_1_5_i,temp_m2_1_7_r,temp_m2_1_7_i,temp_m2_3_5_r,temp_m2_3_5_i,temp_m2_3_7_r,temp_m2_3_7_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly69 (clk,temp_m2_1_5_r,temp_m2_1_5_i,temp_m2_1_7_r,temp_m2_1_7_i,temp_m2_3_5_r,temp_m2_3_5_i,temp_m2_3_7_r,temp_m2_3_7_i,temp_b2_1_5_r,temp_b2_1_5_i,temp_b2_1_7_r,temp_b2_1_7_i,temp_b2_3_5_r,temp_b2_3_5_i,temp_b2_3_7_r,temp_b2_3_7_i);
MULT MULT70 (clk,temp_b1_1_6_r,temp_b1_1_6_i,temp_b1_1_8_r,temp_b1_1_8_i,temp_b1_3_6_r,temp_b1_3_6_i,temp_b1_3_8_r,temp_b1_3_8_i,temp_m2_1_6_r,temp_m2_1_6_i,temp_m2_1_8_r,temp_m2_1_8_i,temp_m2_3_6_r,temp_m2_3_6_i,temp_m2_3_8_r,temp_m2_3_8_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly70 (clk,temp_m2_1_6_r,temp_m2_1_6_i,temp_m2_1_8_r,temp_m2_1_8_i,temp_m2_3_6_r,temp_m2_3_6_i,temp_m2_3_8_r,temp_m2_3_8_i,temp_b2_1_6_r,temp_b2_1_6_i,temp_b2_1_8_r,temp_b2_1_8_i,temp_b2_3_6_r,temp_b2_3_6_i,temp_b2_3_8_r,temp_b2_3_8_i);
MULT MULT71 (clk,temp_b1_2_5_r,temp_b1_2_5_i,temp_b1_2_7_r,temp_b1_2_7_i,temp_b1_4_5_r,temp_b1_4_5_i,temp_b1_4_7_r,temp_b1_4_7_i,temp_m2_2_5_r,temp_m2_2_5_i,temp_m2_2_7_r,temp_m2_2_7_i,temp_m2_4_5_r,temp_m2_4_5_i,temp_m2_4_7_r,temp_m2_4_7_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly71 (clk,temp_m2_2_5_r,temp_m2_2_5_i,temp_m2_2_7_r,temp_m2_2_7_i,temp_m2_4_5_r,temp_m2_4_5_i,temp_m2_4_7_r,temp_m2_4_7_i,temp_b2_2_5_r,temp_b2_2_5_i,temp_b2_2_7_r,temp_b2_2_7_i,temp_b2_4_5_r,temp_b2_4_5_i,temp_b2_4_7_r,temp_b2_4_7_i);
MULT MULT72 (clk,temp_b1_2_6_r,temp_b1_2_6_i,temp_b1_2_8_r,temp_b1_2_8_i,temp_b1_4_6_r,temp_b1_4_6_i,temp_b1_4_8_r,temp_b1_4_8_i,temp_m2_2_6_r,temp_m2_2_6_i,temp_m2_2_8_r,temp_m2_2_8_i,temp_m2_4_6_r,temp_m2_4_6_i,temp_m2_4_8_r,temp_m2_4_8_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly72 (clk,temp_m2_2_6_r,temp_m2_2_6_i,temp_m2_2_8_r,temp_m2_2_8_i,temp_m2_4_6_r,temp_m2_4_6_i,temp_m2_4_8_r,temp_m2_4_8_i,temp_b2_2_6_r,temp_b2_2_6_i,temp_b2_2_8_r,temp_b2_2_8_i,temp_b2_4_6_r,temp_b2_4_6_i,temp_b2_4_8_r,temp_b2_4_8_i);
MULT MULT73 (clk,temp_b1_1_9_r,temp_b1_1_9_i,temp_b1_1_11_r,temp_b1_1_11_i,temp_b1_3_9_r,temp_b1_3_9_i,temp_b1_3_11_r,temp_b1_3_11_i,temp_m2_1_9_r,temp_m2_1_9_i,temp_m2_1_11_r,temp_m2_1_11_i,temp_m2_3_9_r,temp_m2_3_9_i,temp_m2_3_11_r,temp_m2_3_11_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly73 (clk,temp_m2_1_9_r,temp_m2_1_9_i,temp_m2_1_11_r,temp_m2_1_11_i,temp_m2_3_9_r,temp_m2_3_9_i,temp_m2_3_11_r,temp_m2_3_11_i,temp_b2_1_9_r,temp_b2_1_9_i,temp_b2_1_11_r,temp_b2_1_11_i,temp_b2_3_9_r,temp_b2_3_9_i,temp_b2_3_11_r,temp_b2_3_11_i);
MULT MULT74 (clk,temp_b1_1_10_r,temp_b1_1_10_i,temp_b1_1_12_r,temp_b1_1_12_i,temp_b1_3_10_r,temp_b1_3_10_i,temp_b1_3_12_r,temp_b1_3_12_i,temp_m2_1_10_r,temp_m2_1_10_i,temp_m2_1_12_r,temp_m2_1_12_i,temp_m2_3_10_r,temp_m2_3_10_i,temp_m2_3_12_r,temp_m2_3_12_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly74 (clk,temp_m2_1_10_r,temp_m2_1_10_i,temp_m2_1_12_r,temp_m2_1_12_i,temp_m2_3_10_r,temp_m2_3_10_i,temp_m2_3_12_r,temp_m2_3_12_i,temp_b2_1_10_r,temp_b2_1_10_i,temp_b2_1_12_r,temp_b2_1_12_i,temp_b2_3_10_r,temp_b2_3_10_i,temp_b2_3_12_r,temp_b2_3_12_i);
MULT MULT75 (clk,temp_b1_2_9_r,temp_b1_2_9_i,temp_b1_2_11_r,temp_b1_2_11_i,temp_b1_4_9_r,temp_b1_4_9_i,temp_b1_4_11_r,temp_b1_4_11_i,temp_m2_2_9_r,temp_m2_2_9_i,temp_m2_2_11_r,temp_m2_2_11_i,temp_m2_4_9_r,temp_m2_4_9_i,temp_m2_4_11_r,temp_m2_4_11_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly75 (clk,temp_m2_2_9_r,temp_m2_2_9_i,temp_m2_2_11_r,temp_m2_2_11_i,temp_m2_4_9_r,temp_m2_4_9_i,temp_m2_4_11_r,temp_m2_4_11_i,temp_b2_2_9_r,temp_b2_2_9_i,temp_b2_2_11_r,temp_b2_2_11_i,temp_b2_4_9_r,temp_b2_4_9_i,temp_b2_4_11_r,temp_b2_4_11_i);
MULT MULT76 (clk,temp_b1_2_10_r,temp_b1_2_10_i,temp_b1_2_12_r,temp_b1_2_12_i,temp_b1_4_10_r,temp_b1_4_10_i,temp_b1_4_12_r,temp_b1_4_12_i,temp_m2_2_10_r,temp_m2_2_10_i,temp_m2_2_12_r,temp_m2_2_12_i,temp_m2_4_10_r,temp_m2_4_10_i,temp_m2_4_12_r,temp_m2_4_12_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly76 (clk,temp_m2_2_10_r,temp_m2_2_10_i,temp_m2_2_12_r,temp_m2_2_12_i,temp_m2_4_10_r,temp_m2_4_10_i,temp_m2_4_12_r,temp_m2_4_12_i,temp_b2_2_10_r,temp_b2_2_10_i,temp_b2_2_12_r,temp_b2_2_12_i,temp_b2_4_10_r,temp_b2_4_10_i,temp_b2_4_12_r,temp_b2_4_12_i);
MULT MULT77 (clk,temp_b1_1_13_r,temp_b1_1_13_i,temp_b1_1_15_r,temp_b1_1_15_i,temp_b1_3_13_r,temp_b1_3_13_i,temp_b1_3_15_r,temp_b1_3_15_i,temp_m2_1_13_r,temp_m2_1_13_i,temp_m2_1_15_r,temp_m2_1_15_i,temp_m2_3_13_r,temp_m2_3_13_i,temp_m2_3_15_r,temp_m2_3_15_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly77 (clk,temp_m2_1_13_r,temp_m2_1_13_i,temp_m2_1_15_r,temp_m2_1_15_i,temp_m2_3_13_r,temp_m2_3_13_i,temp_m2_3_15_r,temp_m2_3_15_i,temp_b2_1_13_r,temp_b2_1_13_i,temp_b2_1_15_r,temp_b2_1_15_i,temp_b2_3_13_r,temp_b2_3_13_i,temp_b2_3_15_r,temp_b2_3_15_i);
MULT MULT78 (clk,temp_b1_1_14_r,temp_b1_1_14_i,temp_b1_1_16_r,temp_b1_1_16_i,temp_b1_3_14_r,temp_b1_3_14_i,temp_b1_3_16_r,temp_b1_3_16_i,temp_m2_1_14_r,temp_m2_1_14_i,temp_m2_1_16_r,temp_m2_1_16_i,temp_m2_3_14_r,temp_m2_3_14_i,temp_m2_3_16_r,temp_m2_3_16_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly78 (clk,temp_m2_1_14_r,temp_m2_1_14_i,temp_m2_1_16_r,temp_m2_1_16_i,temp_m2_3_14_r,temp_m2_3_14_i,temp_m2_3_16_r,temp_m2_3_16_i,temp_b2_1_14_r,temp_b2_1_14_i,temp_b2_1_16_r,temp_b2_1_16_i,temp_b2_3_14_r,temp_b2_3_14_i,temp_b2_3_16_r,temp_b2_3_16_i);
MULT MULT79 (clk,temp_b1_2_13_r,temp_b1_2_13_i,temp_b1_2_15_r,temp_b1_2_15_i,temp_b1_4_13_r,temp_b1_4_13_i,temp_b1_4_15_r,temp_b1_4_15_i,temp_m2_2_13_r,temp_m2_2_13_i,temp_m2_2_15_r,temp_m2_2_15_i,temp_m2_4_13_r,temp_m2_4_13_i,temp_m2_4_15_r,temp_m2_4_15_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly79 (clk,temp_m2_2_13_r,temp_m2_2_13_i,temp_m2_2_15_r,temp_m2_2_15_i,temp_m2_4_13_r,temp_m2_4_13_i,temp_m2_4_15_r,temp_m2_4_15_i,temp_b2_2_13_r,temp_b2_2_13_i,temp_b2_2_15_r,temp_b2_2_15_i,temp_b2_4_13_r,temp_b2_4_13_i,temp_b2_4_15_r,temp_b2_4_15_i);
MULT MULT80 (clk,temp_b1_2_14_r,temp_b1_2_14_i,temp_b1_2_16_r,temp_b1_2_16_i,temp_b1_4_14_r,temp_b1_4_14_i,temp_b1_4_16_r,temp_b1_4_16_i,temp_m2_2_14_r,temp_m2_2_14_i,temp_m2_2_16_r,temp_m2_2_16_i,temp_m2_4_14_r,temp_m2_4_14_i,temp_m2_4_16_r,temp_m2_4_16_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly80 (clk,temp_m2_2_14_r,temp_m2_2_14_i,temp_m2_2_16_r,temp_m2_2_16_i,temp_m2_4_14_r,temp_m2_4_14_i,temp_m2_4_16_r,temp_m2_4_16_i,temp_b2_2_14_r,temp_b2_2_14_i,temp_b2_2_16_r,temp_b2_2_16_i,temp_b2_4_14_r,temp_b2_4_14_i,temp_b2_4_16_r,temp_b2_4_16_i);
MULT MULT81 (clk,temp_b1_5_1_r,temp_b1_5_1_i,temp_b1_5_3_r,temp_b1_5_3_i,temp_b1_7_1_r,temp_b1_7_1_i,temp_b1_7_3_r,temp_b1_7_3_i,temp_m2_5_1_r,temp_m2_5_1_i,temp_m2_5_3_r,temp_m2_5_3_i,temp_m2_7_1_r,temp_m2_7_1_i,temp_m2_7_3_r,temp_m2_7_3_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly81 (clk,temp_m2_5_1_r,temp_m2_5_1_i,temp_m2_5_3_r,temp_m2_5_3_i,temp_m2_7_1_r,temp_m2_7_1_i,temp_m2_7_3_r,temp_m2_7_3_i,temp_b2_5_1_r,temp_b2_5_1_i,temp_b2_5_3_r,temp_b2_5_3_i,temp_b2_7_1_r,temp_b2_7_1_i,temp_b2_7_3_r,temp_b2_7_3_i);
MULT MULT82 (clk,temp_b1_5_2_r,temp_b1_5_2_i,temp_b1_5_4_r,temp_b1_5_4_i,temp_b1_7_2_r,temp_b1_7_2_i,temp_b1_7_4_r,temp_b1_7_4_i,temp_m2_5_2_r,temp_m2_5_2_i,temp_m2_5_4_r,temp_m2_5_4_i,temp_m2_7_2_r,temp_m2_7_2_i,temp_m2_7_4_r,temp_m2_7_4_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly82 (clk,temp_m2_5_2_r,temp_m2_5_2_i,temp_m2_5_4_r,temp_m2_5_4_i,temp_m2_7_2_r,temp_m2_7_2_i,temp_m2_7_4_r,temp_m2_7_4_i,temp_b2_5_2_r,temp_b2_5_2_i,temp_b2_5_4_r,temp_b2_5_4_i,temp_b2_7_2_r,temp_b2_7_2_i,temp_b2_7_4_r,temp_b2_7_4_i);
MULT MULT83 (clk,temp_b1_6_1_r,temp_b1_6_1_i,temp_b1_6_3_r,temp_b1_6_3_i,temp_b1_8_1_r,temp_b1_8_1_i,temp_b1_8_3_r,temp_b1_8_3_i,temp_m2_6_1_r,temp_m2_6_1_i,temp_m2_6_3_r,temp_m2_6_3_i,temp_m2_8_1_r,temp_m2_8_1_i,temp_m2_8_3_r,temp_m2_8_3_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly83 (clk,temp_m2_6_1_r,temp_m2_6_1_i,temp_m2_6_3_r,temp_m2_6_3_i,temp_m2_8_1_r,temp_m2_8_1_i,temp_m2_8_3_r,temp_m2_8_3_i,temp_b2_6_1_r,temp_b2_6_1_i,temp_b2_6_3_r,temp_b2_6_3_i,temp_b2_8_1_r,temp_b2_8_1_i,temp_b2_8_3_r,temp_b2_8_3_i);
MULT MULT84 (clk,temp_b1_6_2_r,temp_b1_6_2_i,temp_b1_6_4_r,temp_b1_6_4_i,temp_b1_8_2_r,temp_b1_8_2_i,temp_b1_8_4_r,temp_b1_8_4_i,temp_m2_6_2_r,temp_m2_6_2_i,temp_m2_6_4_r,temp_m2_6_4_i,temp_m2_8_2_r,temp_m2_8_2_i,temp_m2_8_4_r,temp_m2_8_4_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly84 (clk,temp_m2_6_2_r,temp_m2_6_2_i,temp_m2_6_4_r,temp_m2_6_4_i,temp_m2_8_2_r,temp_m2_8_2_i,temp_m2_8_4_r,temp_m2_8_4_i,temp_b2_6_2_r,temp_b2_6_2_i,temp_b2_6_4_r,temp_b2_6_4_i,temp_b2_8_2_r,temp_b2_8_2_i,temp_b2_8_4_r,temp_b2_8_4_i);
MULT MULT85 (clk,temp_b1_5_5_r,temp_b1_5_5_i,temp_b1_5_7_r,temp_b1_5_7_i,temp_b1_7_5_r,temp_b1_7_5_i,temp_b1_7_7_r,temp_b1_7_7_i,temp_m2_5_5_r,temp_m2_5_5_i,temp_m2_5_7_r,temp_m2_5_7_i,temp_m2_7_5_r,temp_m2_7_5_i,temp_m2_7_7_r,temp_m2_7_7_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly85 (clk,temp_m2_5_5_r,temp_m2_5_5_i,temp_m2_5_7_r,temp_m2_5_7_i,temp_m2_7_5_r,temp_m2_7_5_i,temp_m2_7_7_r,temp_m2_7_7_i,temp_b2_5_5_r,temp_b2_5_5_i,temp_b2_5_7_r,temp_b2_5_7_i,temp_b2_7_5_r,temp_b2_7_5_i,temp_b2_7_7_r,temp_b2_7_7_i);
MULT MULT86 (clk,temp_b1_5_6_r,temp_b1_5_6_i,temp_b1_5_8_r,temp_b1_5_8_i,temp_b1_7_6_r,temp_b1_7_6_i,temp_b1_7_8_r,temp_b1_7_8_i,temp_m2_5_6_r,temp_m2_5_6_i,temp_m2_5_8_r,temp_m2_5_8_i,temp_m2_7_6_r,temp_m2_7_6_i,temp_m2_7_8_r,temp_m2_7_8_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly86 (clk,temp_m2_5_6_r,temp_m2_5_6_i,temp_m2_5_8_r,temp_m2_5_8_i,temp_m2_7_6_r,temp_m2_7_6_i,temp_m2_7_8_r,temp_m2_7_8_i,temp_b2_5_6_r,temp_b2_5_6_i,temp_b2_5_8_r,temp_b2_5_8_i,temp_b2_7_6_r,temp_b2_7_6_i,temp_b2_7_8_r,temp_b2_7_8_i);
MULT MULT87 (clk,temp_b1_6_5_r,temp_b1_6_5_i,temp_b1_6_7_r,temp_b1_6_7_i,temp_b1_8_5_r,temp_b1_8_5_i,temp_b1_8_7_r,temp_b1_8_7_i,temp_m2_6_5_r,temp_m2_6_5_i,temp_m2_6_7_r,temp_m2_6_7_i,temp_m2_8_5_r,temp_m2_8_5_i,temp_m2_8_7_r,temp_m2_8_7_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly87 (clk,temp_m2_6_5_r,temp_m2_6_5_i,temp_m2_6_7_r,temp_m2_6_7_i,temp_m2_8_5_r,temp_m2_8_5_i,temp_m2_8_7_r,temp_m2_8_7_i,temp_b2_6_5_r,temp_b2_6_5_i,temp_b2_6_7_r,temp_b2_6_7_i,temp_b2_8_5_r,temp_b2_8_5_i,temp_b2_8_7_r,temp_b2_8_7_i);
MULT MULT88 (clk,temp_b1_6_6_r,temp_b1_6_6_i,temp_b1_6_8_r,temp_b1_6_8_i,temp_b1_8_6_r,temp_b1_8_6_i,temp_b1_8_8_r,temp_b1_8_8_i,temp_m2_6_6_r,temp_m2_6_6_i,temp_m2_6_8_r,temp_m2_6_8_i,temp_m2_8_6_r,temp_m2_8_6_i,temp_m2_8_8_r,temp_m2_8_8_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly88 (clk,temp_m2_6_6_r,temp_m2_6_6_i,temp_m2_6_8_r,temp_m2_6_8_i,temp_m2_8_6_r,temp_m2_8_6_i,temp_m2_8_8_r,temp_m2_8_8_i,temp_b2_6_6_r,temp_b2_6_6_i,temp_b2_6_8_r,temp_b2_6_8_i,temp_b2_8_6_r,temp_b2_8_6_i,temp_b2_8_8_r,temp_b2_8_8_i);
MULT MULT89 (clk,temp_b1_5_9_r,temp_b1_5_9_i,temp_b1_5_11_r,temp_b1_5_11_i,temp_b1_7_9_r,temp_b1_7_9_i,temp_b1_7_11_r,temp_b1_7_11_i,temp_m2_5_9_r,temp_m2_5_9_i,temp_m2_5_11_r,temp_m2_5_11_i,temp_m2_7_9_r,temp_m2_7_9_i,temp_m2_7_11_r,temp_m2_7_11_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly89 (clk,temp_m2_5_9_r,temp_m2_5_9_i,temp_m2_5_11_r,temp_m2_5_11_i,temp_m2_7_9_r,temp_m2_7_9_i,temp_m2_7_11_r,temp_m2_7_11_i,temp_b2_5_9_r,temp_b2_5_9_i,temp_b2_5_11_r,temp_b2_5_11_i,temp_b2_7_9_r,temp_b2_7_9_i,temp_b2_7_11_r,temp_b2_7_11_i);
MULT MULT90 (clk,temp_b1_5_10_r,temp_b1_5_10_i,temp_b1_5_12_r,temp_b1_5_12_i,temp_b1_7_10_r,temp_b1_7_10_i,temp_b1_7_12_r,temp_b1_7_12_i,temp_m2_5_10_r,temp_m2_5_10_i,temp_m2_5_12_r,temp_m2_5_12_i,temp_m2_7_10_r,temp_m2_7_10_i,temp_m2_7_12_r,temp_m2_7_12_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly90 (clk,temp_m2_5_10_r,temp_m2_5_10_i,temp_m2_5_12_r,temp_m2_5_12_i,temp_m2_7_10_r,temp_m2_7_10_i,temp_m2_7_12_r,temp_m2_7_12_i,temp_b2_5_10_r,temp_b2_5_10_i,temp_b2_5_12_r,temp_b2_5_12_i,temp_b2_7_10_r,temp_b2_7_10_i,temp_b2_7_12_r,temp_b2_7_12_i);
MULT MULT91 (clk,temp_b1_6_9_r,temp_b1_6_9_i,temp_b1_6_11_r,temp_b1_6_11_i,temp_b1_8_9_r,temp_b1_8_9_i,temp_b1_8_11_r,temp_b1_8_11_i,temp_m2_6_9_r,temp_m2_6_9_i,temp_m2_6_11_r,temp_m2_6_11_i,temp_m2_8_9_r,temp_m2_8_9_i,temp_m2_8_11_r,temp_m2_8_11_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly91 (clk,temp_m2_6_9_r,temp_m2_6_9_i,temp_m2_6_11_r,temp_m2_6_11_i,temp_m2_8_9_r,temp_m2_8_9_i,temp_m2_8_11_r,temp_m2_8_11_i,temp_b2_6_9_r,temp_b2_6_9_i,temp_b2_6_11_r,temp_b2_6_11_i,temp_b2_8_9_r,temp_b2_8_9_i,temp_b2_8_11_r,temp_b2_8_11_i);
MULT MULT92 (clk,temp_b1_6_10_r,temp_b1_6_10_i,temp_b1_6_12_r,temp_b1_6_12_i,temp_b1_8_10_r,temp_b1_8_10_i,temp_b1_8_12_r,temp_b1_8_12_i,temp_m2_6_10_r,temp_m2_6_10_i,temp_m2_6_12_r,temp_m2_6_12_i,temp_m2_8_10_r,temp_m2_8_10_i,temp_m2_8_12_r,temp_m2_8_12_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly92 (clk,temp_m2_6_10_r,temp_m2_6_10_i,temp_m2_6_12_r,temp_m2_6_12_i,temp_m2_8_10_r,temp_m2_8_10_i,temp_m2_8_12_r,temp_m2_8_12_i,temp_b2_6_10_r,temp_b2_6_10_i,temp_b2_6_12_r,temp_b2_6_12_i,temp_b2_8_10_r,temp_b2_8_10_i,temp_b2_8_12_r,temp_b2_8_12_i);
MULT MULT93 (clk,temp_b1_5_13_r,temp_b1_5_13_i,temp_b1_5_15_r,temp_b1_5_15_i,temp_b1_7_13_r,temp_b1_7_13_i,temp_b1_7_15_r,temp_b1_7_15_i,temp_m2_5_13_r,temp_m2_5_13_i,temp_m2_5_15_r,temp_m2_5_15_i,temp_m2_7_13_r,temp_m2_7_13_i,temp_m2_7_15_r,temp_m2_7_15_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly93 (clk,temp_m2_5_13_r,temp_m2_5_13_i,temp_m2_5_15_r,temp_m2_5_15_i,temp_m2_7_13_r,temp_m2_7_13_i,temp_m2_7_15_r,temp_m2_7_15_i,temp_b2_5_13_r,temp_b2_5_13_i,temp_b2_5_15_r,temp_b2_5_15_i,temp_b2_7_13_r,temp_b2_7_13_i,temp_b2_7_15_r,temp_b2_7_15_i);
MULT MULT94 (clk,temp_b1_5_14_r,temp_b1_5_14_i,temp_b1_5_16_r,temp_b1_5_16_i,temp_b1_7_14_r,temp_b1_7_14_i,temp_b1_7_16_r,temp_b1_7_16_i,temp_m2_5_14_r,temp_m2_5_14_i,temp_m2_5_16_r,temp_m2_5_16_i,temp_m2_7_14_r,temp_m2_7_14_i,temp_m2_7_16_r,temp_m2_7_16_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly94 (clk,temp_m2_5_14_r,temp_m2_5_14_i,temp_m2_5_16_r,temp_m2_5_16_i,temp_m2_7_14_r,temp_m2_7_14_i,temp_m2_7_16_r,temp_m2_7_16_i,temp_b2_5_14_r,temp_b2_5_14_i,temp_b2_5_16_r,temp_b2_5_16_i,temp_b2_7_14_r,temp_b2_7_14_i,temp_b2_7_16_r,temp_b2_7_16_i);
MULT MULT95 (clk,temp_b1_6_13_r,temp_b1_6_13_i,temp_b1_6_15_r,temp_b1_6_15_i,temp_b1_8_13_r,temp_b1_8_13_i,temp_b1_8_15_r,temp_b1_8_15_i,temp_m2_6_13_r,temp_m2_6_13_i,temp_m2_6_15_r,temp_m2_6_15_i,temp_m2_8_13_r,temp_m2_8_13_i,temp_m2_8_15_r,temp_m2_8_15_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly95 (clk,temp_m2_6_13_r,temp_m2_6_13_i,temp_m2_6_15_r,temp_m2_6_15_i,temp_m2_8_13_r,temp_m2_8_13_i,temp_m2_8_15_r,temp_m2_8_15_i,temp_b2_6_13_r,temp_b2_6_13_i,temp_b2_6_15_r,temp_b2_6_15_i,temp_b2_8_13_r,temp_b2_8_13_i,temp_b2_8_15_r,temp_b2_8_15_i);
MULT MULT96 (clk,temp_b1_6_14_r,temp_b1_6_14_i,temp_b1_6_16_r,temp_b1_6_16_i,temp_b1_8_14_r,temp_b1_8_14_i,temp_b1_8_16_r,temp_b1_8_16_i,temp_m2_6_14_r,temp_m2_6_14_i,temp_m2_6_16_r,temp_m2_6_16_i,temp_m2_8_14_r,temp_m2_8_14_i,temp_m2_8_16_r,temp_m2_8_16_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly96 (clk,temp_m2_6_14_r,temp_m2_6_14_i,temp_m2_6_16_r,temp_m2_6_16_i,temp_m2_8_14_r,temp_m2_8_14_i,temp_m2_8_16_r,temp_m2_8_16_i,temp_b2_6_14_r,temp_b2_6_14_i,temp_b2_6_16_r,temp_b2_6_16_i,temp_b2_8_14_r,temp_b2_8_14_i,temp_b2_8_16_r,temp_b2_8_16_i);
MULT MULT97 (clk,temp_b1_9_1_r,temp_b1_9_1_i,temp_b1_9_3_r,temp_b1_9_3_i,temp_b1_11_1_r,temp_b1_11_1_i,temp_b1_11_3_r,temp_b1_11_3_i,temp_m2_9_1_r,temp_m2_9_1_i,temp_m2_9_3_r,temp_m2_9_3_i,temp_m2_11_1_r,temp_m2_11_1_i,temp_m2_11_3_r,temp_m2_11_3_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly97 (clk,temp_m2_9_1_r,temp_m2_9_1_i,temp_m2_9_3_r,temp_m2_9_3_i,temp_m2_11_1_r,temp_m2_11_1_i,temp_m2_11_3_r,temp_m2_11_3_i,temp_b2_9_1_r,temp_b2_9_1_i,temp_b2_9_3_r,temp_b2_9_3_i,temp_b2_11_1_r,temp_b2_11_1_i,temp_b2_11_3_r,temp_b2_11_3_i);
MULT MULT98 (clk,temp_b1_9_2_r,temp_b1_9_2_i,temp_b1_9_4_r,temp_b1_9_4_i,temp_b1_11_2_r,temp_b1_11_2_i,temp_b1_11_4_r,temp_b1_11_4_i,temp_m2_9_2_r,temp_m2_9_2_i,temp_m2_9_4_r,temp_m2_9_4_i,temp_m2_11_2_r,temp_m2_11_2_i,temp_m2_11_4_r,temp_m2_11_4_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly98 (clk,temp_m2_9_2_r,temp_m2_9_2_i,temp_m2_9_4_r,temp_m2_9_4_i,temp_m2_11_2_r,temp_m2_11_2_i,temp_m2_11_4_r,temp_m2_11_4_i,temp_b2_9_2_r,temp_b2_9_2_i,temp_b2_9_4_r,temp_b2_9_4_i,temp_b2_11_2_r,temp_b2_11_2_i,temp_b2_11_4_r,temp_b2_11_4_i);
MULT MULT99 (clk,temp_b1_10_1_r,temp_b1_10_1_i,temp_b1_10_3_r,temp_b1_10_3_i,temp_b1_12_1_r,temp_b1_12_1_i,temp_b1_12_3_r,temp_b1_12_3_i,temp_m2_10_1_r,temp_m2_10_1_i,temp_m2_10_3_r,temp_m2_10_3_i,temp_m2_12_1_r,temp_m2_12_1_i,temp_m2_12_3_r,temp_m2_12_3_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly99 (clk,temp_m2_10_1_r,temp_m2_10_1_i,temp_m2_10_3_r,temp_m2_10_3_i,temp_m2_12_1_r,temp_m2_12_1_i,temp_m2_12_3_r,temp_m2_12_3_i,temp_b2_10_1_r,temp_b2_10_1_i,temp_b2_10_3_r,temp_b2_10_3_i,temp_b2_12_1_r,temp_b2_12_1_i,temp_b2_12_3_r,temp_b2_12_3_i);
MULT MULT100 (clk,temp_b1_10_2_r,temp_b1_10_2_i,temp_b1_10_4_r,temp_b1_10_4_i,temp_b1_12_2_r,temp_b1_12_2_i,temp_b1_12_4_r,temp_b1_12_4_i,temp_m2_10_2_r,temp_m2_10_2_i,temp_m2_10_4_r,temp_m2_10_4_i,temp_m2_12_2_r,temp_m2_12_2_i,temp_m2_12_4_r,temp_m2_12_4_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly100 (clk,temp_m2_10_2_r,temp_m2_10_2_i,temp_m2_10_4_r,temp_m2_10_4_i,temp_m2_12_2_r,temp_m2_12_2_i,temp_m2_12_4_r,temp_m2_12_4_i,temp_b2_10_2_r,temp_b2_10_2_i,temp_b2_10_4_r,temp_b2_10_4_i,temp_b2_12_2_r,temp_b2_12_2_i,temp_b2_12_4_r,temp_b2_12_4_i);
MULT MULT101 (clk,temp_b1_9_5_r,temp_b1_9_5_i,temp_b1_9_7_r,temp_b1_9_7_i,temp_b1_11_5_r,temp_b1_11_5_i,temp_b1_11_7_r,temp_b1_11_7_i,temp_m2_9_5_r,temp_m2_9_5_i,temp_m2_9_7_r,temp_m2_9_7_i,temp_m2_11_5_r,temp_m2_11_5_i,temp_m2_11_7_r,temp_m2_11_7_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly101 (clk,temp_m2_9_5_r,temp_m2_9_5_i,temp_m2_9_7_r,temp_m2_9_7_i,temp_m2_11_5_r,temp_m2_11_5_i,temp_m2_11_7_r,temp_m2_11_7_i,temp_b2_9_5_r,temp_b2_9_5_i,temp_b2_9_7_r,temp_b2_9_7_i,temp_b2_11_5_r,temp_b2_11_5_i,temp_b2_11_7_r,temp_b2_11_7_i);
MULT MULT102 (clk,temp_b1_9_6_r,temp_b1_9_6_i,temp_b1_9_8_r,temp_b1_9_8_i,temp_b1_11_6_r,temp_b1_11_6_i,temp_b1_11_8_r,temp_b1_11_8_i,temp_m2_9_6_r,temp_m2_9_6_i,temp_m2_9_8_r,temp_m2_9_8_i,temp_m2_11_6_r,temp_m2_11_6_i,temp_m2_11_8_r,temp_m2_11_8_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly102 (clk,temp_m2_9_6_r,temp_m2_9_6_i,temp_m2_9_8_r,temp_m2_9_8_i,temp_m2_11_6_r,temp_m2_11_6_i,temp_m2_11_8_r,temp_m2_11_8_i,temp_b2_9_6_r,temp_b2_9_6_i,temp_b2_9_8_r,temp_b2_9_8_i,temp_b2_11_6_r,temp_b2_11_6_i,temp_b2_11_8_r,temp_b2_11_8_i);
MULT MULT103 (clk,temp_b1_10_5_r,temp_b1_10_5_i,temp_b1_10_7_r,temp_b1_10_7_i,temp_b1_12_5_r,temp_b1_12_5_i,temp_b1_12_7_r,temp_b1_12_7_i,temp_m2_10_5_r,temp_m2_10_5_i,temp_m2_10_7_r,temp_m2_10_7_i,temp_m2_12_5_r,temp_m2_12_5_i,temp_m2_12_7_r,temp_m2_12_7_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly103 (clk,temp_m2_10_5_r,temp_m2_10_5_i,temp_m2_10_7_r,temp_m2_10_7_i,temp_m2_12_5_r,temp_m2_12_5_i,temp_m2_12_7_r,temp_m2_12_7_i,temp_b2_10_5_r,temp_b2_10_5_i,temp_b2_10_7_r,temp_b2_10_7_i,temp_b2_12_5_r,temp_b2_12_5_i,temp_b2_12_7_r,temp_b2_12_7_i);
MULT MULT104 (clk,temp_b1_10_6_r,temp_b1_10_6_i,temp_b1_10_8_r,temp_b1_10_8_i,temp_b1_12_6_r,temp_b1_12_6_i,temp_b1_12_8_r,temp_b1_12_8_i,temp_m2_10_6_r,temp_m2_10_6_i,temp_m2_10_8_r,temp_m2_10_8_i,temp_m2_12_6_r,temp_m2_12_6_i,temp_m2_12_8_r,temp_m2_12_8_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly104 (clk,temp_m2_10_6_r,temp_m2_10_6_i,temp_m2_10_8_r,temp_m2_10_8_i,temp_m2_12_6_r,temp_m2_12_6_i,temp_m2_12_8_r,temp_m2_12_8_i,temp_b2_10_6_r,temp_b2_10_6_i,temp_b2_10_8_r,temp_b2_10_8_i,temp_b2_12_6_r,temp_b2_12_6_i,temp_b2_12_8_r,temp_b2_12_8_i);
MULT MULT105 (clk,temp_b1_9_9_r,temp_b1_9_9_i,temp_b1_9_11_r,temp_b1_9_11_i,temp_b1_11_9_r,temp_b1_11_9_i,temp_b1_11_11_r,temp_b1_11_11_i,temp_m2_9_9_r,temp_m2_9_9_i,temp_m2_9_11_r,temp_m2_9_11_i,temp_m2_11_9_r,temp_m2_11_9_i,temp_m2_11_11_r,temp_m2_11_11_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly105 (clk,temp_m2_9_9_r,temp_m2_9_9_i,temp_m2_9_11_r,temp_m2_9_11_i,temp_m2_11_9_r,temp_m2_11_9_i,temp_m2_11_11_r,temp_m2_11_11_i,temp_b2_9_9_r,temp_b2_9_9_i,temp_b2_9_11_r,temp_b2_9_11_i,temp_b2_11_9_r,temp_b2_11_9_i,temp_b2_11_11_r,temp_b2_11_11_i);
MULT MULT106 (clk,temp_b1_9_10_r,temp_b1_9_10_i,temp_b1_9_12_r,temp_b1_9_12_i,temp_b1_11_10_r,temp_b1_11_10_i,temp_b1_11_12_r,temp_b1_11_12_i,temp_m2_9_10_r,temp_m2_9_10_i,temp_m2_9_12_r,temp_m2_9_12_i,temp_m2_11_10_r,temp_m2_11_10_i,temp_m2_11_12_r,temp_m2_11_12_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly106 (clk,temp_m2_9_10_r,temp_m2_9_10_i,temp_m2_9_12_r,temp_m2_9_12_i,temp_m2_11_10_r,temp_m2_11_10_i,temp_m2_11_12_r,temp_m2_11_12_i,temp_b2_9_10_r,temp_b2_9_10_i,temp_b2_9_12_r,temp_b2_9_12_i,temp_b2_11_10_r,temp_b2_11_10_i,temp_b2_11_12_r,temp_b2_11_12_i);
MULT MULT107 (clk,temp_b1_10_9_r,temp_b1_10_9_i,temp_b1_10_11_r,temp_b1_10_11_i,temp_b1_12_9_r,temp_b1_12_9_i,temp_b1_12_11_r,temp_b1_12_11_i,temp_m2_10_9_r,temp_m2_10_9_i,temp_m2_10_11_r,temp_m2_10_11_i,temp_m2_12_9_r,temp_m2_12_9_i,temp_m2_12_11_r,temp_m2_12_11_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly107 (clk,temp_m2_10_9_r,temp_m2_10_9_i,temp_m2_10_11_r,temp_m2_10_11_i,temp_m2_12_9_r,temp_m2_12_9_i,temp_m2_12_11_r,temp_m2_12_11_i,temp_b2_10_9_r,temp_b2_10_9_i,temp_b2_10_11_r,temp_b2_10_11_i,temp_b2_12_9_r,temp_b2_12_9_i,temp_b2_12_11_r,temp_b2_12_11_i);
MULT MULT108 (clk,temp_b1_10_10_r,temp_b1_10_10_i,temp_b1_10_12_r,temp_b1_10_12_i,temp_b1_12_10_r,temp_b1_12_10_i,temp_b1_12_12_r,temp_b1_12_12_i,temp_m2_10_10_r,temp_m2_10_10_i,temp_m2_10_12_r,temp_m2_10_12_i,temp_m2_12_10_r,temp_m2_12_10_i,temp_m2_12_12_r,temp_m2_12_12_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly108 (clk,temp_m2_10_10_r,temp_m2_10_10_i,temp_m2_10_12_r,temp_m2_10_12_i,temp_m2_12_10_r,temp_m2_12_10_i,temp_m2_12_12_r,temp_m2_12_12_i,temp_b2_10_10_r,temp_b2_10_10_i,temp_b2_10_12_r,temp_b2_10_12_i,temp_b2_12_10_r,temp_b2_12_10_i,temp_b2_12_12_r,temp_b2_12_12_i);
MULT MULT109 (clk,temp_b1_9_13_r,temp_b1_9_13_i,temp_b1_9_15_r,temp_b1_9_15_i,temp_b1_11_13_r,temp_b1_11_13_i,temp_b1_11_15_r,temp_b1_11_15_i,temp_m2_9_13_r,temp_m2_9_13_i,temp_m2_9_15_r,temp_m2_9_15_i,temp_m2_11_13_r,temp_m2_11_13_i,temp_m2_11_15_r,temp_m2_11_15_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly109 (clk,temp_m2_9_13_r,temp_m2_9_13_i,temp_m2_9_15_r,temp_m2_9_15_i,temp_m2_11_13_r,temp_m2_11_13_i,temp_m2_11_15_r,temp_m2_11_15_i,temp_b2_9_13_r,temp_b2_9_13_i,temp_b2_9_15_r,temp_b2_9_15_i,temp_b2_11_13_r,temp_b2_11_13_i,temp_b2_11_15_r,temp_b2_11_15_i);
MULT MULT110 (clk,temp_b1_9_14_r,temp_b1_9_14_i,temp_b1_9_16_r,temp_b1_9_16_i,temp_b1_11_14_r,temp_b1_11_14_i,temp_b1_11_16_r,temp_b1_11_16_i,temp_m2_9_14_r,temp_m2_9_14_i,temp_m2_9_16_r,temp_m2_9_16_i,temp_m2_11_14_r,temp_m2_11_14_i,temp_m2_11_16_r,temp_m2_11_16_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly110 (clk,temp_m2_9_14_r,temp_m2_9_14_i,temp_m2_9_16_r,temp_m2_9_16_i,temp_m2_11_14_r,temp_m2_11_14_i,temp_m2_11_16_r,temp_m2_11_16_i,temp_b2_9_14_r,temp_b2_9_14_i,temp_b2_9_16_r,temp_b2_9_16_i,temp_b2_11_14_r,temp_b2_11_14_i,temp_b2_11_16_r,temp_b2_11_16_i);
MULT MULT111 (clk,temp_b1_10_13_r,temp_b1_10_13_i,temp_b1_10_15_r,temp_b1_10_15_i,temp_b1_12_13_r,temp_b1_12_13_i,temp_b1_12_15_r,temp_b1_12_15_i,temp_m2_10_13_r,temp_m2_10_13_i,temp_m2_10_15_r,temp_m2_10_15_i,temp_m2_12_13_r,temp_m2_12_13_i,temp_m2_12_15_r,temp_m2_12_15_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly111 (clk,temp_m2_10_13_r,temp_m2_10_13_i,temp_m2_10_15_r,temp_m2_10_15_i,temp_m2_12_13_r,temp_m2_12_13_i,temp_m2_12_15_r,temp_m2_12_15_i,temp_b2_10_13_r,temp_b2_10_13_i,temp_b2_10_15_r,temp_b2_10_15_i,temp_b2_12_13_r,temp_b2_12_13_i,temp_b2_12_15_r,temp_b2_12_15_i);
MULT MULT112 (clk,temp_b1_10_14_r,temp_b1_10_14_i,temp_b1_10_16_r,temp_b1_10_16_i,temp_b1_12_14_r,temp_b1_12_14_i,temp_b1_12_16_r,temp_b1_12_16_i,temp_m2_10_14_r,temp_m2_10_14_i,temp_m2_10_16_r,temp_m2_10_16_i,temp_m2_12_14_r,temp_m2_12_14_i,temp_m2_12_16_r,temp_m2_12_16_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly112 (clk,temp_m2_10_14_r,temp_m2_10_14_i,temp_m2_10_16_r,temp_m2_10_16_i,temp_m2_12_14_r,temp_m2_12_14_i,temp_m2_12_16_r,temp_m2_12_16_i,temp_b2_10_14_r,temp_b2_10_14_i,temp_b2_10_16_r,temp_b2_10_16_i,temp_b2_12_14_r,temp_b2_12_14_i,temp_b2_12_16_r,temp_b2_12_16_i);
MULT MULT113 (clk,temp_b1_13_1_r,temp_b1_13_1_i,temp_b1_13_3_r,temp_b1_13_3_i,temp_b1_15_1_r,temp_b1_15_1_i,temp_b1_15_3_r,temp_b1_15_3_i,temp_m2_13_1_r,temp_m2_13_1_i,temp_m2_13_3_r,temp_m2_13_3_i,temp_m2_15_1_r,temp_m2_15_1_i,temp_m2_15_3_r,temp_m2_15_3_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly113 (clk,temp_m2_13_1_r,temp_m2_13_1_i,temp_m2_13_3_r,temp_m2_13_3_i,temp_m2_15_1_r,temp_m2_15_1_i,temp_m2_15_3_r,temp_m2_15_3_i,temp_b2_13_1_r,temp_b2_13_1_i,temp_b2_13_3_r,temp_b2_13_3_i,temp_b2_15_1_r,temp_b2_15_1_i,temp_b2_15_3_r,temp_b2_15_3_i);
MULT MULT114 (clk,temp_b1_13_2_r,temp_b1_13_2_i,temp_b1_13_4_r,temp_b1_13_4_i,temp_b1_15_2_r,temp_b1_15_2_i,temp_b1_15_4_r,temp_b1_15_4_i,temp_m2_13_2_r,temp_m2_13_2_i,temp_m2_13_4_r,temp_m2_13_4_i,temp_m2_15_2_r,temp_m2_15_2_i,temp_m2_15_4_r,temp_m2_15_4_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly114 (clk,temp_m2_13_2_r,temp_m2_13_2_i,temp_m2_13_4_r,temp_m2_13_4_i,temp_m2_15_2_r,temp_m2_15_2_i,temp_m2_15_4_r,temp_m2_15_4_i,temp_b2_13_2_r,temp_b2_13_2_i,temp_b2_13_4_r,temp_b2_13_4_i,temp_b2_15_2_r,temp_b2_15_2_i,temp_b2_15_4_r,temp_b2_15_4_i);
MULT MULT115 (clk,temp_b1_14_1_r,temp_b1_14_1_i,temp_b1_14_3_r,temp_b1_14_3_i,temp_b1_16_1_r,temp_b1_16_1_i,temp_b1_16_3_r,temp_b1_16_3_i,temp_m2_14_1_r,temp_m2_14_1_i,temp_m2_14_3_r,temp_m2_14_3_i,temp_m2_16_1_r,temp_m2_16_1_i,temp_m2_16_3_r,temp_m2_16_3_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly115 (clk,temp_m2_14_1_r,temp_m2_14_1_i,temp_m2_14_3_r,temp_m2_14_3_i,temp_m2_16_1_r,temp_m2_16_1_i,temp_m2_16_3_r,temp_m2_16_3_i,temp_b2_14_1_r,temp_b2_14_1_i,temp_b2_14_3_r,temp_b2_14_3_i,temp_b2_16_1_r,temp_b2_16_1_i,temp_b2_16_3_r,temp_b2_16_3_i);
MULT MULT116 (clk,temp_b1_14_2_r,temp_b1_14_2_i,temp_b1_14_4_r,temp_b1_14_4_i,temp_b1_16_2_r,temp_b1_16_2_i,temp_b1_16_4_r,temp_b1_16_4_i,temp_m2_14_2_r,temp_m2_14_2_i,temp_m2_14_4_r,temp_m2_14_4_i,temp_m2_16_2_r,temp_m2_16_2_i,temp_m2_16_4_r,temp_m2_16_4_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly116 (clk,temp_m2_14_2_r,temp_m2_14_2_i,temp_m2_14_4_r,temp_m2_14_4_i,temp_m2_16_2_r,temp_m2_16_2_i,temp_m2_16_4_r,temp_m2_16_4_i,temp_b2_14_2_r,temp_b2_14_2_i,temp_b2_14_4_r,temp_b2_14_4_i,temp_b2_16_2_r,temp_b2_16_2_i,temp_b2_16_4_r,temp_b2_16_4_i);
MULT MULT117 (clk,temp_b1_13_5_r,temp_b1_13_5_i,temp_b1_13_7_r,temp_b1_13_7_i,temp_b1_15_5_r,temp_b1_15_5_i,temp_b1_15_7_r,temp_b1_15_7_i,temp_m2_13_5_r,temp_m2_13_5_i,temp_m2_13_7_r,temp_m2_13_7_i,temp_m2_15_5_r,temp_m2_15_5_i,temp_m2_15_7_r,temp_m2_15_7_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly117 (clk,temp_m2_13_5_r,temp_m2_13_5_i,temp_m2_13_7_r,temp_m2_13_7_i,temp_m2_15_5_r,temp_m2_15_5_i,temp_m2_15_7_r,temp_m2_15_7_i,temp_b2_13_5_r,temp_b2_13_5_i,temp_b2_13_7_r,temp_b2_13_7_i,temp_b2_15_5_r,temp_b2_15_5_i,temp_b2_15_7_r,temp_b2_15_7_i);
MULT MULT118 (clk,temp_b1_13_6_r,temp_b1_13_6_i,temp_b1_13_8_r,temp_b1_13_8_i,temp_b1_15_6_r,temp_b1_15_6_i,temp_b1_15_8_r,temp_b1_15_8_i,temp_m2_13_6_r,temp_m2_13_6_i,temp_m2_13_8_r,temp_m2_13_8_i,temp_m2_15_6_r,temp_m2_15_6_i,temp_m2_15_8_r,temp_m2_15_8_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly118 (clk,temp_m2_13_6_r,temp_m2_13_6_i,temp_m2_13_8_r,temp_m2_13_8_i,temp_m2_15_6_r,temp_m2_15_6_i,temp_m2_15_8_r,temp_m2_15_8_i,temp_b2_13_6_r,temp_b2_13_6_i,temp_b2_13_8_r,temp_b2_13_8_i,temp_b2_15_6_r,temp_b2_15_6_i,temp_b2_15_8_r,temp_b2_15_8_i);
MULT MULT119 (clk,temp_b1_14_5_r,temp_b1_14_5_i,temp_b1_14_7_r,temp_b1_14_7_i,temp_b1_16_5_r,temp_b1_16_5_i,temp_b1_16_7_r,temp_b1_16_7_i,temp_m2_14_5_r,temp_m2_14_5_i,temp_m2_14_7_r,temp_m2_14_7_i,temp_m2_16_5_r,temp_m2_16_5_i,temp_m2_16_7_r,temp_m2_16_7_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly119 (clk,temp_m2_14_5_r,temp_m2_14_5_i,temp_m2_14_7_r,temp_m2_14_7_i,temp_m2_16_5_r,temp_m2_16_5_i,temp_m2_16_7_r,temp_m2_16_7_i,temp_b2_14_5_r,temp_b2_14_5_i,temp_b2_14_7_r,temp_b2_14_7_i,temp_b2_16_5_r,temp_b2_16_5_i,temp_b2_16_7_r,temp_b2_16_7_i);
MULT MULT120 (clk,temp_b1_14_6_r,temp_b1_14_6_i,temp_b1_14_8_r,temp_b1_14_8_i,temp_b1_16_6_r,temp_b1_16_6_i,temp_b1_16_8_r,temp_b1_16_8_i,temp_m2_14_6_r,temp_m2_14_6_i,temp_m2_14_8_r,temp_m2_14_8_i,temp_m2_16_6_r,temp_m2_16_6_i,temp_m2_16_8_r,temp_m2_16_8_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly120 (clk,temp_m2_14_6_r,temp_m2_14_6_i,temp_m2_14_8_r,temp_m2_14_8_i,temp_m2_16_6_r,temp_m2_16_6_i,temp_m2_16_8_r,temp_m2_16_8_i,temp_b2_14_6_r,temp_b2_14_6_i,temp_b2_14_8_r,temp_b2_14_8_i,temp_b2_16_6_r,temp_b2_16_6_i,temp_b2_16_8_r,temp_b2_16_8_i);
MULT MULT121 (clk,temp_b1_13_9_r,temp_b1_13_9_i,temp_b1_13_11_r,temp_b1_13_11_i,temp_b1_15_9_r,temp_b1_15_9_i,temp_b1_15_11_r,temp_b1_15_11_i,temp_m2_13_9_r,temp_m2_13_9_i,temp_m2_13_11_r,temp_m2_13_11_i,temp_m2_15_9_r,temp_m2_15_9_i,temp_m2_15_11_r,temp_m2_15_11_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly121 (clk,temp_m2_13_9_r,temp_m2_13_9_i,temp_m2_13_11_r,temp_m2_13_11_i,temp_m2_15_9_r,temp_m2_15_9_i,temp_m2_15_11_r,temp_m2_15_11_i,temp_b2_13_9_r,temp_b2_13_9_i,temp_b2_13_11_r,temp_b2_13_11_i,temp_b2_15_9_r,temp_b2_15_9_i,temp_b2_15_11_r,temp_b2_15_11_i);
MULT MULT122 (clk,temp_b1_13_10_r,temp_b1_13_10_i,temp_b1_13_12_r,temp_b1_13_12_i,temp_b1_15_10_r,temp_b1_15_10_i,temp_b1_15_12_r,temp_b1_15_12_i,temp_m2_13_10_r,temp_m2_13_10_i,temp_m2_13_12_r,temp_m2_13_12_i,temp_m2_15_10_r,temp_m2_15_10_i,temp_m2_15_12_r,temp_m2_15_12_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly122 (clk,temp_m2_13_10_r,temp_m2_13_10_i,temp_m2_13_12_r,temp_m2_13_12_i,temp_m2_15_10_r,temp_m2_15_10_i,temp_m2_15_12_r,temp_m2_15_12_i,temp_b2_13_10_r,temp_b2_13_10_i,temp_b2_13_12_r,temp_b2_13_12_i,temp_b2_15_10_r,temp_b2_15_10_i,temp_b2_15_12_r,temp_b2_15_12_i);
MULT MULT123 (clk,temp_b1_14_9_r,temp_b1_14_9_i,temp_b1_14_11_r,temp_b1_14_11_i,temp_b1_16_9_r,temp_b1_16_9_i,temp_b1_16_11_r,temp_b1_16_11_i,temp_m2_14_9_r,temp_m2_14_9_i,temp_m2_14_11_r,temp_m2_14_11_i,temp_m2_16_9_r,temp_m2_16_9_i,temp_m2_16_11_r,temp_m2_16_11_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly123 (clk,temp_m2_14_9_r,temp_m2_14_9_i,temp_m2_14_11_r,temp_m2_14_11_i,temp_m2_16_9_r,temp_m2_16_9_i,temp_m2_16_11_r,temp_m2_16_11_i,temp_b2_14_9_r,temp_b2_14_9_i,temp_b2_14_11_r,temp_b2_14_11_i,temp_b2_16_9_r,temp_b2_16_9_i,temp_b2_16_11_r,temp_b2_16_11_i);
MULT MULT124 (clk,temp_b1_14_10_r,temp_b1_14_10_i,temp_b1_14_12_r,temp_b1_14_12_i,temp_b1_16_10_r,temp_b1_16_10_i,temp_b1_16_12_r,temp_b1_16_12_i,temp_m2_14_10_r,temp_m2_14_10_i,temp_m2_14_12_r,temp_m2_14_12_i,temp_m2_16_10_r,temp_m2_16_10_i,temp_m2_16_12_r,temp_m2_16_12_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly124 (clk,temp_m2_14_10_r,temp_m2_14_10_i,temp_m2_14_12_r,temp_m2_14_12_i,temp_m2_16_10_r,temp_m2_16_10_i,temp_m2_16_12_r,temp_m2_16_12_i,temp_b2_14_10_r,temp_b2_14_10_i,temp_b2_14_12_r,temp_b2_14_12_i,temp_b2_16_10_r,temp_b2_16_10_i,temp_b2_16_12_r,temp_b2_16_12_i);
MULT MULT125 (clk,temp_b1_13_13_r,temp_b1_13_13_i,temp_b1_13_15_r,temp_b1_13_15_i,temp_b1_15_13_r,temp_b1_15_13_i,temp_b1_15_15_r,temp_b1_15_15_i,temp_m2_13_13_r,temp_m2_13_13_i,temp_m2_13_15_r,temp_m2_13_15_i,temp_m2_15_13_r,temp_m2_15_13_i,temp_m2_15_15_r,temp_m2_15_15_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly125 (clk,temp_m2_13_13_r,temp_m2_13_13_i,temp_m2_13_15_r,temp_m2_13_15_i,temp_m2_15_13_r,temp_m2_15_13_i,temp_m2_15_15_r,temp_m2_15_15_i,temp_b2_13_13_r,temp_b2_13_13_i,temp_b2_13_15_r,temp_b2_13_15_i,temp_b2_15_13_r,temp_b2_15_13_i,temp_b2_15_15_r,temp_b2_15_15_i);
MULT MULT126 (clk,temp_b1_13_14_r,temp_b1_13_14_i,temp_b1_13_16_r,temp_b1_13_16_i,temp_b1_15_14_r,temp_b1_15_14_i,temp_b1_15_16_r,temp_b1_15_16_i,temp_m2_13_14_r,temp_m2_13_14_i,temp_m2_13_16_r,temp_m2_13_16_i,temp_m2_15_14_r,temp_m2_15_14_i,temp_m2_15_16_r,temp_m2_15_16_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly126 (clk,temp_m2_13_14_r,temp_m2_13_14_i,temp_m2_13_16_r,temp_m2_13_16_i,temp_m2_15_14_r,temp_m2_15_14_i,temp_m2_15_16_r,temp_m2_15_16_i,temp_b2_13_14_r,temp_b2_13_14_i,temp_b2_13_16_r,temp_b2_13_16_i,temp_b2_15_14_r,temp_b2_15_14_i,temp_b2_15_16_r,temp_b2_15_16_i);
MULT MULT127 (clk,temp_b1_14_13_r,temp_b1_14_13_i,temp_b1_14_15_r,temp_b1_14_15_i,temp_b1_16_13_r,temp_b1_16_13_i,temp_b1_16_15_r,temp_b1_16_15_i,temp_m2_14_13_r,temp_m2_14_13_i,temp_m2_14_15_r,temp_m2_14_15_i,temp_m2_16_13_r,temp_m2_16_13_i,temp_m2_16_15_r,temp_m2_16_15_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly127 (clk,temp_m2_14_13_r,temp_m2_14_13_i,temp_m2_14_15_r,temp_m2_14_15_i,temp_m2_16_13_r,temp_m2_16_13_i,temp_m2_16_15_r,temp_m2_16_15_i,temp_b2_14_13_r,temp_b2_14_13_i,temp_b2_14_15_r,temp_b2_14_15_i,temp_b2_16_13_r,temp_b2_16_13_i,temp_b2_16_15_r,temp_b2_16_15_i);
MULT MULT128 (clk,temp_b1_14_14_r,temp_b1_14_14_i,temp_b1_14_16_r,temp_b1_14_16_i,temp_b1_16_14_r,temp_b1_16_14_i,temp_b1_16_16_r,temp_b1_16_16_i,temp_m2_14_14_r,temp_m2_14_14_i,temp_m2_14_16_r,temp_m2_14_16_i,temp_m2_16_14_r,temp_m2_16_14_i,temp_m2_16_16_r,temp_m2_16_16_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly128 (clk,temp_m2_14_14_r,temp_m2_14_14_i,temp_m2_14_16_r,temp_m2_14_16_i,temp_m2_16_14_r,temp_m2_16_14_i,temp_m2_16_16_r,temp_m2_16_16_i,temp_b2_14_14_r,temp_b2_14_14_i,temp_b2_14_16_r,temp_b2_14_16_i,temp_b2_16_14_r,temp_b2_16_14_i,temp_b2_16_16_r,temp_b2_16_16_i);
MULT MULT129 (clk,temp_b2_1_1_r,temp_b2_1_1_i,temp_b2_1_5_r,temp_b2_1_5_i,temp_b2_5_1_r,temp_b2_5_1_i,temp_b2_5_5_r,temp_b2_5_5_i,temp_m3_1_1_r,temp_m3_1_1_i,temp_m3_1_5_r,temp_m3_1_5_i,temp_m3_5_1_r,temp_m3_5_1_i,temp_m3_5_5_r,temp_m3_5_5_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly129 (clk,temp_m3_1_1_r,temp_m3_1_1_i,temp_m3_1_5_r,temp_m3_1_5_i,temp_m3_5_1_r,temp_m3_5_1_i,temp_m3_5_5_r,temp_m3_5_5_i,temp_b3_1_1_r,temp_b3_1_1_i,temp_b3_1_5_r,temp_b3_1_5_i,temp_b3_5_1_r,temp_b3_5_1_i,temp_b3_5_5_r,temp_b3_5_5_i);
MULT MULT130 (clk,temp_b2_1_2_r,temp_b2_1_2_i,temp_b2_1_6_r,temp_b2_1_6_i,temp_b2_5_2_r,temp_b2_5_2_i,temp_b2_5_6_r,temp_b2_5_6_i,temp_m3_1_2_r,temp_m3_1_2_i,temp_m3_1_6_r,temp_m3_1_6_i,temp_m3_5_2_r,temp_m3_5_2_i,temp_m3_5_6_r,temp_m3_5_6_i,`W2_real,`W2_imag,`W0_real,`W0_imag,`W2_real,`W2_imag);
butterfly butterfly130 (clk,temp_m3_1_2_r,temp_m3_1_2_i,temp_m3_1_6_r,temp_m3_1_6_i,temp_m3_5_2_r,temp_m3_5_2_i,temp_m3_5_6_r,temp_m3_5_6_i,temp_b3_1_2_r,temp_b3_1_2_i,temp_b3_1_6_r,temp_b3_1_6_i,temp_b3_5_2_r,temp_b3_5_2_i,temp_b3_5_6_r,temp_b3_5_6_i);
MULT MULT131 (clk,temp_b2_1_3_r,temp_b2_1_3_i,temp_b2_1_7_r,temp_b2_1_7_i,temp_b2_5_3_r,temp_b2_5_3_i,temp_b2_5_7_r,temp_b2_5_7_i,temp_m3_1_3_r,temp_m3_1_3_i,temp_m3_1_7_r,temp_m3_1_7_i,temp_m3_5_3_r,temp_m3_5_3_i,temp_m3_5_7_r,temp_m3_5_7_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly131 (clk,temp_m3_1_3_r,temp_m3_1_3_i,temp_m3_1_7_r,temp_m3_1_7_i,temp_m3_5_3_r,temp_m3_5_3_i,temp_m3_5_7_r,temp_m3_5_7_i,temp_b3_1_3_r,temp_b3_1_3_i,temp_b3_1_7_r,temp_b3_1_7_i,temp_b3_5_3_r,temp_b3_5_3_i,temp_b3_5_7_r,temp_b3_5_7_i);
MULT MULT132 (clk,temp_b2_1_4_r,temp_b2_1_4_i,temp_b2_1_8_r,temp_b2_1_8_i,temp_b2_5_4_r,temp_b2_5_4_i,temp_b2_5_8_r,temp_b2_5_8_i,temp_m3_1_4_r,temp_m3_1_4_i,temp_m3_1_8_r,temp_m3_1_8_i,temp_m3_5_4_r,temp_m3_5_4_i,temp_m3_5_8_r,temp_m3_5_8_i,`W6_real,`W6_imag,`W0_real,`W0_imag,`W6_real,`W6_imag);
butterfly butterfly132 (clk,temp_m3_1_4_r,temp_m3_1_4_i,temp_m3_1_8_r,temp_m3_1_8_i,temp_m3_5_4_r,temp_m3_5_4_i,temp_m3_5_8_r,temp_m3_5_8_i,temp_b3_1_4_r,temp_b3_1_4_i,temp_b3_1_8_r,temp_b3_1_8_i,temp_b3_5_4_r,temp_b3_5_4_i,temp_b3_5_8_r,temp_b3_5_8_i);
MULT MULT133 (clk,temp_b2_2_1_r,temp_b2_2_1_i,temp_b2_2_5_r,temp_b2_2_5_i,temp_b2_6_1_r,temp_b2_6_1_i,temp_b2_6_5_r,temp_b2_6_5_i,temp_m3_2_1_r,temp_m3_2_1_i,temp_m3_2_5_r,temp_m3_2_5_i,temp_m3_6_1_r,temp_m3_6_1_i,temp_m3_6_5_r,temp_m3_6_5_i,`W0_real,`W0_imag,`W2_real,`W2_imag,`W2_real,`W2_imag);
butterfly butterfly133 (clk,temp_m3_2_1_r,temp_m3_2_1_i,temp_m3_2_5_r,temp_m3_2_5_i,temp_m3_6_1_r,temp_m3_6_1_i,temp_m3_6_5_r,temp_m3_6_5_i,temp_b3_2_1_r,temp_b3_2_1_i,temp_b3_2_5_r,temp_b3_2_5_i,temp_b3_6_1_r,temp_b3_6_1_i,temp_b3_6_5_r,temp_b3_6_5_i);
MULT MULT134 (clk,temp_b2_2_2_r,temp_b2_2_2_i,temp_b2_2_6_r,temp_b2_2_6_i,temp_b2_6_2_r,temp_b2_6_2_i,temp_b2_6_6_r,temp_b2_6_6_i,temp_m3_2_2_r,temp_m3_2_2_i,temp_m3_2_6_r,temp_m3_2_6_i,temp_m3_6_2_r,temp_m3_6_2_i,temp_m3_6_6_r,temp_m3_6_6_i,`W2_real,`W2_imag,`W2_real,`W2_imag,`W4_real,`W4_imag);
butterfly butterfly134 (clk,temp_m3_2_2_r,temp_m3_2_2_i,temp_m3_2_6_r,temp_m3_2_6_i,temp_m3_6_2_r,temp_m3_6_2_i,temp_m3_6_6_r,temp_m3_6_6_i,temp_b3_2_2_r,temp_b3_2_2_i,temp_b3_2_6_r,temp_b3_2_6_i,temp_b3_6_2_r,temp_b3_6_2_i,temp_b3_6_6_r,temp_b3_6_6_i);
MULT MULT135 (clk,temp_b2_2_3_r,temp_b2_2_3_i,temp_b2_2_7_r,temp_b2_2_7_i,temp_b2_6_3_r,temp_b2_6_3_i,temp_b2_6_7_r,temp_b2_6_7_i,temp_m3_2_3_r,temp_m3_2_3_i,temp_m3_2_7_r,temp_m3_2_7_i,temp_m3_6_3_r,temp_m3_6_3_i,temp_m3_6_7_r,temp_m3_6_7_i,`W4_real,`W4_imag,`W2_real,`W2_imag,`W6_real,`W6_imag);
butterfly butterfly135 (clk,temp_m3_2_3_r,temp_m3_2_3_i,temp_m3_2_7_r,temp_m3_2_7_i,temp_m3_6_3_r,temp_m3_6_3_i,temp_m3_6_7_r,temp_m3_6_7_i,temp_b3_2_3_r,temp_b3_2_3_i,temp_b3_2_7_r,temp_b3_2_7_i,temp_b3_6_3_r,temp_b3_6_3_i,temp_b3_6_7_r,temp_b3_6_7_i);
MULT MULT136 (clk,temp_b2_2_4_r,temp_b2_2_4_i,temp_b2_2_8_r,temp_b2_2_8_i,temp_b2_6_4_r,temp_b2_6_4_i,temp_b2_6_8_r,temp_b2_6_8_i,temp_m3_2_4_r,temp_m3_2_4_i,temp_m3_2_8_r,temp_m3_2_8_i,temp_m3_6_4_r,temp_m3_6_4_i,temp_m3_6_8_r,temp_m3_6_8_i,`W6_real,`W6_imag,`W2_real,`W2_imag,`W8_real,`W8_imag);
butterfly butterfly136 (clk,temp_m3_2_4_r,temp_m3_2_4_i,temp_m3_2_8_r,temp_m3_2_8_i,temp_m3_6_4_r,temp_m3_6_4_i,temp_m3_6_8_r,temp_m3_6_8_i,temp_b3_2_4_r,temp_b3_2_4_i,temp_b3_2_8_r,temp_b3_2_8_i,temp_b3_6_4_r,temp_b3_6_4_i,temp_b3_6_8_r,temp_b3_6_8_i);
MULT MULT137 (clk,temp_b2_3_1_r,temp_b2_3_1_i,temp_b2_3_5_r,temp_b2_3_5_i,temp_b2_7_1_r,temp_b2_7_1_i,temp_b2_7_5_r,temp_b2_7_5_i,temp_m3_3_1_r,temp_m3_3_1_i,temp_m3_3_5_r,temp_m3_3_5_i,temp_m3_7_1_r,temp_m3_7_1_i,temp_m3_7_5_r,temp_m3_7_5_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly137 (clk,temp_m3_3_1_r,temp_m3_3_1_i,temp_m3_3_5_r,temp_m3_3_5_i,temp_m3_7_1_r,temp_m3_7_1_i,temp_m3_7_5_r,temp_m3_7_5_i,temp_b3_3_1_r,temp_b3_3_1_i,temp_b3_3_5_r,temp_b3_3_5_i,temp_b3_7_1_r,temp_b3_7_1_i,temp_b3_7_5_r,temp_b3_7_5_i);
MULT MULT138 (clk,temp_b2_3_2_r,temp_b2_3_2_i,temp_b2_3_6_r,temp_b2_3_6_i,temp_b2_7_2_r,temp_b2_7_2_i,temp_b2_7_6_r,temp_b2_7_6_i,temp_m3_3_2_r,temp_m3_3_2_i,temp_m3_3_6_r,temp_m3_3_6_i,temp_m3_7_2_r,temp_m3_7_2_i,temp_m3_7_6_r,temp_m3_7_6_i,`W2_real,`W2_imag,`W4_real,`W4_imag,`W6_real,`W6_imag);
butterfly butterfly138 (clk,temp_m3_3_2_r,temp_m3_3_2_i,temp_m3_3_6_r,temp_m3_3_6_i,temp_m3_7_2_r,temp_m3_7_2_i,temp_m3_7_6_r,temp_m3_7_6_i,temp_b3_3_2_r,temp_b3_3_2_i,temp_b3_3_6_r,temp_b3_3_6_i,temp_b3_7_2_r,temp_b3_7_2_i,temp_b3_7_6_r,temp_b3_7_6_i);
MULT MULT139 (clk,temp_b2_3_3_r,temp_b2_3_3_i,temp_b2_3_7_r,temp_b2_3_7_i,temp_b2_7_3_r,temp_b2_7_3_i,temp_b2_7_7_r,temp_b2_7_7_i,temp_m3_3_3_r,temp_m3_3_3_i,temp_m3_3_7_r,temp_m3_3_7_i,temp_m3_7_3_r,temp_m3_7_3_i,temp_m3_7_7_r,temp_m3_7_7_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly139 (clk,temp_m3_3_3_r,temp_m3_3_3_i,temp_m3_3_7_r,temp_m3_3_7_i,temp_m3_7_3_r,temp_m3_7_3_i,temp_m3_7_7_r,temp_m3_7_7_i,temp_b3_3_3_r,temp_b3_3_3_i,temp_b3_3_7_r,temp_b3_3_7_i,temp_b3_7_3_r,temp_b3_7_3_i,temp_b3_7_7_r,temp_b3_7_7_i);
MULT MULT140 (clk,temp_b2_3_4_r,temp_b2_3_4_i,temp_b2_3_8_r,temp_b2_3_8_i,temp_b2_7_4_r,temp_b2_7_4_i,temp_b2_7_8_r,temp_b2_7_8_i,temp_m3_3_4_r,temp_m3_3_4_i,temp_m3_3_8_r,temp_m3_3_8_i,temp_m3_7_4_r,temp_m3_7_4_i,temp_m3_7_8_r,temp_m3_7_8_i,`W6_real,`W6_imag,`W4_real,`W4_imag,`W10_real,`W10_imag);
butterfly butterfly140 (clk,temp_m3_3_4_r,temp_m3_3_4_i,temp_m3_3_8_r,temp_m3_3_8_i,temp_m3_7_4_r,temp_m3_7_4_i,temp_m3_7_8_r,temp_m3_7_8_i,temp_b3_3_4_r,temp_b3_3_4_i,temp_b3_3_8_r,temp_b3_3_8_i,temp_b3_7_4_r,temp_b3_7_4_i,temp_b3_7_8_r,temp_b3_7_8_i);
MULT MULT141 (clk,temp_b2_4_1_r,temp_b2_4_1_i,temp_b2_4_5_r,temp_b2_4_5_i,temp_b2_8_1_r,temp_b2_8_1_i,temp_b2_8_5_r,temp_b2_8_5_i,temp_m3_4_1_r,temp_m3_4_1_i,temp_m3_4_5_r,temp_m3_4_5_i,temp_m3_8_1_r,temp_m3_8_1_i,temp_m3_8_5_r,temp_m3_8_5_i,`W0_real,`W0_imag,`W6_real,`W6_imag,`W6_real,`W6_imag);
butterfly butterfly141 (clk,temp_m3_4_1_r,temp_m3_4_1_i,temp_m3_4_5_r,temp_m3_4_5_i,temp_m3_8_1_r,temp_m3_8_1_i,temp_m3_8_5_r,temp_m3_8_5_i,temp_b3_4_1_r,temp_b3_4_1_i,temp_b3_4_5_r,temp_b3_4_5_i,temp_b3_8_1_r,temp_b3_8_1_i,temp_b3_8_5_r,temp_b3_8_5_i);
MULT MULT142 (clk,temp_b2_4_2_r,temp_b2_4_2_i,temp_b2_4_6_r,temp_b2_4_6_i,temp_b2_8_2_r,temp_b2_8_2_i,temp_b2_8_6_r,temp_b2_8_6_i,temp_m3_4_2_r,temp_m3_4_2_i,temp_m3_4_6_r,temp_m3_4_6_i,temp_m3_8_2_r,temp_m3_8_2_i,temp_m3_8_6_r,temp_m3_8_6_i,`W2_real,`W2_imag,`W6_real,`W6_imag,`W8_real,`W8_imag);
butterfly butterfly142 (clk,temp_m3_4_2_r,temp_m3_4_2_i,temp_m3_4_6_r,temp_m3_4_6_i,temp_m3_8_2_r,temp_m3_8_2_i,temp_m3_8_6_r,temp_m3_8_6_i,temp_b3_4_2_r,temp_b3_4_2_i,temp_b3_4_6_r,temp_b3_4_6_i,temp_b3_8_2_r,temp_b3_8_2_i,temp_b3_8_6_r,temp_b3_8_6_i);
MULT MULT143 (clk,temp_b2_4_3_r,temp_b2_4_3_i,temp_b2_4_7_r,temp_b2_4_7_i,temp_b2_8_3_r,temp_b2_8_3_i,temp_b2_8_7_r,temp_b2_8_7_i,temp_m3_4_3_r,temp_m3_4_3_i,temp_m3_4_7_r,temp_m3_4_7_i,temp_m3_8_3_r,temp_m3_8_3_i,temp_m3_8_7_r,temp_m3_8_7_i,`W4_real,`W4_imag,`W6_real,`W6_imag,`W10_real,`W10_imag);
butterfly butterfly143 (clk,temp_m3_4_3_r,temp_m3_4_3_i,temp_m3_4_7_r,temp_m3_4_7_i,temp_m3_8_3_r,temp_m3_8_3_i,temp_m3_8_7_r,temp_m3_8_7_i,temp_b3_4_3_r,temp_b3_4_3_i,temp_b3_4_7_r,temp_b3_4_7_i,temp_b3_8_3_r,temp_b3_8_3_i,temp_b3_8_7_r,temp_b3_8_7_i);
MULT MULT144 (clk,temp_b2_4_4_r,temp_b2_4_4_i,temp_b2_4_8_r,temp_b2_4_8_i,temp_b2_8_4_r,temp_b2_8_4_i,temp_b2_8_8_r,temp_b2_8_8_i,temp_m3_4_4_r,temp_m3_4_4_i,temp_m3_4_8_r,temp_m3_4_8_i,temp_m3_8_4_r,temp_m3_8_4_i,temp_m3_8_8_r,temp_m3_8_8_i,`W6_real,`W6_imag,`W6_real,`W6_imag,`W12_real,`W12_imag);
butterfly butterfly144 (clk,temp_m3_4_4_r,temp_m3_4_4_i,temp_m3_4_8_r,temp_m3_4_8_i,temp_m3_8_4_r,temp_m3_8_4_i,temp_m3_8_8_r,temp_m3_8_8_i,temp_b3_4_4_r,temp_b3_4_4_i,temp_b3_4_8_r,temp_b3_4_8_i,temp_b3_8_4_r,temp_b3_8_4_i,temp_b3_8_8_r,temp_b3_8_8_i);
MULT MULT145 (clk,temp_b2_1_9_r,temp_b2_1_9_i,temp_b2_1_13_r,temp_b2_1_13_i,temp_b2_5_9_r,temp_b2_5_9_i,temp_b2_5_13_r,temp_b2_5_13_i,temp_m3_1_9_r,temp_m3_1_9_i,temp_m3_1_13_r,temp_m3_1_13_i,temp_m3_5_9_r,temp_m3_5_9_i,temp_m3_5_13_r,temp_m3_5_13_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly145 (clk,temp_m3_1_9_r,temp_m3_1_9_i,temp_m3_1_13_r,temp_m3_1_13_i,temp_m3_5_9_r,temp_m3_5_9_i,temp_m3_5_13_r,temp_m3_5_13_i,temp_b3_1_9_r,temp_b3_1_9_i,temp_b3_1_13_r,temp_b3_1_13_i,temp_b3_5_9_r,temp_b3_5_9_i,temp_b3_5_13_r,temp_b3_5_13_i);
MULT MULT146 (clk,temp_b2_1_10_r,temp_b2_1_10_i,temp_b2_1_14_r,temp_b2_1_14_i,temp_b2_5_10_r,temp_b2_5_10_i,temp_b2_5_14_r,temp_b2_5_14_i,temp_m3_1_10_r,temp_m3_1_10_i,temp_m3_1_14_r,temp_m3_1_14_i,temp_m3_5_10_r,temp_m3_5_10_i,temp_m3_5_14_r,temp_m3_5_14_i,`W2_real,`W2_imag,`W0_real,`W0_imag,`W2_real,`W2_imag);
butterfly butterfly146 (clk,temp_m3_1_10_r,temp_m3_1_10_i,temp_m3_1_14_r,temp_m3_1_14_i,temp_m3_5_10_r,temp_m3_5_10_i,temp_m3_5_14_r,temp_m3_5_14_i,temp_b3_1_10_r,temp_b3_1_10_i,temp_b3_1_14_r,temp_b3_1_14_i,temp_b3_5_10_r,temp_b3_5_10_i,temp_b3_5_14_r,temp_b3_5_14_i);
MULT MULT147 (clk,temp_b2_1_11_r,temp_b2_1_11_i,temp_b2_1_15_r,temp_b2_1_15_i,temp_b2_5_11_r,temp_b2_5_11_i,temp_b2_5_15_r,temp_b2_5_15_i,temp_m3_1_11_r,temp_m3_1_11_i,temp_m3_1_15_r,temp_m3_1_15_i,temp_m3_5_11_r,temp_m3_5_11_i,temp_m3_5_15_r,temp_m3_5_15_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly147 (clk,temp_m3_1_11_r,temp_m3_1_11_i,temp_m3_1_15_r,temp_m3_1_15_i,temp_m3_5_11_r,temp_m3_5_11_i,temp_m3_5_15_r,temp_m3_5_15_i,temp_b3_1_11_r,temp_b3_1_11_i,temp_b3_1_15_r,temp_b3_1_15_i,temp_b3_5_11_r,temp_b3_5_11_i,temp_b3_5_15_r,temp_b3_5_15_i);
MULT MULT148 (clk,temp_b2_1_12_r,temp_b2_1_12_i,temp_b2_1_16_r,temp_b2_1_16_i,temp_b2_5_12_r,temp_b2_5_12_i,temp_b2_5_16_r,temp_b2_5_16_i,temp_m3_1_12_r,temp_m3_1_12_i,temp_m3_1_16_r,temp_m3_1_16_i,temp_m3_5_12_r,temp_m3_5_12_i,temp_m3_5_16_r,temp_m3_5_16_i,`W6_real,`W6_imag,`W0_real,`W0_imag,`W6_real,`W6_imag);
butterfly butterfly148 (clk,temp_m3_1_12_r,temp_m3_1_12_i,temp_m3_1_16_r,temp_m3_1_16_i,temp_m3_5_12_r,temp_m3_5_12_i,temp_m3_5_16_r,temp_m3_5_16_i,temp_b3_1_12_r,temp_b3_1_12_i,temp_b3_1_16_r,temp_b3_1_16_i,temp_b3_5_12_r,temp_b3_5_12_i,temp_b3_5_16_r,temp_b3_5_16_i);
MULT MULT149 (clk,temp_b2_2_9_r,temp_b2_2_9_i,temp_b2_2_13_r,temp_b2_2_13_i,temp_b2_6_9_r,temp_b2_6_9_i,temp_b2_6_13_r,temp_b2_6_13_i,temp_m3_2_9_r,temp_m3_2_9_i,temp_m3_2_13_r,temp_m3_2_13_i,temp_m3_6_9_r,temp_m3_6_9_i,temp_m3_6_13_r,temp_m3_6_13_i,`W0_real,`W0_imag,`W2_real,`W2_imag,`W2_real,`W2_imag);
butterfly butterfly149 (clk,temp_m3_2_9_r,temp_m3_2_9_i,temp_m3_2_13_r,temp_m3_2_13_i,temp_m3_6_9_r,temp_m3_6_9_i,temp_m3_6_13_r,temp_m3_6_13_i,temp_b3_2_9_r,temp_b3_2_9_i,temp_b3_2_13_r,temp_b3_2_13_i,temp_b3_6_9_r,temp_b3_6_9_i,temp_b3_6_13_r,temp_b3_6_13_i);
MULT MULT150 (clk,temp_b2_2_10_r,temp_b2_2_10_i,temp_b2_2_14_r,temp_b2_2_14_i,temp_b2_6_10_r,temp_b2_6_10_i,temp_b2_6_14_r,temp_b2_6_14_i,temp_m3_2_10_r,temp_m3_2_10_i,temp_m3_2_14_r,temp_m3_2_14_i,temp_m3_6_10_r,temp_m3_6_10_i,temp_m3_6_14_r,temp_m3_6_14_i,`W2_real,`W2_imag,`W2_real,`W2_imag,`W4_real,`W4_imag);
butterfly butterfly150 (clk,temp_m3_2_10_r,temp_m3_2_10_i,temp_m3_2_14_r,temp_m3_2_14_i,temp_m3_6_10_r,temp_m3_6_10_i,temp_m3_6_14_r,temp_m3_6_14_i,temp_b3_2_10_r,temp_b3_2_10_i,temp_b3_2_14_r,temp_b3_2_14_i,temp_b3_6_10_r,temp_b3_6_10_i,temp_b3_6_14_r,temp_b3_6_14_i);
MULT MULT151 (clk,temp_b2_2_11_r,temp_b2_2_11_i,temp_b2_2_15_r,temp_b2_2_15_i,temp_b2_6_11_r,temp_b2_6_11_i,temp_b2_6_15_r,temp_b2_6_15_i,temp_m3_2_11_r,temp_m3_2_11_i,temp_m3_2_15_r,temp_m3_2_15_i,temp_m3_6_11_r,temp_m3_6_11_i,temp_m3_6_15_r,temp_m3_6_15_i,`W4_real,`W4_imag,`W2_real,`W2_imag,`W6_real,`W6_imag);
butterfly butterfly151 (clk,temp_m3_2_11_r,temp_m3_2_11_i,temp_m3_2_15_r,temp_m3_2_15_i,temp_m3_6_11_r,temp_m3_6_11_i,temp_m3_6_15_r,temp_m3_6_15_i,temp_b3_2_11_r,temp_b3_2_11_i,temp_b3_2_15_r,temp_b3_2_15_i,temp_b3_6_11_r,temp_b3_6_11_i,temp_b3_6_15_r,temp_b3_6_15_i);
MULT MULT152 (clk,temp_b2_2_12_r,temp_b2_2_12_i,temp_b2_2_16_r,temp_b2_2_16_i,temp_b2_6_12_r,temp_b2_6_12_i,temp_b2_6_16_r,temp_b2_6_16_i,temp_m3_2_12_r,temp_m3_2_12_i,temp_m3_2_16_r,temp_m3_2_16_i,temp_m3_6_12_r,temp_m3_6_12_i,temp_m3_6_16_r,temp_m3_6_16_i,`W6_real,`W6_imag,`W2_real,`W2_imag,`W8_real,`W8_imag);
butterfly butterfly152 (clk,temp_m3_2_12_r,temp_m3_2_12_i,temp_m3_2_16_r,temp_m3_2_16_i,temp_m3_6_12_r,temp_m3_6_12_i,temp_m3_6_16_r,temp_m3_6_16_i,temp_b3_2_12_r,temp_b3_2_12_i,temp_b3_2_16_r,temp_b3_2_16_i,temp_b3_6_12_r,temp_b3_6_12_i,temp_b3_6_16_r,temp_b3_6_16_i);
MULT MULT153 (clk,temp_b2_3_9_r,temp_b2_3_9_i,temp_b2_3_13_r,temp_b2_3_13_i,temp_b2_7_9_r,temp_b2_7_9_i,temp_b2_7_13_r,temp_b2_7_13_i,temp_m3_3_9_r,temp_m3_3_9_i,temp_m3_3_13_r,temp_m3_3_13_i,temp_m3_7_9_r,temp_m3_7_9_i,temp_m3_7_13_r,temp_m3_7_13_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly153 (clk,temp_m3_3_9_r,temp_m3_3_9_i,temp_m3_3_13_r,temp_m3_3_13_i,temp_m3_7_9_r,temp_m3_7_9_i,temp_m3_7_13_r,temp_m3_7_13_i,temp_b3_3_9_r,temp_b3_3_9_i,temp_b3_3_13_r,temp_b3_3_13_i,temp_b3_7_9_r,temp_b3_7_9_i,temp_b3_7_13_r,temp_b3_7_13_i);
MULT MULT154 (clk,temp_b2_3_10_r,temp_b2_3_10_i,temp_b2_3_14_r,temp_b2_3_14_i,temp_b2_7_10_r,temp_b2_7_10_i,temp_b2_7_14_r,temp_b2_7_14_i,temp_m3_3_10_r,temp_m3_3_10_i,temp_m3_3_14_r,temp_m3_3_14_i,temp_m3_7_10_r,temp_m3_7_10_i,temp_m3_7_14_r,temp_m3_7_14_i,`W2_real,`W2_imag,`W4_real,`W4_imag,`W6_real,`W6_imag);
butterfly butterfly154 (clk,temp_m3_3_10_r,temp_m3_3_10_i,temp_m3_3_14_r,temp_m3_3_14_i,temp_m3_7_10_r,temp_m3_7_10_i,temp_m3_7_14_r,temp_m3_7_14_i,temp_b3_3_10_r,temp_b3_3_10_i,temp_b3_3_14_r,temp_b3_3_14_i,temp_b3_7_10_r,temp_b3_7_10_i,temp_b3_7_14_r,temp_b3_7_14_i);
MULT MULT155 (clk,temp_b2_3_11_r,temp_b2_3_11_i,temp_b2_3_15_r,temp_b2_3_15_i,temp_b2_7_11_r,temp_b2_7_11_i,temp_b2_7_15_r,temp_b2_7_15_i,temp_m3_3_11_r,temp_m3_3_11_i,temp_m3_3_15_r,temp_m3_3_15_i,temp_m3_7_11_r,temp_m3_7_11_i,temp_m3_7_15_r,temp_m3_7_15_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly155 (clk,temp_m3_3_11_r,temp_m3_3_11_i,temp_m3_3_15_r,temp_m3_3_15_i,temp_m3_7_11_r,temp_m3_7_11_i,temp_m3_7_15_r,temp_m3_7_15_i,temp_b3_3_11_r,temp_b3_3_11_i,temp_b3_3_15_r,temp_b3_3_15_i,temp_b3_7_11_r,temp_b3_7_11_i,temp_b3_7_15_r,temp_b3_7_15_i);
MULT MULT156 (clk,temp_b2_3_12_r,temp_b2_3_12_i,temp_b2_3_16_r,temp_b2_3_16_i,temp_b2_7_12_r,temp_b2_7_12_i,temp_b2_7_16_r,temp_b2_7_16_i,temp_m3_3_12_r,temp_m3_3_12_i,temp_m3_3_16_r,temp_m3_3_16_i,temp_m3_7_12_r,temp_m3_7_12_i,temp_m3_7_16_r,temp_m3_7_16_i,`W6_real,`W6_imag,`W4_real,`W4_imag,`W10_real,`W10_imag);
butterfly butterfly156 (clk,temp_m3_3_12_r,temp_m3_3_12_i,temp_m3_3_16_r,temp_m3_3_16_i,temp_m3_7_12_r,temp_m3_7_12_i,temp_m3_7_16_r,temp_m3_7_16_i,temp_b3_3_12_r,temp_b3_3_12_i,temp_b3_3_16_r,temp_b3_3_16_i,temp_b3_7_12_r,temp_b3_7_12_i,temp_b3_7_16_r,temp_b3_7_16_i);
MULT MULT157 (clk,temp_b2_4_9_r,temp_b2_4_9_i,temp_b2_4_13_r,temp_b2_4_13_i,temp_b2_8_9_r,temp_b2_8_9_i,temp_b2_8_13_r,temp_b2_8_13_i,temp_m3_4_9_r,temp_m3_4_9_i,temp_m3_4_13_r,temp_m3_4_13_i,temp_m3_8_9_r,temp_m3_8_9_i,temp_m3_8_13_r,temp_m3_8_13_i,`W0_real,`W0_imag,`W6_real,`W6_imag,`W6_real,`W6_imag);
butterfly butterfly157 (clk,temp_m3_4_9_r,temp_m3_4_9_i,temp_m3_4_13_r,temp_m3_4_13_i,temp_m3_8_9_r,temp_m3_8_9_i,temp_m3_8_13_r,temp_m3_8_13_i,temp_b3_4_9_r,temp_b3_4_9_i,temp_b3_4_13_r,temp_b3_4_13_i,temp_b3_8_9_r,temp_b3_8_9_i,temp_b3_8_13_r,temp_b3_8_13_i);
MULT MULT158 (clk,temp_b2_4_10_r,temp_b2_4_10_i,temp_b2_4_14_r,temp_b2_4_14_i,temp_b2_8_10_r,temp_b2_8_10_i,temp_b2_8_14_r,temp_b2_8_14_i,temp_m3_4_10_r,temp_m3_4_10_i,temp_m3_4_14_r,temp_m3_4_14_i,temp_m3_8_10_r,temp_m3_8_10_i,temp_m3_8_14_r,temp_m3_8_14_i,`W2_real,`W2_imag,`W6_real,`W6_imag,`W8_real,`W8_imag);
butterfly butterfly158 (clk,temp_m3_4_10_r,temp_m3_4_10_i,temp_m3_4_14_r,temp_m3_4_14_i,temp_m3_8_10_r,temp_m3_8_10_i,temp_m3_8_14_r,temp_m3_8_14_i,temp_b3_4_10_r,temp_b3_4_10_i,temp_b3_4_14_r,temp_b3_4_14_i,temp_b3_8_10_r,temp_b3_8_10_i,temp_b3_8_14_r,temp_b3_8_14_i);
MULT MULT159 (clk,temp_b2_4_11_r,temp_b2_4_11_i,temp_b2_4_15_r,temp_b2_4_15_i,temp_b2_8_11_r,temp_b2_8_11_i,temp_b2_8_15_r,temp_b2_8_15_i,temp_m3_4_11_r,temp_m3_4_11_i,temp_m3_4_15_r,temp_m3_4_15_i,temp_m3_8_11_r,temp_m3_8_11_i,temp_m3_8_15_r,temp_m3_8_15_i,`W4_real,`W4_imag,`W6_real,`W6_imag,`W10_real,`W10_imag);
butterfly butterfly159 (clk,temp_m3_4_11_r,temp_m3_4_11_i,temp_m3_4_15_r,temp_m3_4_15_i,temp_m3_8_11_r,temp_m3_8_11_i,temp_m3_8_15_r,temp_m3_8_15_i,temp_b3_4_11_r,temp_b3_4_11_i,temp_b3_4_15_r,temp_b3_4_15_i,temp_b3_8_11_r,temp_b3_8_11_i,temp_b3_8_15_r,temp_b3_8_15_i);
MULT MULT160 (clk,temp_b2_4_12_r,temp_b2_4_12_i,temp_b2_4_16_r,temp_b2_4_16_i,temp_b2_8_12_r,temp_b2_8_12_i,temp_b2_8_16_r,temp_b2_8_16_i,temp_m3_4_12_r,temp_m3_4_12_i,temp_m3_4_16_r,temp_m3_4_16_i,temp_m3_8_12_r,temp_m3_8_12_i,temp_m3_8_16_r,temp_m3_8_16_i,`W6_real,`W6_imag,`W6_real,`W6_imag,`W12_real,`W12_imag);
butterfly butterfly160 (clk,temp_m3_4_12_r,temp_m3_4_12_i,temp_m3_4_16_r,temp_m3_4_16_i,temp_m3_8_12_r,temp_m3_8_12_i,temp_m3_8_16_r,temp_m3_8_16_i,temp_b3_4_12_r,temp_b3_4_12_i,temp_b3_4_16_r,temp_b3_4_16_i,temp_b3_8_12_r,temp_b3_8_12_i,temp_b3_8_16_r,temp_b3_8_16_i);
MULT MULT161 (clk,temp_b2_9_1_r,temp_b2_9_1_i,temp_b2_9_5_r,temp_b2_9_5_i,temp_b2_13_1_r,temp_b2_13_1_i,temp_b2_13_5_r,temp_b2_13_5_i,temp_m3_9_1_r,temp_m3_9_1_i,temp_m3_9_5_r,temp_m3_9_5_i,temp_m3_13_1_r,temp_m3_13_1_i,temp_m3_13_5_r,temp_m3_13_5_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly161 (clk,temp_m3_9_1_r,temp_m3_9_1_i,temp_m3_9_5_r,temp_m3_9_5_i,temp_m3_13_1_r,temp_m3_13_1_i,temp_m3_13_5_r,temp_m3_13_5_i,temp_b3_9_1_r,temp_b3_9_1_i,temp_b3_9_5_r,temp_b3_9_5_i,temp_b3_13_1_r,temp_b3_13_1_i,temp_b3_13_5_r,temp_b3_13_5_i);
MULT MULT162 (clk,temp_b2_9_2_r,temp_b2_9_2_i,temp_b2_9_6_r,temp_b2_9_6_i,temp_b2_13_2_r,temp_b2_13_2_i,temp_b2_13_6_r,temp_b2_13_6_i,temp_m3_9_2_r,temp_m3_9_2_i,temp_m3_9_6_r,temp_m3_9_6_i,temp_m3_13_2_r,temp_m3_13_2_i,temp_m3_13_6_r,temp_m3_13_6_i,`W2_real,`W2_imag,`W0_real,`W0_imag,`W2_real,`W2_imag);
butterfly butterfly162 (clk,temp_m3_9_2_r,temp_m3_9_2_i,temp_m3_9_6_r,temp_m3_9_6_i,temp_m3_13_2_r,temp_m3_13_2_i,temp_m3_13_6_r,temp_m3_13_6_i,temp_b3_9_2_r,temp_b3_9_2_i,temp_b3_9_6_r,temp_b3_9_6_i,temp_b3_13_2_r,temp_b3_13_2_i,temp_b3_13_6_r,temp_b3_13_6_i);
MULT MULT163 (clk,temp_b2_9_3_r,temp_b2_9_3_i,temp_b2_9_7_r,temp_b2_9_7_i,temp_b2_13_3_r,temp_b2_13_3_i,temp_b2_13_7_r,temp_b2_13_7_i,temp_m3_9_3_r,temp_m3_9_3_i,temp_m3_9_7_r,temp_m3_9_7_i,temp_m3_13_3_r,temp_m3_13_3_i,temp_m3_13_7_r,temp_m3_13_7_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly163 (clk,temp_m3_9_3_r,temp_m3_9_3_i,temp_m3_9_7_r,temp_m3_9_7_i,temp_m3_13_3_r,temp_m3_13_3_i,temp_m3_13_7_r,temp_m3_13_7_i,temp_b3_9_3_r,temp_b3_9_3_i,temp_b3_9_7_r,temp_b3_9_7_i,temp_b3_13_3_r,temp_b3_13_3_i,temp_b3_13_7_r,temp_b3_13_7_i);
MULT MULT164 (clk,temp_b2_9_4_r,temp_b2_9_4_i,temp_b2_9_8_r,temp_b2_9_8_i,temp_b2_13_4_r,temp_b2_13_4_i,temp_b2_13_8_r,temp_b2_13_8_i,temp_m3_9_4_r,temp_m3_9_4_i,temp_m3_9_8_r,temp_m3_9_8_i,temp_m3_13_4_r,temp_m3_13_4_i,temp_m3_13_8_r,temp_m3_13_8_i,`W6_real,`W6_imag,`W0_real,`W0_imag,`W6_real,`W6_imag);
butterfly butterfly164 (clk,temp_m3_9_4_r,temp_m3_9_4_i,temp_m3_9_8_r,temp_m3_9_8_i,temp_m3_13_4_r,temp_m3_13_4_i,temp_m3_13_8_r,temp_m3_13_8_i,temp_b3_9_4_r,temp_b3_9_4_i,temp_b3_9_8_r,temp_b3_9_8_i,temp_b3_13_4_r,temp_b3_13_4_i,temp_b3_13_8_r,temp_b3_13_8_i);
MULT MULT165 (clk,temp_b2_10_1_r,temp_b2_10_1_i,temp_b2_10_5_r,temp_b2_10_5_i,temp_b2_14_1_r,temp_b2_14_1_i,temp_b2_14_5_r,temp_b2_14_5_i,temp_m3_10_1_r,temp_m3_10_1_i,temp_m3_10_5_r,temp_m3_10_5_i,temp_m3_14_1_r,temp_m3_14_1_i,temp_m3_14_5_r,temp_m3_14_5_i,`W0_real,`W0_imag,`W2_real,`W2_imag,`W2_real,`W2_imag);
butterfly butterfly165 (clk,temp_m3_10_1_r,temp_m3_10_1_i,temp_m3_10_5_r,temp_m3_10_5_i,temp_m3_14_1_r,temp_m3_14_1_i,temp_m3_14_5_r,temp_m3_14_5_i,temp_b3_10_1_r,temp_b3_10_1_i,temp_b3_10_5_r,temp_b3_10_5_i,temp_b3_14_1_r,temp_b3_14_1_i,temp_b3_14_5_r,temp_b3_14_5_i);
MULT MULT166 (clk,temp_b2_10_2_r,temp_b2_10_2_i,temp_b2_10_6_r,temp_b2_10_6_i,temp_b2_14_2_r,temp_b2_14_2_i,temp_b2_14_6_r,temp_b2_14_6_i,temp_m3_10_2_r,temp_m3_10_2_i,temp_m3_10_6_r,temp_m3_10_6_i,temp_m3_14_2_r,temp_m3_14_2_i,temp_m3_14_6_r,temp_m3_14_6_i,`W2_real,`W2_imag,`W2_real,`W2_imag,`W4_real,`W4_imag);
butterfly butterfly166 (clk,temp_m3_10_2_r,temp_m3_10_2_i,temp_m3_10_6_r,temp_m3_10_6_i,temp_m3_14_2_r,temp_m3_14_2_i,temp_m3_14_6_r,temp_m3_14_6_i,temp_b3_10_2_r,temp_b3_10_2_i,temp_b3_10_6_r,temp_b3_10_6_i,temp_b3_14_2_r,temp_b3_14_2_i,temp_b3_14_6_r,temp_b3_14_6_i);
MULT MULT167 (clk,temp_b2_10_3_r,temp_b2_10_3_i,temp_b2_10_7_r,temp_b2_10_7_i,temp_b2_14_3_r,temp_b2_14_3_i,temp_b2_14_7_r,temp_b2_14_7_i,temp_m3_10_3_r,temp_m3_10_3_i,temp_m3_10_7_r,temp_m3_10_7_i,temp_m3_14_3_r,temp_m3_14_3_i,temp_m3_14_7_r,temp_m3_14_7_i,`W4_real,`W4_imag,`W2_real,`W2_imag,`W6_real,`W6_imag);
butterfly butterfly167 (clk,temp_m3_10_3_r,temp_m3_10_3_i,temp_m3_10_7_r,temp_m3_10_7_i,temp_m3_14_3_r,temp_m3_14_3_i,temp_m3_14_7_r,temp_m3_14_7_i,temp_b3_10_3_r,temp_b3_10_3_i,temp_b3_10_7_r,temp_b3_10_7_i,temp_b3_14_3_r,temp_b3_14_3_i,temp_b3_14_7_r,temp_b3_14_7_i);
MULT MULT168 (clk,temp_b2_10_4_r,temp_b2_10_4_i,temp_b2_10_8_r,temp_b2_10_8_i,temp_b2_14_4_r,temp_b2_14_4_i,temp_b2_14_8_r,temp_b2_14_8_i,temp_m3_10_4_r,temp_m3_10_4_i,temp_m3_10_8_r,temp_m3_10_8_i,temp_m3_14_4_r,temp_m3_14_4_i,temp_m3_14_8_r,temp_m3_14_8_i,`W6_real,`W6_imag,`W2_real,`W2_imag,`W8_real,`W8_imag);
butterfly butterfly168 (clk,temp_m3_10_4_r,temp_m3_10_4_i,temp_m3_10_8_r,temp_m3_10_8_i,temp_m3_14_4_r,temp_m3_14_4_i,temp_m3_14_8_r,temp_m3_14_8_i,temp_b3_10_4_r,temp_b3_10_4_i,temp_b3_10_8_r,temp_b3_10_8_i,temp_b3_14_4_r,temp_b3_14_4_i,temp_b3_14_8_r,temp_b3_14_8_i);
MULT MULT169 (clk,temp_b2_11_1_r,temp_b2_11_1_i,temp_b2_11_5_r,temp_b2_11_5_i,temp_b2_15_1_r,temp_b2_15_1_i,temp_b2_15_5_r,temp_b2_15_5_i,temp_m3_11_1_r,temp_m3_11_1_i,temp_m3_11_5_r,temp_m3_11_5_i,temp_m3_15_1_r,temp_m3_15_1_i,temp_m3_15_5_r,temp_m3_15_5_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly169 (clk,temp_m3_11_1_r,temp_m3_11_1_i,temp_m3_11_5_r,temp_m3_11_5_i,temp_m3_15_1_r,temp_m3_15_1_i,temp_m3_15_5_r,temp_m3_15_5_i,temp_b3_11_1_r,temp_b3_11_1_i,temp_b3_11_5_r,temp_b3_11_5_i,temp_b3_15_1_r,temp_b3_15_1_i,temp_b3_15_5_r,temp_b3_15_5_i);
MULT MULT170 (clk,temp_b2_11_2_r,temp_b2_11_2_i,temp_b2_11_6_r,temp_b2_11_6_i,temp_b2_15_2_r,temp_b2_15_2_i,temp_b2_15_6_r,temp_b2_15_6_i,temp_m3_11_2_r,temp_m3_11_2_i,temp_m3_11_6_r,temp_m3_11_6_i,temp_m3_15_2_r,temp_m3_15_2_i,temp_m3_15_6_r,temp_m3_15_6_i,`W2_real,`W2_imag,`W4_real,`W4_imag,`W6_real,`W6_imag);
butterfly butterfly170 (clk,temp_m3_11_2_r,temp_m3_11_2_i,temp_m3_11_6_r,temp_m3_11_6_i,temp_m3_15_2_r,temp_m3_15_2_i,temp_m3_15_6_r,temp_m3_15_6_i,temp_b3_11_2_r,temp_b3_11_2_i,temp_b3_11_6_r,temp_b3_11_6_i,temp_b3_15_2_r,temp_b3_15_2_i,temp_b3_15_6_r,temp_b3_15_6_i);
MULT MULT171 (clk,temp_b2_11_3_r,temp_b2_11_3_i,temp_b2_11_7_r,temp_b2_11_7_i,temp_b2_15_3_r,temp_b2_15_3_i,temp_b2_15_7_r,temp_b2_15_7_i,temp_m3_11_3_r,temp_m3_11_3_i,temp_m3_11_7_r,temp_m3_11_7_i,temp_m3_15_3_r,temp_m3_15_3_i,temp_m3_15_7_r,temp_m3_15_7_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly171 (clk,temp_m3_11_3_r,temp_m3_11_3_i,temp_m3_11_7_r,temp_m3_11_7_i,temp_m3_15_3_r,temp_m3_15_3_i,temp_m3_15_7_r,temp_m3_15_7_i,temp_b3_11_3_r,temp_b3_11_3_i,temp_b3_11_7_r,temp_b3_11_7_i,temp_b3_15_3_r,temp_b3_15_3_i,temp_b3_15_7_r,temp_b3_15_7_i);
MULT MULT172 (clk,temp_b2_11_4_r,temp_b2_11_4_i,temp_b2_11_8_r,temp_b2_11_8_i,temp_b2_15_4_r,temp_b2_15_4_i,temp_b2_15_8_r,temp_b2_15_8_i,temp_m3_11_4_r,temp_m3_11_4_i,temp_m3_11_8_r,temp_m3_11_8_i,temp_m3_15_4_r,temp_m3_15_4_i,temp_m3_15_8_r,temp_m3_15_8_i,`W6_real,`W6_imag,`W4_real,`W4_imag,`W10_real,`W10_imag);
butterfly butterfly172 (clk,temp_m3_11_4_r,temp_m3_11_4_i,temp_m3_11_8_r,temp_m3_11_8_i,temp_m3_15_4_r,temp_m3_15_4_i,temp_m3_15_8_r,temp_m3_15_8_i,temp_b3_11_4_r,temp_b3_11_4_i,temp_b3_11_8_r,temp_b3_11_8_i,temp_b3_15_4_r,temp_b3_15_4_i,temp_b3_15_8_r,temp_b3_15_8_i);
MULT MULT173 (clk,temp_b2_12_1_r,temp_b2_12_1_i,temp_b2_12_5_r,temp_b2_12_5_i,temp_b2_16_1_r,temp_b2_16_1_i,temp_b2_16_5_r,temp_b2_16_5_i,temp_m3_12_1_r,temp_m3_12_1_i,temp_m3_12_5_r,temp_m3_12_5_i,temp_m3_16_1_r,temp_m3_16_1_i,temp_m3_16_5_r,temp_m3_16_5_i,`W0_real,`W0_imag,`W6_real,`W6_imag,`W6_real,`W6_imag);
butterfly butterfly173 (clk,temp_m3_12_1_r,temp_m3_12_1_i,temp_m3_12_5_r,temp_m3_12_5_i,temp_m3_16_1_r,temp_m3_16_1_i,temp_m3_16_5_r,temp_m3_16_5_i,temp_b3_12_1_r,temp_b3_12_1_i,temp_b3_12_5_r,temp_b3_12_5_i,temp_b3_16_1_r,temp_b3_16_1_i,temp_b3_16_5_r,temp_b3_16_5_i);
MULT MULT174 (clk,temp_b2_12_2_r,temp_b2_12_2_i,temp_b2_12_6_r,temp_b2_12_6_i,temp_b2_16_2_r,temp_b2_16_2_i,temp_b2_16_6_r,temp_b2_16_6_i,temp_m3_12_2_r,temp_m3_12_2_i,temp_m3_12_6_r,temp_m3_12_6_i,temp_m3_16_2_r,temp_m3_16_2_i,temp_m3_16_6_r,temp_m3_16_6_i,`W2_real,`W2_imag,`W6_real,`W6_imag,`W8_real,`W8_imag);
butterfly butterfly174 (clk,temp_m3_12_2_r,temp_m3_12_2_i,temp_m3_12_6_r,temp_m3_12_6_i,temp_m3_16_2_r,temp_m3_16_2_i,temp_m3_16_6_r,temp_m3_16_6_i,temp_b3_12_2_r,temp_b3_12_2_i,temp_b3_12_6_r,temp_b3_12_6_i,temp_b3_16_2_r,temp_b3_16_2_i,temp_b3_16_6_r,temp_b3_16_6_i);
MULT MULT175 (clk,temp_b2_12_3_r,temp_b2_12_3_i,temp_b2_12_7_r,temp_b2_12_7_i,temp_b2_16_3_r,temp_b2_16_3_i,temp_b2_16_7_r,temp_b2_16_7_i,temp_m3_12_3_r,temp_m3_12_3_i,temp_m3_12_7_r,temp_m3_12_7_i,temp_m3_16_3_r,temp_m3_16_3_i,temp_m3_16_7_r,temp_m3_16_7_i,`W4_real,`W4_imag,`W6_real,`W6_imag,`W10_real,`W10_imag);
butterfly butterfly175 (clk,temp_m3_12_3_r,temp_m3_12_3_i,temp_m3_12_7_r,temp_m3_12_7_i,temp_m3_16_3_r,temp_m3_16_3_i,temp_m3_16_7_r,temp_m3_16_7_i,temp_b3_12_3_r,temp_b3_12_3_i,temp_b3_12_7_r,temp_b3_12_7_i,temp_b3_16_3_r,temp_b3_16_3_i,temp_b3_16_7_r,temp_b3_16_7_i);
MULT MULT176 (clk,temp_b2_12_4_r,temp_b2_12_4_i,temp_b2_12_8_r,temp_b2_12_8_i,temp_b2_16_4_r,temp_b2_16_4_i,temp_b2_16_8_r,temp_b2_16_8_i,temp_m3_12_4_r,temp_m3_12_4_i,temp_m3_12_8_r,temp_m3_12_8_i,temp_m3_16_4_r,temp_m3_16_4_i,temp_m3_16_8_r,temp_m3_16_8_i,`W6_real,`W6_imag,`W6_real,`W6_imag,`W12_real,`W12_imag);
butterfly butterfly176 (clk,temp_m3_12_4_r,temp_m3_12_4_i,temp_m3_12_8_r,temp_m3_12_8_i,temp_m3_16_4_r,temp_m3_16_4_i,temp_m3_16_8_r,temp_m3_16_8_i,temp_b3_12_4_r,temp_b3_12_4_i,temp_b3_12_8_r,temp_b3_12_8_i,temp_b3_16_4_r,temp_b3_16_4_i,temp_b3_16_8_r,temp_b3_16_8_i);
MULT MULT177 (clk,temp_b2_9_9_r,temp_b2_9_9_i,temp_b2_9_13_r,temp_b2_9_13_i,temp_b2_13_9_r,temp_b2_13_9_i,temp_b2_13_13_r,temp_b2_13_13_i,temp_m3_9_9_r,temp_m3_9_9_i,temp_m3_9_13_r,temp_m3_9_13_i,temp_m3_13_9_r,temp_m3_13_9_i,temp_m3_13_13_r,temp_m3_13_13_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly177 (clk,temp_m3_9_9_r,temp_m3_9_9_i,temp_m3_9_13_r,temp_m3_9_13_i,temp_m3_13_9_r,temp_m3_13_9_i,temp_m3_13_13_r,temp_m3_13_13_i,temp_b3_9_9_r,temp_b3_9_9_i,temp_b3_9_13_r,temp_b3_9_13_i,temp_b3_13_9_r,temp_b3_13_9_i,temp_b3_13_13_r,temp_b3_13_13_i);
MULT MULT178 (clk,temp_b2_9_10_r,temp_b2_9_10_i,temp_b2_9_14_r,temp_b2_9_14_i,temp_b2_13_10_r,temp_b2_13_10_i,temp_b2_13_14_r,temp_b2_13_14_i,temp_m3_9_10_r,temp_m3_9_10_i,temp_m3_9_14_r,temp_m3_9_14_i,temp_m3_13_10_r,temp_m3_13_10_i,temp_m3_13_14_r,temp_m3_13_14_i,`W2_real,`W2_imag,`W0_real,`W0_imag,`W2_real,`W2_imag);
butterfly butterfly178 (clk,temp_m3_9_10_r,temp_m3_9_10_i,temp_m3_9_14_r,temp_m3_9_14_i,temp_m3_13_10_r,temp_m3_13_10_i,temp_m3_13_14_r,temp_m3_13_14_i,temp_b3_9_10_r,temp_b3_9_10_i,temp_b3_9_14_r,temp_b3_9_14_i,temp_b3_13_10_r,temp_b3_13_10_i,temp_b3_13_14_r,temp_b3_13_14_i);
MULT MULT179 (clk,temp_b2_9_11_r,temp_b2_9_11_i,temp_b2_9_15_r,temp_b2_9_15_i,temp_b2_13_11_r,temp_b2_13_11_i,temp_b2_13_15_r,temp_b2_13_15_i,temp_m3_9_11_r,temp_m3_9_11_i,temp_m3_9_15_r,temp_m3_9_15_i,temp_m3_13_11_r,temp_m3_13_11_i,temp_m3_13_15_r,temp_m3_13_15_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly179 (clk,temp_m3_9_11_r,temp_m3_9_11_i,temp_m3_9_15_r,temp_m3_9_15_i,temp_m3_13_11_r,temp_m3_13_11_i,temp_m3_13_15_r,temp_m3_13_15_i,temp_b3_9_11_r,temp_b3_9_11_i,temp_b3_9_15_r,temp_b3_9_15_i,temp_b3_13_11_r,temp_b3_13_11_i,temp_b3_13_15_r,temp_b3_13_15_i);
MULT MULT180 (clk,temp_b2_9_12_r,temp_b2_9_12_i,temp_b2_9_16_r,temp_b2_9_16_i,temp_b2_13_12_r,temp_b2_13_12_i,temp_b2_13_16_r,temp_b2_13_16_i,temp_m3_9_12_r,temp_m3_9_12_i,temp_m3_9_16_r,temp_m3_9_16_i,temp_m3_13_12_r,temp_m3_13_12_i,temp_m3_13_16_r,temp_m3_13_16_i,`W6_real,`W6_imag,`W0_real,`W0_imag,`W6_real,`W6_imag);
butterfly butterfly180 (clk,temp_m3_9_12_r,temp_m3_9_12_i,temp_m3_9_16_r,temp_m3_9_16_i,temp_m3_13_12_r,temp_m3_13_12_i,temp_m3_13_16_r,temp_m3_13_16_i,temp_b3_9_12_r,temp_b3_9_12_i,temp_b3_9_16_r,temp_b3_9_16_i,temp_b3_13_12_r,temp_b3_13_12_i,temp_b3_13_16_r,temp_b3_13_16_i);
MULT MULT181 (clk,temp_b2_10_9_r,temp_b2_10_9_i,temp_b2_10_13_r,temp_b2_10_13_i,temp_b2_14_9_r,temp_b2_14_9_i,temp_b2_14_13_r,temp_b2_14_13_i,temp_m3_10_9_r,temp_m3_10_9_i,temp_m3_10_13_r,temp_m3_10_13_i,temp_m3_14_9_r,temp_m3_14_9_i,temp_m3_14_13_r,temp_m3_14_13_i,`W0_real,`W0_imag,`W2_real,`W2_imag,`W2_real,`W2_imag);
butterfly butterfly181 (clk,temp_m3_10_9_r,temp_m3_10_9_i,temp_m3_10_13_r,temp_m3_10_13_i,temp_m3_14_9_r,temp_m3_14_9_i,temp_m3_14_13_r,temp_m3_14_13_i,temp_b3_10_9_r,temp_b3_10_9_i,temp_b3_10_13_r,temp_b3_10_13_i,temp_b3_14_9_r,temp_b3_14_9_i,temp_b3_14_13_r,temp_b3_14_13_i);
MULT MULT182 (clk,temp_b2_10_10_r,temp_b2_10_10_i,temp_b2_10_14_r,temp_b2_10_14_i,temp_b2_14_10_r,temp_b2_14_10_i,temp_b2_14_14_r,temp_b2_14_14_i,temp_m3_10_10_r,temp_m3_10_10_i,temp_m3_10_14_r,temp_m3_10_14_i,temp_m3_14_10_r,temp_m3_14_10_i,temp_m3_14_14_r,temp_m3_14_14_i,`W2_real,`W2_imag,`W2_real,`W2_imag,`W4_real,`W4_imag);
butterfly butterfly182 (clk,temp_m3_10_10_r,temp_m3_10_10_i,temp_m3_10_14_r,temp_m3_10_14_i,temp_m3_14_10_r,temp_m3_14_10_i,temp_m3_14_14_r,temp_m3_14_14_i,temp_b3_10_10_r,temp_b3_10_10_i,temp_b3_10_14_r,temp_b3_10_14_i,temp_b3_14_10_r,temp_b3_14_10_i,temp_b3_14_14_r,temp_b3_14_14_i);
MULT MULT183 (clk,temp_b2_10_11_r,temp_b2_10_11_i,temp_b2_10_15_r,temp_b2_10_15_i,temp_b2_14_11_r,temp_b2_14_11_i,temp_b2_14_15_r,temp_b2_14_15_i,temp_m3_10_11_r,temp_m3_10_11_i,temp_m3_10_15_r,temp_m3_10_15_i,temp_m3_14_11_r,temp_m3_14_11_i,temp_m3_14_15_r,temp_m3_14_15_i,`W4_real,`W4_imag,`W2_real,`W2_imag,`W6_real,`W6_imag);
butterfly butterfly183 (clk,temp_m3_10_11_r,temp_m3_10_11_i,temp_m3_10_15_r,temp_m3_10_15_i,temp_m3_14_11_r,temp_m3_14_11_i,temp_m3_14_15_r,temp_m3_14_15_i,temp_b3_10_11_r,temp_b3_10_11_i,temp_b3_10_15_r,temp_b3_10_15_i,temp_b3_14_11_r,temp_b3_14_11_i,temp_b3_14_15_r,temp_b3_14_15_i);
MULT MULT184 (clk,temp_b2_10_12_r,temp_b2_10_12_i,temp_b2_10_16_r,temp_b2_10_16_i,temp_b2_14_12_r,temp_b2_14_12_i,temp_b2_14_16_r,temp_b2_14_16_i,temp_m3_10_12_r,temp_m3_10_12_i,temp_m3_10_16_r,temp_m3_10_16_i,temp_m3_14_12_r,temp_m3_14_12_i,temp_m3_14_16_r,temp_m3_14_16_i,`W6_real,`W6_imag,`W2_real,`W2_imag,`W8_real,`W8_imag);
butterfly butterfly184 (clk,temp_m3_10_12_r,temp_m3_10_12_i,temp_m3_10_16_r,temp_m3_10_16_i,temp_m3_14_12_r,temp_m3_14_12_i,temp_m3_14_16_r,temp_m3_14_16_i,temp_b3_10_12_r,temp_b3_10_12_i,temp_b3_10_16_r,temp_b3_10_16_i,temp_b3_14_12_r,temp_b3_14_12_i,temp_b3_14_16_r,temp_b3_14_16_i);
MULT MULT185 (clk,temp_b2_11_9_r,temp_b2_11_9_i,temp_b2_11_13_r,temp_b2_11_13_i,temp_b2_15_9_r,temp_b2_15_9_i,temp_b2_15_13_r,temp_b2_15_13_i,temp_m3_11_9_r,temp_m3_11_9_i,temp_m3_11_13_r,temp_m3_11_13_i,temp_m3_15_9_r,temp_m3_15_9_i,temp_m3_15_13_r,temp_m3_15_13_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly185 (clk,temp_m3_11_9_r,temp_m3_11_9_i,temp_m3_11_13_r,temp_m3_11_13_i,temp_m3_15_9_r,temp_m3_15_9_i,temp_m3_15_13_r,temp_m3_15_13_i,temp_b3_11_9_r,temp_b3_11_9_i,temp_b3_11_13_r,temp_b3_11_13_i,temp_b3_15_9_r,temp_b3_15_9_i,temp_b3_15_13_r,temp_b3_15_13_i);
MULT MULT186 (clk,temp_b2_11_10_r,temp_b2_11_10_i,temp_b2_11_14_r,temp_b2_11_14_i,temp_b2_15_10_r,temp_b2_15_10_i,temp_b2_15_14_r,temp_b2_15_14_i,temp_m3_11_10_r,temp_m3_11_10_i,temp_m3_11_14_r,temp_m3_11_14_i,temp_m3_15_10_r,temp_m3_15_10_i,temp_m3_15_14_r,temp_m3_15_14_i,`W2_real,`W2_imag,`W4_real,`W4_imag,`W6_real,`W6_imag);
butterfly butterfly186 (clk,temp_m3_11_10_r,temp_m3_11_10_i,temp_m3_11_14_r,temp_m3_11_14_i,temp_m3_15_10_r,temp_m3_15_10_i,temp_m3_15_14_r,temp_m3_15_14_i,temp_b3_11_10_r,temp_b3_11_10_i,temp_b3_11_14_r,temp_b3_11_14_i,temp_b3_15_10_r,temp_b3_15_10_i,temp_b3_15_14_r,temp_b3_15_14_i);
MULT MULT187 (clk,temp_b2_11_11_r,temp_b2_11_11_i,temp_b2_11_15_r,temp_b2_11_15_i,temp_b2_15_11_r,temp_b2_15_11_i,temp_b2_15_15_r,temp_b2_15_15_i,temp_m3_11_11_r,temp_m3_11_11_i,temp_m3_11_15_r,temp_m3_11_15_i,temp_m3_15_11_r,temp_m3_15_11_i,temp_m3_15_15_r,temp_m3_15_15_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly187 (clk,temp_m3_11_11_r,temp_m3_11_11_i,temp_m3_11_15_r,temp_m3_11_15_i,temp_m3_15_11_r,temp_m3_15_11_i,temp_m3_15_15_r,temp_m3_15_15_i,temp_b3_11_11_r,temp_b3_11_11_i,temp_b3_11_15_r,temp_b3_11_15_i,temp_b3_15_11_r,temp_b3_15_11_i,temp_b3_15_15_r,temp_b3_15_15_i);
MULT MULT188 (clk,temp_b2_11_12_r,temp_b2_11_12_i,temp_b2_11_16_r,temp_b2_11_16_i,temp_b2_15_12_r,temp_b2_15_12_i,temp_b2_15_16_r,temp_b2_15_16_i,temp_m3_11_12_r,temp_m3_11_12_i,temp_m3_11_16_r,temp_m3_11_16_i,temp_m3_15_12_r,temp_m3_15_12_i,temp_m3_15_16_r,temp_m3_15_16_i,`W6_real,`W6_imag,`W4_real,`W4_imag,`W10_real,`W10_imag);
butterfly butterfly188 (clk,temp_m3_11_12_r,temp_m3_11_12_i,temp_m3_11_16_r,temp_m3_11_16_i,temp_m3_15_12_r,temp_m3_15_12_i,temp_m3_15_16_r,temp_m3_15_16_i,temp_b3_11_12_r,temp_b3_11_12_i,temp_b3_11_16_r,temp_b3_11_16_i,temp_b3_15_12_r,temp_b3_15_12_i,temp_b3_15_16_r,temp_b3_15_16_i);
MULT MULT189 (clk,temp_b2_12_9_r,temp_b2_12_9_i,temp_b2_12_13_r,temp_b2_12_13_i,temp_b2_16_9_r,temp_b2_16_9_i,temp_b2_16_13_r,temp_b2_16_13_i,temp_m3_12_9_r,temp_m3_12_9_i,temp_m3_12_13_r,temp_m3_12_13_i,temp_m3_16_9_r,temp_m3_16_9_i,temp_m3_16_13_r,temp_m3_16_13_i,`W0_real,`W0_imag,`W6_real,`W6_imag,`W6_real,`W6_imag);
butterfly butterfly189 (clk,temp_m3_12_9_r,temp_m3_12_9_i,temp_m3_12_13_r,temp_m3_12_13_i,temp_m3_16_9_r,temp_m3_16_9_i,temp_m3_16_13_r,temp_m3_16_13_i,temp_b3_12_9_r,temp_b3_12_9_i,temp_b3_12_13_r,temp_b3_12_13_i,temp_b3_16_9_r,temp_b3_16_9_i,temp_b3_16_13_r,temp_b3_16_13_i);
MULT MULT190 (clk,temp_b2_12_10_r,temp_b2_12_10_i,temp_b2_12_14_r,temp_b2_12_14_i,temp_b2_16_10_r,temp_b2_16_10_i,temp_b2_16_14_r,temp_b2_16_14_i,temp_m3_12_10_r,temp_m3_12_10_i,temp_m3_12_14_r,temp_m3_12_14_i,temp_m3_16_10_r,temp_m3_16_10_i,temp_m3_16_14_r,temp_m3_16_14_i,`W2_real,`W2_imag,`W6_real,`W6_imag,`W8_real,`W8_imag);
butterfly butterfly190 (clk,temp_m3_12_10_r,temp_m3_12_10_i,temp_m3_12_14_r,temp_m3_12_14_i,temp_m3_16_10_r,temp_m3_16_10_i,temp_m3_16_14_r,temp_m3_16_14_i,temp_b3_12_10_r,temp_b3_12_10_i,temp_b3_12_14_r,temp_b3_12_14_i,temp_b3_16_10_r,temp_b3_16_10_i,temp_b3_16_14_r,temp_b3_16_14_i);
MULT MULT191 (clk,temp_b2_12_11_r,temp_b2_12_11_i,temp_b2_12_15_r,temp_b2_12_15_i,temp_b2_16_11_r,temp_b2_16_11_i,temp_b2_16_15_r,temp_b2_16_15_i,temp_m3_12_11_r,temp_m3_12_11_i,temp_m3_12_15_r,temp_m3_12_15_i,temp_m3_16_11_r,temp_m3_16_11_i,temp_m3_16_15_r,temp_m3_16_15_i,`W4_real,`W4_imag,`W6_real,`W6_imag,`W10_real,`W10_imag);
butterfly butterfly191 (clk,temp_m3_12_11_r,temp_m3_12_11_i,temp_m3_12_15_r,temp_m3_12_15_i,temp_m3_16_11_r,temp_m3_16_11_i,temp_m3_16_15_r,temp_m3_16_15_i,temp_b3_12_11_r,temp_b3_12_11_i,temp_b3_12_15_r,temp_b3_12_15_i,temp_b3_16_11_r,temp_b3_16_11_i,temp_b3_16_15_r,temp_b3_16_15_i);
MULT MULT192 (clk,temp_b2_12_12_r,temp_b2_12_12_i,temp_b2_12_16_r,temp_b2_12_16_i,temp_b2_16_12_r,temp_b2_16_12_i,temp_b2_16_16_r,temp_b2_16_16_i,temp_m3_12_12_r,temp_m3_12_12_i,temp_m3_12_16_r,temp_m3_12_16_i,temp_m3_16_12_r,temp_m3_16_12_i,temp_m3_16_16_r,temp_m3_16_16_i,`W6_real,`W6_imag,`W6_real,`W6_imag,`W12_real,`W12_imag);
butterfly butterfly192 (clk,temp_m3_12_12_r,temp_m3_12_12_i,temp_m3_12_16_r,temp_m3_12_16_i,temp_m3_16_12_r,temp_m3_16_12_i,temp_m3_16_16_r,temp_m3_16_16_i,temp_b3_12_12_r,temp_b3_12_12_i,temp_b3_12_16_r,temp_b3_12_16_i,temp_b3_16_12_r,temp_b3_16_12_i,temp_b3_16_16_r,temp_b3_16_16_i);
MULT MULT193 (clk,temp_b3_1_1_r,temp_b3_1_1_i,temp_b3_1_9_r,temp_b3_1_9_i,temp_b3_9_1_r,temp_b3_9_1_i,temp_b3_9_9_r,temp_b3_9_9_i,temp_m4_1_1_r,temp_m4_1_1_i,temp_m4_1_9_r,temp_m4_1_9_i,temp_m4_9_1_r,temp_m4_9_1_i,temp_m4_9_9_r,temp_m4_9_9_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly193 (clk,temp_m4_1_1_r,temp_m4_1_1_i,temp_m4_1_9_r,temp_m4_1_9_i,temp_m4_9_1_r,temp_m4_9_1_i,temp_m4_9_9_r,temp_m4_9_9_i,temp_b4_1_1_r,temp_b4_1_1_i,temp_b4_1_9_r,temp_b4_1_9_i,temp_b4_9_1_r,temp_b4_9_1_i,temp_b4_9_9_r,temp_b4_9_9_i);
MULT MULT194 (clk,temp_b3_1_2_r,temp_b3_1_2_i,temp_b3_1_10_r,temp_b3_1_10_i,temp_b3_9_2_r,temp_b3_9_2_i,temp_b3_9_10_r,temp_b3_9_10_i,temp_m4_1_2_r,temp_m4_1_2_i,temp_m4_1_10_r,temp_m4_1_10_i,temp_m4_9_2_r,temp_m4_9_2_i,temp_m4_9_10_r,temp_m4_9_10_i,`W1_real,`W1_imag,`W0_real,`W0_imag,`W1_real,`W1_imag);
butterfly butterfly194 (clk,temp_m4_1_2_r,temp_m4_1_2_i,temp_m4_1_10_r,temp_m4_1_10_i,temp_m4_9_2_r,temp_m4_9_2_i,temp_m4_9_10_r,temp_m4_9_10_i,temp_b4_1_2_r,temp_b4_1_2_i,temp_b4_1_10_r,temp_b4_1_10_i,temp_b4_9_2_r,temp_b4_9_2_i,temp_b4_9_10_r,temp_b4_9_10_i);
MULT MULT195 (clk,temp_b3_1_3_r,temp_b3_1_3_i,temp_b3_1_11_r,temp_b3_1_11_i,temp_b3_9_3_r,temp_b3_9_3_i,temp_b3_9_11_r,temp_b3_9_11_i,temp_m4_1_3_r,temp_m4_1_3_i,temp_m4_1_11_r,temp_m4_1_11_i,temp_m4_9_3_r,temp_m4_9_3_i,temp_m4_9_11_r,temp_m4_9_11_i,`W2_real,`W2_imag,`W0_real,`W0_imag,`W2_real,`W2_imag);
butterfly butterfly195 (clk,temp_m4_1_3_r,temp_m4_1_3_i,temp_m4_1_11_r,temp_m4_1_11_i,temp_m4_9_3_r,temp_m4_9_3_i,temp_m4_9_11_r,temp_m4_9_11_i,temp_b4_1_3_r,temp_b4_1_3_i,temp_b4_1_11_r,temp_b4_1_11_i,temp_b4_9_3_r,temp_b4_9_3_i,temp_b4_9_11_r,temp_b4_9_11_i);
MULT MULT196 (clk,temp_b3_1_4_r,temp_b3_1_4_i,temp_b3_1_12_r,temp_b3_1_12_i,temp_b3_9_4_r,temp_b3_9_4_i,temp_b3_9_12_r,temp_b3_9_12_i,temp_m4_1_4_r,temp_m4_1_4_i,temp_m4_1_12_r,temp_m4_1_12_i,temp_m4_9_4_r,temp_m4_9_4_i,temp_m4_9_12_r,temp_m4_9_12_i,`W3_real,`W3_imag,`W0_real,`W0_imag,`W3_real,`W3_imag);
butterfly butterfly196 (clk,temp_m4_1_4_r,temp_m4_1_4_i,temp_m4_1_12_r,temp_m4_1_12_i,temp_m4_9_4_r,temp_m4_9_4_i,temp_m4_9_12_r,temp_m4_9_12_i,temp_b4_1_4_r,temp_b4_1_4_i,temp_b4_1_12_r,temp_b4_1_12_i,temp_b4_9_4_r,temp_b4_9_4_i,temp_b4_9_12_r,temp_b4_9_12_i);
MULT MULT197 (clk,temp_b3_1_5_r,temp_b3_1_5_i,temp_b3_1_13_r,temp_b3_1_13_i,temp_b3_9_5_r,temp_b3_9_5_i,temp_b3_9_13_r,temp_b3_9_13_i,temp_m4_1_5_r,temp_m4_1_5_i,temp_m4_1_13_r,temp_m4_1_13_i,temp_m4_9_5_r,temp_m4_9_5_i,temp_m4_9_13_r,temp_m4_9_13_i,`W4_real,`W4_imag,`W0_real,`W0_imag,`W4_real,`W4_imag);
butterfly butterfly197 (clk,temp_m4_1_5_r,temp_m4_1_5_i,temp_m4_1_13_r,temp_m4_1_13_i,temp_m4_9_5_r,temp_m4_9_5_i,temp_m4_9_13_r,temp_m4_9_13_i,temp_b4_1_5_r,temp_b4_1_5_i,temp_b4_1_13_r,temp_b4_1_13_i,temp_b4_9_5_r,temp_b4_9_5_i,temp_b4_9_13_r,temp_b4_9_13_i);
MULT MULT198 (clk,temp_b3_1_6_r,temp_b3_1_6_i,temp_b3_1_14_r,temp_b3_1_14_i,temp_b3_9_6_r,temp_b3_9_6_i,temp_b3_9_14_r,temp_b3_9_14_i,temp_m4_1_6_r,temp_m4_1_6_i,temp_m4_1_14_r,temp_m4_1_14_i,temp_m4_9_6_r,temp_m4_9_6_i,temp_m4_9_14_r,temp_m4_9_14_i,`W5_real,`W5_imag,`W0_real,`W0_imag,`W5_real,`W5_imag);
butterfly butterfly198 (clk,temp_m4_1_6_r,temp_m4_1_6_i,temp_m4_1_14_r,temp_m4_1_14_i,temp_m4_9_6_r,temp_m4_9_6_i,temp_m4_9_14_r,temp_m4_9_14_i,temp_b4_1_6_r,temp_b4_1_6_i,temp_b4_1_14_r,temp_b4_1_14_i,temp_b4_9_6_r,temp_b4_9_6_i,temp_b4_9_14_r,temp_b4_9_14_i);
MULT MULT199 (clk,temp_b3_1_7_r,temp_b3_1_7_i,temp_b3_1_15_r,temp_b3_1_15_i,temp_b3_9_7_r,temp_b3_9_7_i,temp_b3_9_15_r,temp_b3_9_15_i,temp_m4_1_7_r,temp_m4_1_7_i,temp_m4_1_15_r,temp_m4_1_15_i,temp_m4_9_7_r,temp_m4_9_7_i,temp_m4_9_15_r,temp_m4_9_15_i,`W6_real,`W6_imag,`W0_real,`W0_imag,`W6_real,`W6_imag);
butterfly butterfly199 (clk,temp_m4_1_7_r,temp_m4_1_7_i,temp_m4_1_15_r,temp_m4_1_15_i,temp_m4_9_7_r,temp_m4_9_7_i,temp_m4_9_15_r,temp_m4_9_15_i,temp_b4_1_7_r,temp_b4_1_7_i,temp_b4_1_15_r,temp_b4_1_15_i,temp_b4_9_7_r,temp_b4_9_7_i,temp_b4_9_15_r,temp_b4_9_15_i);
MULT MULT200 (clk,temp_b3_1_8_r,temp_b3_1_8_i,temp_b3_1_16_r,temp_b3_1_16_i,temp_b3_9_8_r,temp_b3_9_8_i,temp_b3_9_16_r,temp_b3_9_16_i,temp_m4_1_8_r,temp_m4_1_8_i,temp_m4_1_16_r,temp_m4_1_16_i,temp_m4_9_8_r,temp_m4_9_8_i,temp_m4_9_16_r,temp_m4_9_16_i,`W7_real,`W7_imag,`W0_real,`W0_imag,`W7_real,`W7_imag);
butterfly butterfly200 (clk,temp_m4_1_8_r,temp_m4_1_8_i,temp_m4_1_16_r,temp_m4_1_16_i,temp_m4_9_8_r,temp_m4_9_8_i,temp_m4_9_16_r,temp_m4_9_16_i,temp_b4_1_8_r,temp_b4_1_8_i,temp_b4_1_16_r,temp_b4_1_16_i,temp_b4_9_8_r,temp_b4_9_8_i,temp_b4_9_16_r,temp_b4_9_16_i);
MULT MULT201 (clk,temp_b3_2_1_r,temp_b3_2_1_i,temp_b3_2_9_r,temp_b3_2_9_i,temp_b3_10_1_r,temp_b3_10_1_i,temp_b3_10_9_r,temp_b3_10_9_i,temp_m4_2_1_r,temp_m4_2_1_i,temp_m4_2_9_r,temp_m4_2_9_i,temp_m4_10_1_r,temp_m4_10_1_i,temp_m4_10_9_r,temp_m4_10_9_i,`W0_real,`W0_imag,`W1_real,`W1_imag,`W1_real,`W1_imag);
butterfly butterfly201 (clk,temp_m4_2_1_r,temp_m4_2_1_i,temp_m4_2_9_r,temp_m4_2_9_i,temp_m4_10_1_r,temp_m4_10_1_i,temp_m4_10_9_r,temp_m4_10_9_i,temp_b4_2_1_r,temp_b4_2_1_i,temp_b4_2_9_r,temp_b4_2_9_i,temp_b4_10_1_r,temp_b4_10_1_i,temp_b4_10_9_r,temp_b4_10_9_i);
MULT MULT202 (clk,temp_b3_2_2_r,temp_b3_2_2_i,temp_b3_2_10_r,temp_b3_2_10_i,temp_b3_10_2_r,temp_b3_10_2_i,temp_b3_10_10_r,temp_b3_10_10_i,temp_m4_2_2_r,temp_m4_2_2_i,temp_m4_2_10_r,temp_m4_2_10_i,temp_m4_10_2_r,temp_m4_10_2_i,temp_m4_10_10_r,temp_m4_10_10_i,`W1_real,`W1_imag,`W1_real,`W1_imag,`W2_real,`W2_imag);
butterfly butterfly202 (clk,temp_m4_2_2_r,temp_m4_2_2_i,temp_m4_2_10_r,temp_m4_2_10_i,temp_m4_10_2_r,temp_m4_10_2_i,temp_m4_10_10_r,temp_m4_10_10_i,temp_b4_2_2_r,temp_b4_2_2_i,temp_b4_2_10_r,temp_b4_2_10_i,temp_b4_10_2_r,temp_b4_10_2_i,temp_b4_10_10_r,temp_b4_10_10_i);
MULT MULT203 (clk,temp_b3_2_3_r,temp_b3_2_3_i,temp_b3_2_11_r,temp_b3_2_11_i,temp_b3_10_3_r,temp_b3_10_3_i,temp_b3_10_11_r,temp_b3_10_11_i,temp_m4_2_3_r,temp_m4_2_3_i,temp_m4_2_11_r,temp_m4_2_11_i,temp_m4_10_3_r,temp_m4_10_3_i,temp_m4_10_11_r,temp_m4_10_11_i,`W2_real,`W2_imag,`W1_real,`W1_imag,`W3_real,`W3_imag);
butterfly butterfly203 (clk,temp_m4_2_3_r,temp_m4_2_3_i,temp_m4_2_11_r,temp_m4_2_11_i,temp_m4_10_3_r,temp_m4_10_3_i,temp_m4_10_11_r,temp_m4_10_11_i,temp_b4_2_3_r,temp_b4_2_3_i,temp_b4_2_11_r,temp_b4_2_11_i,temp_b4_10_3_r,temp_b4_10_3_i,temp_b4_10_11_r,temp_b4_10_11_i);
MULT MULT204 (clk,temp_b3_2_4_r,temp_b3_2_4_i,temp_b3_2_12_r,temp_b3_2_12_i,temp_b3_10_4_r,temp_b3_10_4_i,temp_b3_10_12_r,temp_b3_10_12_i,temp_m4_2_4_r,temp_m4_2_4_i,temp_m4_2_12_r,temp_m4_2_12_i,temp_m4_10_4_r,temp_m4_10_4_i,temp_m4_10_12_r,temp_m4_10_12_i,`W3_real,`W3_imag,`W1_real,`W1_imag,`W4_real,`W4_imag);
butterfly butterfly204 (clk,temp_m4_2_4_r,temp_m4_2_4_i,temp_m4_2_12_r,temp_m4_2_12_i,temp_m4_10_4_r,temp_m4_10_4_i,temp_m4_10_12_r,temp_m4_10_12_i,temp_b4_2_4_r,temp_b4_2_4_i,temp_b4_2_12_r,temp_b4_2_12_i,temp_b4_10_4_r,temp_b4_10_4_i,temp_b4_10_12_r,temp_b4_10_12_i);
MULT MULT205 (clk,temp_b3_2_5_r,temp_b3_2_5_i,temp_b3_2_13_r,temp_b3_2_13_i,temp_b3_10_5_r,temp_b3_10_5_i,temp_b3_10_13_r,temp_b3_10_13_i,temp_m4_2_5_r,temp_m4_2_5_i,temp_m4_2_13_r,temp_m4_2_13_i,temp_m4_10_5_r,temp_m4_10_5_i,temp_m4_10_13_r,temp_m4_10_13_i,`W4_real,`W4_imag,`W1_real,`W1_imag,`W5_real,`W5_imag);
butterfly butterfly205 (clk,temp_m4_2_5_r,temp_m4_2_5_i,temp_m4_2_13_r,temp_m4_2_13_i,temp_m4_10_5_r,temp_m4_10_5_i,temp_m4_10_13_r,temp_m4_10_13_i,temp_b4_2_5_r,temp_b4_2_5_i,temp_b4_2_13_r,temp_b4_2_13_i,temp_b4_10_5_r,temp_b4_10_5_i,temp_b4_10_13_r,temp_b4_10_13_i);
MULT MULT206 (clk,temp_b3_2_6_r,temp_b3_2_6_i,temp_b3_2_14_r,temp_b3_2_14_i,temp_b3_10_6_r,temp_b3_10_6_i,temp_b3_10_14_r,temp_b3_10_14_i,temp_m4_2_6_r,temp_m4_2_6_i,temp_m4_2_14_r,temp_m4_2_14_i,temp_m4_10_6_r,temp_m4_10_6_i,temp_m4_10_14_r,temp_m4_10_14_i,`W5_real,`W5_imag,`W1_real,`W1_imag,`W6_real,`W6_imag);
butterfly butterfly206 (clk,temp_m4_2_6_r,temp_m4_2_6_i,temp_m4_2_14_r,temp_m4_2_14_i,temp_m4_10_6_r,temp_m4_10_6_i,temp_m4_10_14_r,temp_m4_10_14_i,temp_b4_2_6_r,temp_b4_2_6_i,temp_b4_2_14_r,temp_b4_2_14_i,temp_b4_10_6_r,temp_b4_10_6_i,temp_b4_10_14_r,temp_b4_10_14_i);
MULT MULT207 (clk,temp_b3_2_7_r,temp_b3_2_7_i,temp_b3_2_15_r,temp_b3_2_15_i,temp_b3_10_7_r,temp_b3_10_7_i,temp_b3_10_15_r,temp_b3_10_15_i,temp_m4_2_7_r,temp_m4_2_7_i,temp_m4_2_15_r,temp_m4_2_15_i,temp_m4_10_7_r,temp_m4_10_7_i,temp_m4_10_15_r,temp_m4_10_15_i,`W6_real,`W6_imag,`W1_real,`W1_imag,`W7_real,`W7_imag);
butterfly butterfly207 (clk,temp_m4_2_7_r,temp_m4_2_7_i,temp_m4_2_15_r,temp_m4_2_15_i,temp_m4_10_7_r,temp_m4_10_7_i,temp_m4_10_15_r,temp_m4_10_15_i,temp_b4_2_7_r,temp_b4_2_7_i,temp_b4_2_15_r,temp_b4_2_15_i,temp_b4_10_7_r,temp_b4_10_7_i,temp_b4_10_15_r,temp_b4_10_15_i);
MULT MULT208 (clk,temp_b3_2_8_r,temp_b3_2_8_i,temp_b3_2_16_r,temp_b3_2_16_i,temp_b3_10_8_r,temp_b3_10_8_i,temp_b3_10_16_r,temp_b3_10_16_i,temp_m4_2_8_r,temp_m4_2_8_i,temp_m4_2_16_r,temp_m4_2_16_i,temp_m4_10_8_r,temp_m4_10_8_i,temp_m4_10_16_r,temp_m4_10_16_i,`W7_real,`W7_imag,`W1_real,`W1_imag,`W8_real,`W8_imag);
butterfly butterfly208 (clk,temp_m4_2_8_r,temp_m4_2_8_i,temp_m4_2_16_r,temp_m4_2_16_i,temp_m4_10_8_r,temp_m4_10_8_i,temp_m4_10_16_r,temp_m4_10_16_i,temp_b4_2_8_r,temp_b4_2_8_i,temp_b4_2_16_r,temp_b4_2_16_i,temp_b4_10_8_r,temp_b4_10_8_i,temp_b4_10_16_r,temp_b4_10_16_i);
MULT MULT209 (clk,temp_b3_3_1_r,temp_b3_3_1_i,temp_b3_3_9_r,temp_b3_3_9_i,temp_b3_11_1_r,temp_b3_11_1_i,temp_b3_11_9_r,temp_b3_11_9_i,temp_m4_3_1_r,temp_m4_3_1_i,temp_m4_3_9_r,temp_m4_3_9_i,temp_m4_11_1_r,temp_m4_11_1_i,temp_m4_11_9_r,temp_m4_11_9_i,`W0_real,`W0_imag,`W2_real,`W2_imag,`W2_real,`W2_imag);
butterfly butterfly209 (clk,temp_m4_3_1_r,temp_m4_3_1_i,temp_m4_3_9_r,temp_m4_3_9_i,temp_m4_11_1_r,temp_m4_11_1_i,temp_m4_11_9_r,temp_m4_11_9_i,temp_b4_3_1_r,temp_b4_3_1_i,temp_b4_3_9_r,temp_b4_3_9_i,temp_b4_11_1_r,temp_b4_11_1_i,temp_b4_11_9_r,temp_b4_11_9_i);
MULT MULT210 (clk,temp_b3_3_2_r,temp_b3_3_2_i,temp_b3_3_10_r,temp_b3_3_10_i,temp_b3_11_2_r,temp_b3_11_2_i,temp_b3_11_10_r,temp_b3_11_10_i,temp_m4_3_2_r,temp_m4_3_2_i,temp_m4_3_10_r,temp_m4_3_10_i,temp_m4_11_2_r,temp_m4_11_2_i,temp_m4_11_10_r,temp_m4_11_10_i,`W1_real,`W1_imag,`W2_real,`W2_imag,`W3_real,`W3_imag);
butterfly butterfly210 (clk,temp_m4_3_2_r,temp_m4_3_2_i,temp_m4_3_10_r,temp_m4_3_10_i,temp_m4_11_2_r,temp_m4_11_2_i,temp_m4_11_10_r,temp_m4_11_10_i,temp_b4_3_2_r,temp_b4_3_2_i,temp_b4_3_10_r,temp_b4_3_10_i,temp_b4_11_2_r,temp_b4_11_2_i,temp_b4_11_10_r,temp_b4_11_10_i);
MULT MULT211 (clk,temp_b3_3_3_r,temp_b3_3_3_i,temp_b3_3_11_r,temp_b3_3_11_i,temp_b3_11_3_r,temp_b3_11_3_i,temp_b3_11_11_r,temp_b3_11_11_i,temp_m4_3_3_r,temp_m4_3_3_i,temp_m4_3_11_r,temp_m4_3_11_i,temp_m4_11_3_r,temp_m4_11_3_i,temp_m4_11_11_r,temp_m4_11_11_i,`W2_real,`W2_imag,`W2_real,`W2_imag,`W4_real,`W4_imag);
butterfly butterfly211 (clk,temp_m4_3_3_r,temp_m4_3_3_i,temp_m4_3_11_r,temp_m4_3_11_i,temp_m4_11_3_r,temp_m4_11_3_i,temp_m4_11_11_r,temp_m4_11_11_i,temp_b4_3_3_r,temp_b4_3_3_i,temp_b4_3_11_r,temp_b4_3_11_i,temp_b4_11_3_r,temp_b4_11_3_i,temp_b4_11_11_r,temp_b4_11_11_i);
MULT MULT212 (clk,temp_b3_3_4_r,temp_b3_3_4_i,temp_b3_3_12_r,temp_b3_3_12_i,temp_b3_11_4_r,temp_b3_11_4_i,temp_b3_11_12_r,temp_b3_11_12_i,temp_m4_3_4_r,temp_m4_3_4_i,temp_m4_3_12_r,temp_m4_3_12_i,temp_m4_11_4_r,temp_m4_11_4_i,temp_m4_11_12_r,temp_m4_11_12_i,`W3_real,`W3_imag,`W2_real,`W2_imag,`W5_real,`W5_imag);
butterfly butterfly212 (clk,temp_m4_3_4_r,temp_m4_3_4_i,temp_m4_3_12_r,temp_m4_3_12_i,temp_m4_11_4_r,temp_m4_11_4_i,temp_m4_11_12_r,temp_m4_11_12_i,temp_b4_3_4_r,temp_b4_3_4_i,temp_b4_3_12_r,temp_b4_3_12_i,temp_b4_11_4_r,temp_b4_11_4_i,temp_b4_11_12_r,temp_b4_11_12_i);
MULT MULT213 (clk,temp_b3_3_5_r,temp_b3_3_5_i,temp_b3_3_13_r,temp_b3_3_13_i,temp_b3_11_5_r,temp_b3_11_5_i,temp_b3_11_13_r,temp_b3_11_13_i,temp_m4_3_5_r,temp_m4_3_5_i,temp_m4_3_13_r,temp_m4_3_13_i,temp_m4_11_5_r,temp_m4_11_5_i,temp_m4_11_13_r,temp_m4_11_13_i,`W4_real,`W4_imag,`W2_real,`W2_imag,`W6_real,`W6_imag);
butterfly butterfly213 (clk,temp_m4_3_5_r,temp_m4_3_5_i,temp_m4_3_13_r,temp_m4_3_13_i,temp_m4_11_5_r,temp_m4_11_5_i,temp_m4_11_13_r,temp_m4_11_13_i,temp_b4_3_5_r,temp_b4_3_5_i,temp_b4_3_13_r,temp_b4_3_13_i,temp_b4_11_5_r,temp_b4_11_5_i,temp_b4_11_13_r,temp_b4_11_13_i);
MULT MULT214 (clk,temp_b3_3_6_r,temp_b3_3_6_i,temp_b3_3_14_r,temp_b3_3_14_i,temp_b3_11_6_r,temp_b3_11_6_i,temp_b3_11_14_r,temp_b3_11_14_i,temp_m4_3_6_r,temp_m4_3_6_i,temp_m4_3_14_r,temp_m4_3_14_i,temp_m4_11_6_r,temp_m4_11_6_i,temp_m4_11_14_r,temp_m4_11_14_i,`W5_real,`W5_imag,`W2_real,`W2_imag,`W7_real,`W7_imag);
butterfly butterfly214 (clk,temp_m4_3_6_r,temp_m4_3_6_i,temp_m4_3_14_r,temp_m4_3_14_i,temp_m4_11_6_r,temp_m4_11_6_i,temp_m4_11_14_r,temp_m4_11_14_i,temp_b4_3_6_r,temp_b4_3_6_i,temp_b4_3_14_r,temp_b4_3_14_i,temp_b4_11_6_r,temp_b4_11_6_i,temp_b4_11_14_r,temp_b4_11_14_i);
MULT MULT215 (clk,temp_b3_3_7_r,temp_b3_3_7_i,temp_b3_3_15_r,temp_b3_3_15_i,temp_b3_11_7_r,temp_b3_11_7_i,temp_b3_11_15_r,temp_b3_11_15_i,temp_m4_3_7_r,temp_m4_3_7_i,temp_m4_3_15_r,temp_m4_3_15_i,temp_m4_11_7_r,temp_m4_11_7_i,temp_m4_11_15_r,temp_m4_11_15_i,`W6_real,`W6_imag,`W2_real,`W2_imag,`W8_real,`W8_imag);
butterfly butterfly215 (clk,temp_m4_3_7_r,temp_m4_3_7_i,temp_m4_3_15_r,temp_m4_3_15_i,temp_m4_11_7_r,temp_m4_11_7_i,temp_m4_11_15_r,temp_m4_11_15_i,temp_b4_3_7_r,temp_b4_3_7_i,temp_b4_3_15_r,temp_b4_3_15_i,temp_b4_11_7_r,temp_b4_11_7_i,temp_b4_11_15_r,temp_b4_11_15_i);
MULT MULT216 (clk,temp_b3_3_8_r,temp_b3_3_8_i,temp_b3_3_16_r,temp_b3_3_16_i,temp_b3_11_8_r,temp_b3_11_8_i,temp_b3_11_16_r,temp_b3_11_16_i,temp_m4_3_8_r,temp_m4_3_8_i,temp_m4_3_16_r,temp_m4_3_16_i,temp_m4_11_8_r,temp_m4_11_8_i,temp_m4_11_16_r,temp_m4_11_16_i,`W7_real,`W7_imag,`W2_real,`W2_imag,`W9_real,`W9_imag);
butterfly butterfly216 (clk,temp_m4_3_8_r,temp_m4_3_8_i,temp_m4_3_16_r,temp_m4_3_16_i,temp_m4_11_8_r,temp_m4_11_8_i,temp_m4_11_16_r,temp_m4_11_16_i,temp_b4_3_8_r,temp_b4_3_8_i,temp_b4_3_16_r,temp_b4_3_16_i,temp_b4_11_8_r,temp_b4_11_8_i,temp_b4_11_16_r,temp_b4_11_16_i);
MULT MULT217 (clk,temp_b3_4_1_r,temp_b3_4_1_i,temp_b3_4_9_r,temp_b3_4_9_i,temp_b3_12_1_r,temp_b3_12_1_i,temp_b3_12_9_r,temp_b3_12_9_i,temp_m4_4_1_r,temp_m4_4_1_i,temp_m4_4_9_r,temp_m4_4_9_i,temp_m4_12_1_r,temp_m4_12_1_i,temp_m4_12_9_r,temp_m4_12_9_i,`W0_real,`W0_imag,`W3_real,`W3_imag,`W3_real,`W3_imag);
butterfly butterfly217 (clk,temp_m4_4_1_r,temp_m4_4_1_i,temp_m4_4_9_r,temp_m4_4_9_i,temp_m4_12_1_r,temp_m4_12_1_i,temp_m4_12_9_r,temp_m4_12_9_i,temp_b4_4_1_r,temp_b4_4_1_i,temp_b4_4_9_r,temp_b4_4_9_i,temp_b4_12_1_r,temp_b4_12_1_i,temp_b4_12_9_r,temp_b4_12_9_i);
MULT MULT218 (clk,temp_b3_4_2_r,temp_b3_4_2_i,temp_b3_4_10_r,temp_b3_4_10_i,temp_b3_12_2_r,temp_b3_12_2_i,temp_b3_12_10_r,temp_b3_12_10_i,temp_m4_4_2_r,temp_m4_4_2_i,temp_m4_4_10_r,temp_m4_4_10_i,temp_m4_12_2_r,temp_m4_12_2_i,temp_m4_12_10_r,temp_m4_12_10_i,`W1_real,`W1_imag,`W3_real,`W3_imag,`W4_real,`W4_imag);
butterfly butterfly218 (clk,temp_m4_4_2_r,temp_m4_4_2_i,temp_m4_4_10_r,temp_m4_4_10_i,temp_m4_12_2_r,temp_m4_12_2_i,temp_m4_12_10_r,temp_m4_12_10_i,temp_b4_4_2_r,temp_b4_4_2_i,temp_b4_4_10_r,temp_b4_4_10_i,temp_b4_12_2_r,temp_b4_12_2_i,temp_b4_12_10_r,temp_b4_12_10_i);
MULT MULT219 (clk,temp_b3_4_3_r,temp_b3_4_3_i,temp_b3_4_11_r,temp_b3_4_11_i,temp_b3_12_3_r,temp_b3_12_3_i,temp_b3_12_11_r,temp_b3_12_11_i,temp_m4_4_3_r,temp_m4_4_3_i,temp_m4_4_11_r,temp_m4_4_11_i,temp_m4_12_3_r,temp_m4_12_3_i,temp_m4_12_11_r,temp_m4_12_11_i,`W2_real,`W2_imag,`W3_real,`W3_imag,`W5_real,`W5_imag);
butterfly butterfly219 (clk,temp_m4_4_3_r,temp_m4_4_3_i,temp_m4_4_11_r,temp_m4_4_11_i,temp_m4_12_3_r,temp_m4_12_3_i,temp_m4_12_11_r,temp_m4_12_11_i,temp_b4_4_3_r,temp_b4_4_3_i,temp_b4_4_11_r,temp_b4_4_11_i,temp_b4_12_3_r,temp_b4_12_3_i,temp_b4_12_11_r,temp_b4_12_11_i);
MULT MULT220 (clk,temp_b3_4_4_r,temp_b3_4_4_i,temp_b3_4_12_r,temp_b3_4_12_i,temp_b3_12_4_r,temp_b3_12_4_i,temp_b3_12_12_r,temp_b3_12_12_i,temp_m4_4_4_r,temp_m4_4_4_i,temp_m4_4_12_r,temp_m4_4_12_i,temp_m4_12_4_r,temp_m4_12_4_i,temp_m4_12_12_r,temp_m4_12_12_i,`W3_real,`W3_imag,`W3_real,`W3_imag,`W6_real,`W6_imag);
butterfly butterfly220 (clk,temp_m4_4_4_r,temp_m4_4_4_i,temp_m4_4_12_r,temp_m4_4_12_i,temp_m4_12_4_r,temp_m4_12_4_i,temp_m4_12_12_r,temp_m4_12_12_i,temp_b4_4_4_r,temp_b4_4_4_i,temp_b4_4_12_r,temp_b4_4_12_i,temp_b4_12_4_r,temp_b4_12_4_i,temp_b4_12_12_r,temp_b4_12_12_i);
MULT MULT221 (clk,temp_b3_4_5_r,temp_b3_4_5_i,temp_b3_4_13_r,temp_b3_4_13_i,temp_b3_12_5_r,temp_b3_12_5_i,temp_b3_12_13_r,temp_b3_12_13_i,temp_m4_4_5_r,temp_m4_4_5_i,temp_m4_4_13_r,temp_m4_4_13_i,temp_m4_12_5_r,temp_m4_12_5_i,temp_m4_12_13_r,temp_m4_12_13_i,`W4_real,`W4_imag,`W3_real,`W3_imag,`W7_real,`W7_imag);
butterfly butterfly221 (clk,temp_m4_4_5_r,temp_m4_4_5_i,temp_m4_4_13_r,temp_m4_4_13_i,temp_m4_12_5_r,temp_m4_12_5_i,temp_m4_12_13_r,temp_m4_12_13_i,temp_b4_4_5_r,temp_b4_4_5_i,temp_b4_4_13_r,temp_b4_4_13_i,temp_b4_12_5_r,temp_b4_12_5_i,temp_b4_12_13_r,temp_b4_12_13_i);
MULT MULT222 (clk,temp_b3_4_6_r,temp_b3_4_6_i,temp_b3_4_14_r,temp_b3_4_14_i,temp_b3_12_6_r,temp_b3_12_6_i,temp_b3_12_14_r,temp_b3_12_14_i,temp_m4_4_6_r,temp_m4_4_6_i,temp_m4_4_14_r,temp_m4_4_14_i,temp_m4_12_6_r,temp_m4_12_6_i,temp_m4_12_14_r,temp_m4_12_14_i,`W5_real,`W5_imag,`W3_real,`W3_imag,`W8_real,`W8_imag);
butterfly butterfly222 (clk,temp_m4_4_6_r,temp_m4_4_6_i,temp_m4_4_14_r,temp_m4_4_14_i,temp_m4_12_6_r,temp_m4_12_6_i,temp_m4_12_14_r,temp_m4_12_14_i,temp_b4_4_6_r,temp_b4_4_6_i,temp_b4_4_14_r,temp_b4_4_14_i,temp_b4_12_6_r,temp_b4_12_6_i,temp_b4_12_14_r,temp_b4_12_14_i);
MULT MULT223 (clk,temp_b3_4_7_r,temp_b3_4_7_i,temp_b3_4_15_r,temp_b3_4_15_i,temp_b3_12_7_r,temp_b3_12_7_i,temp_b3_12_15_r,temp_b3_12_15_i,temp_m4_4_7_r,temp_m4_4_7_i,temp_m4_4_15_r,temp_m4_4_15_i,temp_m4_12_7_r,temp_m4_12_7_i,temp_m4_12_15_r,temp_m4_12_15_i,`W6_real,`W6_imag,`W3_real,`W3_imag,`W9_real,`W9_imag);
butterfly butterfly223 (clk,temp_m4_4_7_r,temp_m4_4_7_i,temp_m4_4_15_r,temp_m4_4_15_i,temp_m4_12_7_r,temp_m4_12_7_i,temp_m4_12_15_r,temp_m4_12_15_i,temp_b4_4_7_r,temp_b4_4_7_i,temp_b4_4_15_r,temp_b4_4_15_i,temp_b4_12_7_r,temp_b4_12_7_i,temp_b4_12_15_r,temp_b4_12_15_i);
MULT MULT224 (clk,temp_b3_4_8_r,temp_b3_4_8_i,temp_b3_4_16_r,temp_b3_4_16_i,temp_b3_12_8_r,temp_b3_12_8_i,temp_b3_12_16_r,temp_b3_12_16_i,temp_m4_4_8_r,temp_m4_4_8_i,temp_m4_4_16_r,temp_m4_4_16_i,temp_m4_12_8_r,temp_m4_12_8_i,temp_m4_12_16_r,temp_m4_12_16_i,`W7_real,`W7_imag,`W3_real,`W3_imag,`W10_real,`W10_imag);
butterfly butterfly224 (clk,temp_m4_4_8_r,temp_m4_4_8_i,temp_m4_4_16_r,temp_m4_4_16_i,temp_m4_12_8_r,temp_m4_12_8_i,temp_m4_12_16_r,temp_m4_12_16_i,temp_b4_4_8_r,temp_b4_4_8_i,temp_b4_4_16_r,temp_b4_4_16_i,temp_b4_12_8_r,temp_b4_12_8_i,temp_b4_12_16_r,temp_b4_12_16_i);
MULT MULT225 (clk,temp_b3_5_1_r,temp_b3_5_1_i,temp_b3_5_9_r,temp_b3_5_9_i,temp_b3_13_1_r,temp_b3_13_1_i,temp_b3_13_9_r,temp_b3_13_9_i,temp_m4_5_1_r,temp_m4_5_1_i,temp_m4_5_9_r,temp_m4_5_9_i,temp_m4_13_1_r,temp_m4_13_1_i,temp_m4_13_9_r,temp_m4_13_9_i,`W0_real,`W0_imag,`W4_real,`W4_imag,`W4_real,`W4_imag);
butterfly butterfly225 (clk,temp_m4_5_1_r,temp_m4_5_1_i,temp_m4_5_9_r,temp_m4_5_9_i,temp_m4_13_1_r,temp_m4_13_1_i,temp_m4_13_9_r,temp_m4_13_9_i,temp_b4_5_1_r,temp_b4_5_1_i,temp_b4_5_9_r,temp_b4_5_9_i,temp_b4_13_1_r,temp_b4_13_1_i,temp_b4_13_9_r,temp_b4_13_9_i);
MULT MULT226 (clk,temp_b3_5_2_r,temp_b3_5_2_i,temp_b3_5_10_r,temp_b3_5_10_i,temp_b3_13_2_r,temp_b3_13_2_i,temp_b3_13_10_r,temp_b3_13_10_i,temp_m4_5_2_r,temp_m4_5_2_i,temp_m4_5_10_r,temp_m4_5_10_i,temp_m4_13_2_r,temp_m4_13_2_i,temp_m4_13_10_r,temp_m4_13_10_i,`W1_real,`W1_imag,`W4_real,`W4_imag,`W5_real,`W5_imag);
butterfly butterfly226 (clk,temp_m4_5_2_r,temp_m4_5_2_i,temp_m4_5_10_r,temp_m4_5_10_i,temp_m4_13_2_r,temp_m4_13_2_i,temp_m4_13_10_r,temp_m4_13_10_i,temp_b4_5_2_r,temp_b4_5_2_i,temp_b4_5_10_r,temp_b4_5_10_i,temp_b4_13_2_r,temp_b4_13_2_i,temp_b4_13_10_r,temp_b4_13_10_i);
MULT MULT227 (clk,temp_b3_5_3_r,temp_b3_5_3_i,temp_b3_5_11_r,temp_b3_5_11_i,temp_b3_13_3_r,temp_b3_13_3_i,temp_b3_13_11_r,temp_b3_13_11_i,temp_m4_5_3_r,temp_m4_5_3_i,temp_m4_5_11_r,temp_m4_5_11_i,temp_m4_13_3_r,temp_m4_13_3_i,temp_m4_13_11_r,temp_m4_13_11_i,`W2_real,`W2_imag,`W4_real,`W4_imag,`W6_real,`W6_imag);
butterfly butterfly227 (clk,temp_m4_5_3_r,temp_m4_5_3_i,temp_m4_5_11_r,temp_m4_5_11_i,temp_m4_13_3_r,temp_m4_13_3_i,temp_m4_13_11_r,temp_m4_13_11_i,temp_b4_5_3_r,temp_b4_5_3_i,temp_b4_5_11_r,temp_b4_5_11_i,temp_b4_13_3_r,temp_b4_13_3_i,temp_b4_13_11_r,temp_b4_13_11_i);
MULT MULT228 (clk,temp_b3_5_4_r,temp_b3_5_4_i,temp_b3_5_12_r,temp_b3_5_12_i,temp_b3_13_4_r,temp_b3_13_4_i,temp_b3_13_12_r,temp_b3_13_12_i,temp_m4_5_4_r,temp_m4_5_4_i,temp_m4_5_12_r,temp_m4_5_12_i,temp_m4_13_4_r,temp_m4_13_4_i,temp_m4_13_12_r,temp_m4_13_12_i,`W3_real,`W3_imag,`W4_real,`W4_imag,`W7_real,`W7_imag);
butterfly butterfly228 (clk,temp_m4_5_4_r,temp_m4_5_4_i,temp_m4_5_12_r,temp_m4_5_12_i,temp_m4_13_4_r,temp_m4_13_4_i,temp_m4_13_12_r,temp_m4_13_12_i,temp_b4_5_4_r,temp_b4_5_4_i,temp_b4_5_12_r,temp_b4_5_12_i,temp_b4_13_4_r,temp_b4_13_4_i,temp_b4_13_12_r,temp_b4_13_12_i);
MULT MULT229 (clk,temp_b3_5_5_r,temp_b3_5_5_i,temp_b3_5_13_r,temp_b3_5_13_i,temp_b3_13_5_r,temp_b3_13_5_i,temp_b3_13_13_r,temp_b3_13_13_i,temp_m4_5_5_r,temp_m4_5_5_i,temp_m4_5_13_r,temp_m4_5_13_i,temp_m4_13_5_r,temp_m4_13_5_i,temp_m4_13_13_r,temp_m4_13_13_i,`W4_real,`W4_imag,`W4_real,`W4_imag,`W8_real,`W8_imag);
butterfly butterfly229 (clk,temp_m4_5_5_r,temp_m4_5_5_i,temp_m4_5_13_r,temp_m4_5_13_i,temp_m4_13_5_r,temp_m4_13_5_i,temp_m4_13_13_r,temp_m4_13_13_i,temp_b4_5_5_r,temp_b4_5_5_i,temp_b4_5_13_r,temp_b4_5_13_i,temp_b4_13_5_r,temp_b4_13_5_i,temp_b4_13_13_r,temp_b4_13_13_i);
MULT MULT230 (clk,temp_b3_5_6_r,temp_b3_5_6_i,temp_b3_5_14_r,temp_b3_5_14_i,temp_b3_13_6_r,temp_b3_13_6_i,temp_b3_13_14_r,temp_b3_13_14_i,temp_m4_5_6_r,temp_m4_5_6_i,temp_m4_5_14_r,temp_m4_5_14_i,temp_m4_13_6_r,temp_m4_13_6_i,temp_m4_13_14_r,temp_m4_13_14_i,`W5_real,`W5_imag,`W4_real,`W4_imag,`W9_real,`W9_imag);
butterfly butterfly230 (clk,temp_m4_5_6_r,temp_m4_5_6_i,temp_m4_5_14_r,temp_m4_5_14_i,temp_m4_13_6_r,temp_m4_13_6_i,temp_m4_13_14_r,temp_m4_13_14_i,temp_b4_5_6_r,temp_b4_5_6_i,temp_b4_5_14_r,temp_b4_5_14_i,temp_b4_13_6_r,temp_b4_13_6_i,temp_b4_13_14_r,temp_b4_13_14_i);
MULT MULT231 (clk,temp_b3_5_7_r,temp_b3_5_7_i,temp_b3_5_15_r,temp_b3_5_15_i,temp_b3_13_7_r,temp_b3_13_7_i,temp_b3_13_15_r,temp_b3_13_15_i,temp_m4_5_7_r,temp_m4_5_7_i,temp_m4_5_15_r,temp_m4_5_15_i,temp_m4_13_7_r,temp_m4_13_7_i,temp_m4_13_15_r,temp_m4_13_15_i,`W6_real,`W6_imag,`W4_real,`W4_imag,`W10_real,`W10_imag);
butterfly butterfly231 (clk,temp_m4_5_7_r,temp_m4_5_7_i,temp_m4_5_15_r,temp_m4_5_15_i,temp_m4_13_7_r,temp_m4_13_7_i,temp_m4_13_15_r,temp_m4_13_15_i,temp_b4_5_7_r,temp_b4_5_7_i,temp_b4_5_15_r,temp_b4_5_15_i,temp_b4_13_7_r,temp_b4_13_7_i,temp_b4_13_15_r,temp_b4_13_15_i);
MULT MULT232 (clk,temp_b3_5_8_r,temp_b3_5_8_i,temp_b3_5_16_r,temp_b3_5_16_i,temp_b3_13_8_r,temp_b3_13_8_i,temp_b3_13_16_r,temp_b3_13_16_i,temp_m4_5_8_r,temp_m4_5_8_i,temp_m4_5_16_r,temp_m4_5_16_i,temp_m4_13_8_r,temp_m4_13_8_i,temp_m4_13_16_r,temp_m4_13_16_i,`W7_real,`W7_imag,`W4_real,`W4_imag,`W11_real,`W11_imag);
butterfly butterfly232 (clk,temp_m4_5_8_r,temp_m4_5_8_i,temp_m4_5_16_r,temp_m4_5_16_i,temp_m4_13_8_r,temp_m4_13_8_i,temp_m4_13_16_r,temp_m4_13_16_i,temp_b4_5_8_r,temp_b4_5_8_i,temp_b4_5_16_r,temp_b4_5_16_i,temp_b4_13_8_r,temp_b4_13_8_i,temp_b4_13_16_r,temp_b4_13_16_i);
MULT MULT233 (clk,temp_b3_6_1_r,temp_b3_6_1_i,temp_b3_6_9_r,temp_b3_6_9_i,temp_b3_14_1_r,temp_b3_14_1_i,temp_b3_14_9_r,temp_b3_14_9_i,temp_m4_6_1_r,temp_m4_6_1_i,temp_m4_6_9_r,temp_m4_6_9_i,temp_m4_14_1_r,temp_m4_14_1_i,temp_m4_14_9_r,temp_m4_14_9_i,`W0_real,`W0_imag,`W5_real,`W5_imag,`W5_real,`W5_imag);
butterfly butterfly233 (clk,temp_m4_6_1_r,temp_m4_6_1_i,temp_m4_6_9_r,temp_m4_6_9_i,temp_m4_14_1_r,temp_m4_14_1_i,temp_m4_14_9_r,temp_m4_14_9_i,temp_b4_6_1_r,temp_b4_6_1_i,temp_b4_6_9_r,temp_b4_6_9_i,temp_b4_14_1_r,temp_b4_14_1_i,temp_b4_14_9_r,temp_b4_14_9_i);
MULT MULT234 (clk,temp_b3_6_2_r,temp_b3_6_2_i,temp_b3_6_10_r,temp_b3_6_10_i,temp_b3_14_2_r,temp_b3_14_2_i,temp_b3_14_10_r,temp_b3_14_10_i,temp_m4_6_2_r,temp_m4_6_2_i,temp_m4_6_10_r,temp_m4_6_10_i,temp_m4_14_2_r,temp_m4_14_2_i,temp_m4_14_10_r,temp_m4_14_10_i,`W1_real,`W1_imag,`W5_real,`W5_imag,`W6_real,`W6_imag);
butterfly butterfly234 (clk,temp_m4_6_2_r,temp_m4_6_2_i,temp_m4_6_10_r,temp_m4_6_10_i,temp_m4_14_2_r,temp_m4_14_2_i,temp_m4_14_10_r,temp_m4_14_10_i,temp_b4_6_2_r,temp_b4_6_2_i,temp_b4_6_10_r,temp_b4_6_10_i,temp_b4_14_2_r,temp_b4_14_2_i,temp_b4_14_10_r,temp_b4_14_10_i);
MULT MULT235 (clk,temp_b3_6_3_r,temp_b3_6_3_i,temp_b3_6_11_r,temp_b3_6_11_i,temp_b3_14_3_r,temp_b3_14_3_i,temp_b3_14_11_r,temp_b3_14_11_i,temp_m4_6_3_r,temp_m4_6_3_i,temp_m4_6_11_r,temp_m4_6_11_i,temp_m4_14_3_r,temp_m4_14_3_i,temp_m4_14_11_r,temp_m4_14_11_i,`W2_real,`W2_imag,`W5_real,`W5_imag,`W7_real,`W7_imag);
butterfly butterfly235 (clk,temp_m4_6_3_r,temp_m4_6_3_i,temp_m4_6_11_r,temp_m4_6_11_i,temp_m4_14_3_r,temp_m4_14_3_i,temp_m4_14_11_r,temp_m4_14_11_i,temp_b4_6_3_r,temp_b4_6_3_i,temp_b4_6_11_r,temp_b4_6_11_i,temp_b4_14_3_r,temp_b4_14_3_i,temp_b4_14_11_r,temp_b4_14_11_i);
MULT MULT236 (clk,temp_b3_6_4_r,temp_b3_6_4_i,temp_b3_6_12_r,temp_b3_6_12_i,temp_b3_14_4_r,temp_b3_14_4_i,temp_b3_14_12_r,temp_b3_14_12_i,temp_m4_6_4_r,temp_m4_6_4_i,temp_m4_6_12_r,temp_m4_6_12_i,temp_m4_14_4_r,temp_m4_14_4_i,temp_m4_14_12_r,temp_m4_14_12_i,`W3_real,`W3_imag,`W5_real,`W5_imag,`W8_real,`W8_imag);
butterfly butterfly236 (clk,temp_m4_6_4_r,temp_m4_6_4_i,temp_m4_6_12_r,temp_m4_6_12_i,temp_m4_14_4_r,temp_m4_14_4_i,temp_m4_14_12_r,temp_m4_14_12_i,temp_b4_6_4_r,temp_b4_6_4_i,temp_b4_6_12_r,temp_b4_6_12_i,temp_b4_14_4_r,temp_b4_14_4_i,temp_b4_14_12_r,temp_b4_14_12_i);
MULT MULT237 (clk,temp_b3_6_5_r,temp_b3_6_5_i,temp_b3_6_13_r,temp_b3_6_13_i,temp_b3_14_5_r,temp_b3_14_5_i,temp_b3_14_13_r,temp_b3_14_13_i,temp_m4_6_5_r,temp_m4_6_5_i,temp_m4_6_13_r,temp_m4_6_13_i,temp_m4_14_5_r,temp_m4_14_5_i,temp_m4_14_13_r,temp_m4_14_13_i,`W4_real,`W4_imag,`W5_real,`W5_imag,`W9_real,`W9_imag);
butterfly butterfly237 (clk,temp_m4_6_5_r,temp_m4_6_5_i,temp_m4_6_13_r,temp_m4_6_13_i,temp_m4_14_5_r,temp_m4_14_5_i,temp_m4_14_13_r,temp_m4_14_13_i,temp_b4_6_5_r,temp_b4_6_5_i,temp_b4_6_13_r,temp_b4_6_13_i,temp_b4_14_5_r,temp_b4_14_5_i,temp_b4_14_13_r,temp_b4_14_13_i);
MULT MULT238 (clk,temp_b3_6_6_r,temp_b3_6_6_i,temp_b3_6_14_r,temp_b3_6_14_i,temp_b3_14_6_r,temp_b3_14_6_i,temp_b3_14_14_r,temp_b3_14_14_i,temp_m4_6_6_r,temp_m4_6_6_i,temp_m4_6_14_r,temp_m4_6_14_i,temp_m4_14_6_r,temp_m4_14_6_i,temp_m4_14_14_r,temp_m4_14_14_i,`W5_real,`W5_imag,`W5_real,`W5_imag,`W10_real,`W10_imag);
butterfly butterfly238 (clk,temp_m4_6_6_r,temp_m4_6_6_i,temp_m4_6_14_r,temp_m4_6_14_i,temp_m4_14_6_r,temp_m4_14_6_i,temp_m4_14_14_r,temp_m4_14_14_i,temp_b4_6_6_r,temp_b4_6_6_i,temp_b4_6_14_r,temp_b4_6_14_i,temp_b4_14_6_r,temp_b4_14_6_i,temp_b4_14_14_r,temp_b4_14_14_i);
MULT MULT239 (clk,temp_b3_6_7_r,temp_b3_6_7_i,temp_b3_6_15_r,temp_b3_6_15_i,temp_b3_14_7_r,temp_b3_14_7_i,temp_b3_14_15_r,temp_b3_14_15_i,temp_m4_6_7_r,temp_m4_6_7_i,temp_m4_6_15_r,temp_m4_6_15_i,temp_m4_14_7_r,temp_m4_14_7_i,temp_m4_14_15_r,temp_m4_14_15_i,`W6_real,`W6_imag,`W5_real,`W5_imag,`W11_real,`W11_imag);
butterfly butterfly239 (clk,temp_m4_6_7_r,temp_m4_6_7_i,temp_m4_6_15_r,temp_m4_6_15_i,temp_m4_14_7_r,temp_m4_14_7_i,temp_m4_14_15_r,temp_m4_14_15_i,temp_b4_6_7_r,temp_b4_6_7_i,temp_b4_6_15_r,temp_b4_6_15_i,temp_b4_14_7_r,temp_b4_14_7_i,temp_b4_14_15_r,temp_b4_14_15_i);
MULT MULT240 (clk,temp_b3_6_8_r,temp_b3_6_8_i,temp_b3_6_16_r,temp_b3_6_16_i,temp_b3_14_8_r,temp_b3_14_8_i,temp_b3_14_16_r,temp_b3_14_16_i,temp_m4_6_8_r,temp_m4_6_8_i,temp_m4_6_16_r,temp_m4_6_16_i,temp_m4_14_8_r,temp_m4_14_8_i,temp_m4_14_16_r,temp_m4_14_16_i,`W7_real,`W7_imag,`W5_real,`W5_imag,`W12_real,`W12_imag);
butterfly butterfly240 (clk,temp_m4_6_8_r,temp_m4_6_8_i,temp_m4_6_16_r,temp_m4_6_16_i,temp_m4_14_8_r,temp_m4_14_8_i,temp_m4_14_16_r,temp_m4_14_16_i,temp_b4_6_8_r,temp_b4_6_8_i,temp_b4_6_16_r,temp_b4_6_16_i,temp_b4_14_8_r,temp_b4_14_8_i,temp_b4_14_16_r,temp_b4_14_16_i);
MULT MULT241 (clk,temp_b3_7_1_r,temp_b3_7_1_i,temp_b3_7_9_r,temp_b3_7_9_i,temp_b3_15_1_r,temp_b3_15_1_i,temp_b3_15_9_r,temp_b3_15_9_i,temp_m4_7_1_r,temp_m4_7_1_i,temp_m4_7_9_r,temp_m4_7_9_i,temp_m4_15_1_r,temp_m4_15_1_i,temp_m4_15_9_r,temp_m4_15_9_i,`W0_real,`W0_imag,`W6_real,`W6_imag,`W6_real,`W6_imag);
butterfly butterfly241 (clk,temp_m4_7_1_r,temp_m4_7_1_i,temp_m4_7_9_r,temp_m4_7_9_i,temp_m4_15_1_r,temp_m4_15_1_i,temp_m4_15_9_r,temp_m4_15_9_i,temp_b4_7_1_r,temp_b4_7_1_i,temp_b4_7_9_r,temp_b4_7_9_i,temp_b4_15_1_r,temp_b4_15_1_i,temp_b4_15_9_r,temp_b4_15_9_i);
MULT MULT242 (clk,temp_b3_7_2_r,temp_b3_7_2_i,temp_b3_7_10_r,temp_b3_7_10_i,temp_b3_15_2_r,temp_b3_15_2_i,temp_b3_15_10_r,temp_b3_15_10_i,temp_m4_7_2_r,temp_m4_7_2_i,temp_m4_7_10_r,temp_m4_7_10_i,temp_m4_15_2_r,temp_m4_15_2_i,temp_m4_15_10_r,temp_m4_15_10_i,`W1_real,`W1_imag,`W6_real,`W6_imag,`W7_real,`W7_imag);
butterfly butterfly242 (clk,temp_m4_7_2_r,temp_m4_7_2_i,temp_m4_7_10_r,temp_m4_7_10_i,temp_m4_15_2_r,temp_m4_15_2_i,temp_m4_15_10_r,temp_m4_15_10_i,temp_b4_7_2_r,temp_b4_7_2_i,temp_b4_7_10_r,temp_b4_7_10_i,temp_b4_15_2_r,temp_b4_15_2_i,temp_b4_15_10_r,temp_b4_15_10_i);
MULT MULT243 (clk,temp_b3_7_3_r,temp_b3_7_3_i,temp_b3_7_11_r,temp_b3_7_11_i,temp_b3_15_3_r,temp_b3_15_3_i,temp_b3_15_11_r,temp_b3_15_11_i,temp_m4_7_3_r,temp_m4_7_3_i,temp_m4_7_11_r,temp_m4_7_11_i,temp_m4_15_3_r,temp_m4_15_3_i,temp_m4_15_11_r,temp_m4_15_11_i,`W2_real,`W2_imag,`W6_real,`W6_imag,`W8_real,`W8_imag);
butterfly butterfly243 (clk,temp_m4_7_3_r,temp_m4_7_3_i,temp_m4_7_11_r,temp_m4_7_11_i,temp_m4_15_3_r,temp_m4_15_3_i,temp_m4_15_11_r,temp_m4_15_11_i,temp_b4_7_3_r,temp_b4_7_3_i,temp_b4_7_11_r,temp_b4_7_11_i,temp_b4_15_3_r,temp_b4_15_3_i,temp_b4_15_11_r,temp_b4_15_11_i);
MULT MULT244 (clk,temp_b3_7_4_r,temp_b3_7_4_i,temp_b3_7_12_r,temp_b3_7_12_i,temp_b3_15_4_r,temp_b3_15_4_i,temp_b3_15_12_r,temp_b3_15_12_i,temp_m4_7_4_r,temp_m4_7_4_i,temp_m4_7_12_r,temp_m4_7_12_i,temp_m4_15_4_r,temp_m4_15_4_i,temp_m4_15_12_r,temp_m4_15_12_i,`W3_real,`W3_imag,`W6_real,`W6_imag,`W9_real,`W9_imag);
butterfly butterfly244 (clk,temp_m4_7_4_r,temp_m4_7_4_i,temp_m4_7_12_r,temp_m4_7_12_i,temp_m4_15_4_r,temp_m4_15_4_i,temp_m4_15_12_r,temp_m4_15_12_i,temp_b4_7_4_r,temp_b4_7_4_i,temp_b4_7_12_r,temp_b4_7_12_i,temp_b4_15_4_r,temp_b4_15_4_i,temp_b4_15_12_r,temp_b4_15_12_i);
MULT MULT245 (clk,temp_b3_7_5_r,temp_b3_7_5_i,temp_b3_7_13_r,temp_b3_7_13_i,temp_b3_15_5_r,temp_b3_15_5_i,temp_b3_15_13_r,temp_b3_15_13_i,temp_m4_7_5_r,temp_m4_7_5_i,temp_m4_7_13_r,temp_m4_7_13_i,temp_m4_15_5_r,temp_m4_15_5_i,temp_m4_15_13_r,temp_m4_15_13_i,`W4_real,`W4_imag,`W6_real,`W6_imag,`W10_real,`W10_imag);
butterfly butterfly245 (clk,temp_m4_7_5_r,temp_m4_7_5_i,temp_m4_7_13_r,temp_m4_7_13_i,temp_m4_15_5_r,temp_m4_15_5_i,temp_m4_15_13_r,temp_m4_15_13_i,temp_b4_7_5_r,temp_b4_7_5_i,temp_b4_7_13_r,temp_b4_7_13_i,temp_b4_15_5_r,temp_b4_15_5_i,temp_b4_15_13_r,temp_b4_15_13_i);
MULT MULT246 (clk,temp_b3_7_6_r,temp_b3_7_6_i,temp_b3_7_14_r,temp_b3_7_14_i,temp_b3_15_6_r,temp_b3_15_6_i,temp_b3_15_14_r,temp_b3_15_14_i,temp_m4_7_6_r,temp_m4_7_6_i,temp_m4_7_14_r,temp_m4_7_14_i,temp_m4_15_6_r,temp_m4_15_6_i,temp_m4_15_14_r,temp_m4_15_14_i,`W5_real,`W5_imag,`W6_real,`W6_imag,`W11_real,`W11_imag);
butterfly butterfly246 (clk,temp_m4_7_6_r,temp_m4_7_6_i,temp_m4_7_14_r,temp_m4_7_14_i,temp_m4_15_6_r,temp_m4_15_6_i,temp_m4_15_14_r,temp_m4_15_14_i,temp_b4_7_6_r,temp_b4_7_6_i,temp_b4_7_14_r,temp_b4_7_14_i,temp_b4_15_6_r,temp_b4_15_6_i,temp_b4_15_14_r,temp_b4_15_14_i);
MULT MULT247 (clk,temp_b3_7_7_r,temp_b3_7_7_i,temp_b3_7_15_r,temp_b3_7_15_i,temp_b3_15_7_r,temp_b3_15_7_i,temp_b3_15_15_r,temp_b3_15_15_i,temp_m4_7_7_r,temp_m4_7_7_i,temp_m4_7_15_r,temp_m4_7_15_i,temp_m4_15_7_r,temp_m4_15_7_i,temp_m4_15_15_r,temp_m4_15_15_i,`W6_real,`W6_imag,`W6_real,`W6_imag,`W12_real,`W12_imag);
butterfly butterfly247 (clk,temp_m4_7_7_r,temp_m4_7_7_i,temp_m4_7_15_r,temp_m4_7_15_i,temp_m4_15_7_r,temp_m4_15_7_i,temp_m4_15_15_r,temp_m4_15_15_i,temp_b4_7_7_r,temp_b4_7_7_i,temp_b4_7_15_r,temp_b4_7_15_i,temp_b4_15_7_r,temp_b4_15_7_i,temp_b4_15_15_r,temp_b4_15_15_i);
MULT MULT248 (clk,temp_b3_7_8_r,temp_b3_7_8_i,temp_b3_7_16_r,temp_b3_7_16_i,temp_b3_15_8_r,temp_b3_15_8_i,temp_b3_15_16_r,temp_b3_15_16_i,temp_m4_7_8_r,temp_m4_7_8_i,temp_m4_7_16_r,temp_m4_7_16_i,temp_m4_15_8_r,temp_m4_15_8_i,temp_m4_15_16_r,temp_m4_15_16_i,`W7_real,`W7_imag,`W6_real,`W6_imag,`W13_real,`W13_imag);
butterfly butterfly248 (clk,temp_m4_7_8_r,temp_m4_7_8_i,temp_m4_7_16_r,temp_m4_7_16_i,temp_m4_15_8_r,temp_m4_15_8_i,temp_m4_15_16_r,temp_m4_15_16_i,temp_b4_7_8_r,temp_b4_7_8_i,temp_b4_7_16_r,temp_b4_7_16_i,temp_b4_15_8_r,temp_b4_15_8_i,temp_b4_15_16_r,temp_b4_15_16_i);
MULT MULT249 (clk,temp_b3_8_1_r,temp_b3_8_1_i,temp_b3_8_9_r,temp_b3_8_9_i,temp_b3_16_1_r,temp_b3_16_1_i,temp_b3_16_9_r,temp_b3_16_9_i,temp_m4_8_1_r,temp_m4_8_1_i,temp_m4_8_9_r,temp_m4_8_9_i,temp_m4_16_1_r,temp_m4_16_1_i,temp_m4_16_9_r,temp_m4_16_9_i,`W0_real,`W0_imag,`W7_real,`W7_imag,`W7_real,`W7_imag);
butterfly butterfly249 (clk,temp_m4_8_1_r,temp_m4_8_1_i,temp_m4_8_9_r,temp_m4_8_9_i,temp_m4_16_1_r,temp_m4_16_1_i,temp_m4_16_9_r,temp_m4_16_9_i,temp_b4_8_1_r,temp_b4_8_1_i,temp_b4_8_9_r,temp_b4_8_9_i,temp_b4_16_1_r,temp_b4_16_1_i,temp_b4_16_9_r,temp_b4_16_9_i);
MULT MULT250 (clk,temp_b3_8_2_r,temp_b3_8_2_i,temp_b3_8_10_r,temp_b3_8_10_i,temp_b3_16_2_r,temp_b3_16_2_i,temp_b3_16_10_r,temp_b3_16_10_i,temp_m4_8_2_r,temp_m4_8_2_i,temp_m4_8_10_r,temp_m4_8_10_i,temp_m4_16_2_r,temp_m4_16_2_i,temp_m4_16_10_r,temp_m4_16_10_i,`W1_real,`W1_imag,`W7_real,`W7_imag,`W8_real,`W8_imag);
butterfly butterfly250 (clk,temp_m4_8_2_r,temp_m4_8_2_i,temp_m4_8_10_r,temp_m4_8_10_i,temp_m4_16_2_r,temp_m4_16_2_i,temp_m4_16_10_r,temp_m4_16_10_i,temp_b4_8_2_r,temp_b4_8_2_i,temp_b4_8_10_r,temp_b4_8_10_i,temp_b4_16_2_r,temp_b4_16_2_i,temp_b4_16_10_r,temp_b4_16_10_i);
MULT MULT251 (clk,temp_b3_8_3_r,temp_b3_8_3_i,temp_b3_8_11_r,temp_b3_8_11_i,temp_b3_16_3_r,temp_b3_16_3_i,temp_b3_16_11_r,temp_b3_16_11_i,temp_m4_8_3_r,temp_m4_8_3_i,temp_m4_8_11_r,temp_m4_8_11_i,temp_m4_16_3_r,temp_m4_16_3_i,temp_m4_16_11_r,temp_m4_16_11_i,`W2_real,`W2_imag,`W7_real,`W7_imag,`W9_real,`W9_imag);
butterfly butterfly251 (clk,temp_m4_8_3_r,temp_m4_8_3_i,temp_m4_8_11_r,temp_m4_8_11_i,temp_m4_16_3_r,temp_m4_16_3_i,temp_m4_16_11_r,temp_m4_16_11_i,temp_b4_8_3_r,temp_b4_8_3_i,temp_b4_8_11_r,temp_b4_8_11_i,temp_b4_16_3_r,temp_b4_16_3_i,temp_b4_16_11_r,temp_b4_16_11_i);
MULT MULT252 (clk,temp_b3_8_4_r,temp_b3_8_4_i,temp_b3_8_12_r,temp_b3_8_12_i,temp_b3_16_4_r,temp_b3_16_4_i,temp_b3_16_12_r,temp_b3_16_12_i,temp_m4_8_4_r,temp_m4_8_4_i,temp_m4_8_12_r,temp_m4_8_12_i,temp_m4_16_4_r,temp_m4_16_4_i,temp_m4_16_12_r,temp_m4_16_12_i,`W3_real,`W3_imag,`W7_real,`W7_imag,`W10_real,`W10_imag);
butterfly butterfly252 (clk,temp_m4_8_4_r,temp_m4_8_4_i,temp_m4_8_12_r,temp_m4_8_12_i,temp_m4_16_4_r,temp_m4_16_4_i,temp_m4_16_12_r,temp_m4_16_12_i,temp_b4_8_4_r,temp_b4_8_4_i,temp_b4_8_12_r,temp_b4_8_12_i,temp_b4_16_4_r,temp_b4_16_4_i,temp_b4_16_12_r,temp_b4_16_12_i);
MULT MULT253 (clk,temp_b3_8_5_r,temp_b3_8_5_i,temp_b3_8_13_r,temp_b3_8_13_i,temp_b3_16_5_r,temp_b3_16_5_i,temp_b3_16_13_r,temp_b3_16_13_i,temp_m4_8_5_r,temp_m4_8_5_i,temp_m4_8_13_r,temp_m4_8_13_i,temp_m4_16_5_r,temp_m4_16_5_i,temp_m4_16_13_r,temp_m4_16_13_i,`W4_real,`W4_imag,`W7_real,`W7_imag,`W11_real,`W11_imag);
butterfly butterfly253 (clk,temp_m4_8_5_r,temp_m4_8_5_i,temp_m4_8_13_r,temp_m4_8_13_i,temp_m4_16_5_r,temp_m4_16_5_i,temp_m4_16_13_r,temp_m4_16_13_i,temp_b4_8_5_r,temp_b4_8_5_i,temp_b4_8_13_r,temp_b4_8_13_i,temp_b4_16_5_r,temp_b4_16_5_i,temp_b4_16_13_r,temp_b4_16_13_i);
MULT MULT254 (clk,temp_b3_8_6_r,temp_b3_8_6_i,temp_b3_8_14_r,temp_b3_8_14_i,temp_b3_16_6_r,temp_b3_16_6_i,temp_b3_16_14_r,temp_b3_16_14_i,temp_m4_8_6_r,temp_m4_8_6_i,temp_m4_8_14_r,temp_m4_8_14_i,temp_m4_16_6_r,temp_m4_16_6_i,temp_m4_16_14_r,temp_m4_16_14_i,`W5_real,`W5_imag,`W7_real,`W7_imag,`W12_real,`W12_imag);
butterfly butterfly254 (clk,temp_m4_8_6_r,temp_m4_8_6_i,temp_m4_8_14_r,temp_m4_8_14_i,temp_m4_16_6_r,temp_m4_16_6_i,temp_m4_16_14_r,temp_m4_16_14_i,temp_b4_8_6_r,temp_b4_8_6_i,temp_b4_8_14_r,temp_b4_8_14_i,temp_b4_16_6_r,temp_b4_16_6_i,temp_b4_16_14_r,temp_b4_16_14_i);
MULT MULT255 (clk,temp_b3_8_7_r,temp_b3_8_7_i,temp_b3_8_15_r,temp_b3_8_15_i,temp_b3_16_7_r,temp_b3_16_7_i,temp_b3_16_15_r,temp_b3_16_15_i,temp_m4_8_7_r,temp_m4_8_7_i,temp_m4_8_15_r,temp_m4_8_15_i,temp_m4_16_7_r,temp_m4_16_7_i,temp_m4_16_15_r,temp_m4_16_15_i,`W6_real,`W6_imag,`W7_real,`W7_imag,`W13_real,`W13_imag);
butterfly butterfly255 (clk,temp_m4_8_7_r,temp_m4_8_7_i,temp_m4_8_15_r,temp_m4_8_15_i,temp_m4_16_7_r,temp_m4_16_7_i,temp_m4_16_15_r,temp_m4_16_15_i,temp_b4_8_7_r,temp_b4_8_7_i,temp_b4_8_15_r,temp_b4_8_15_i,temp_b4_16_7_r,temp_b4_16_7_i,temp_b4_16_15_r,temp_b4_16_15_i);
MULT MULT256 (clk,temp_b3_8_8_r,temp_b3_8_8_i,temp_b3_8_16_r,temp_b3_8_16_i,temp_b3_16_8_r,temp_b3_16_8_i,temp_b3_16_16_r,temp_b3_16_16_i,temp_m4_8_8_r,temp_m4_8_8_i,temp_m4_8_16_r,temp_m4_8_16_i,temp_m4_16_8_r,temp_m4_16_8_i,temp_m4_16_16_r,temp_m4_16_16_i,`W7_real,`W7_imag,`W7_real,`W7_imag,`W14_real,`W14_imag);
butterfly butterfly256 (clk,temp_m4_8_8_r,temp_m4_8_8_i,temp_m4_8_16_r,temp_m4_8_16_i,temp_m4_16_8_r,temp_m4_16_8_i,temp_m4_16_16_r,temp_m4_16_16_i,temp_b4_8_8_r,temp_b4_8_8_i,temp_b4_8_16_r,temp_b4_8_16_i,temp_b4_16_8_r,temp_b4_16_8_i,temp_b4_16_16_r,temp_b4_16_16_i);

/******************in out assgin*******************/

assign in_1_1_r = in_r;
assign in_1_1_i = in_i;
assign in_1_2_r = in_r;
assign in_1_2_i = in_i;
assign in_1_3_r = in_r;
assign in_1_3_i = in_i;
assign in_1_4_r = in_r;
assign in_1_4_i = in_i;
assign in_1_5_r = in_r;
assign in_1_5_i = in_i;
assign in_1_6_r = in_r;
assign in_1_6_i = in_i;
assign in_1_7_r = in_r;
assign in_1_7_i = in_i;
assign in_1_8_r = in_r;
assign in_1_8_i = in_i;
assign in_1_9_r = in_r;
assign in_1_9_i = in_i;
assign in_1_10_r = in_r;
assign in_1_10_i = in_i;
assign in_1_11_r = in_r;
assign in_1_11_i = in_i;
assign in_1_12_r = in_r;
assign in_1_12_i = in_i;
assign in_1_13_r = in_r;
assign in_1_13_i = in_i;
assign in_1_14_r = in_r;
assign in_1_14_i = in_i;
assign in_1_15_r = in_r;
assign in_1_15_i = in_i;
assign in_1_16_r = in_r;
assign in_1_16_i = in_i;
assign in_2_1_r = in_r;
assign in_2_1_i = in_i;
assign in_2_2_r = in_r;
assign in_2_2_i = in_i;
assign in_2_3_r = in_r;
assign in_2_3_i = in_i;
assign in_2_4_r = in_r;
assign in_2_4_i = in_i;
assign in_2_5_r = in_r;
assign in_2_5_i = in_i;
assign in_2_6_r = in_r;
assign in_2_6_i = in_i;
assign in_2_7_r = in_r;
assign in_2_7_i = in_i;
assign in_2_8_r = in_r;
assign in_2_8_i = in_i;
assign in_2_9_r = in_r;
assign in_2_9_i = in_i;
assign in_2_10_r = in_r;
assign in_2_10_i = in_i;
assign in_2_11_r = in_r;
assign in_2_11_i = in_i;
assign in_2_12_r = in_r;
assign in_2_12_i = in_i;
assign in_2_13_r = in_r;
assign in_2_13_i = in_i;
assign in_2_14_r = in_r;
assign in_2_14_i = in_i;
assign in_2_15_r = in_r;
assign in_2_15_i = in_i;
assign in_2_16_r = in_r;
assign in_2_16_i = in_i;
assign in_3_1_r = in_r;
assign in_3_1_i = in_i;
assign in_3_2_r = in_r;
assign in_3_2_i = in_i;
assign in_3_3_r = in_r;
assign in_3_3_i = in_i;
assign in_3_4_r = in_r;
assign in_3_4_i = in_i;
assign in_3_5_r = in_r;
assign in_3_5_i = in_i;
assign in_3_6_r = in_r;
assign in_3_6_i = in_i;
assign in_3_7_r = in_r;
assign in_3_7_i = in_i;
assign in_3_8_r = in_r;
assign in_3_8_i = in_i;
assign in_3_9_r = in_r;
assign in_3_9_i = in_i;
assign in_3_10_r = in_r;
assign in_3_10_i = in_i;
assign in_3_11_r = in_r;
assign in_3_11_i = in_i;
assign in_3_12_r = in_r;
assign in_3_12_i = in_i;
assign in_3_13_r = in_r;
assign in_3_13_i = in_i;
assign in_3_14_r = in_r;
assign in_3_14_i = in_i;
assign in_3_15_r = in_r;
assign in_3_15_i = in_i;
assign in_3_16_r = in_r;
assign in_3_16_i = in_i;
assign in_4_1_r = in_r;
assign in_4_1_i = in_i;
assign in_4_2_r = in_r;
assign in_4_2_i = in_i;
assign in_4_3_r = in_r;
assign in_4_3_i = in_i;
assign in_4_4_r = in_r;
assign in_4_4_i = in_i;
assign in_4_5_r = in_r;
assign in_4_5_i = in_i;
assign in_4_6_r = in_r;
assign in_4_6_i = in_i;
assign in_4_7_r = in_r;
assign in_4_7_i = in_i;
assign in_4_8_r = in_r;
assign in_4_8_i = in_i;
assign in_4_9_r = in_r;
assign in_4_9_i = in_i;
assign in_4_10_r = in_r;
assign in_4_10_i = in_i;
assign in_4_11_r = in_r;
assign in_4_11_i = in_i;
assign in_4_12_r = in_r;
assign in_4_12_i = in_i;
assign in_4_13_r = in_r;
assign in_4_13_i = in_i;
assign in_4_14_r = in_r;
assign in_4_14_i = in_i;
assign in_4_15_r = in_r;
assign in_4_15_i = in_i;
assign in_4_16_r = in_r;
assign in_4_16_i = in_i;
assign in_5_1_r = in_r;
assign in_5_1_i = in_i;
assign in_5_2_r = in_r;
assign in_5_2_i = in_i;
assign in_5_3_r = in_r;
assign in_5_3_i = in_i;
assign in_5_4_r = in_r;
assign in_5_4_i = in_i;
assign in_5_5_r = in_r;
assign in_5_5_i = in_i;
assign in_5_6_r = in_r;
assign in_5_6_i = in_i;
assign in_5_7_r = in_r;
assign in_5_7_i = in_i;
assign in_5_8_r = in_r;
assign in_5_8_i = in_i;
assign in_5_9_r = in_r;
assign in_5_9_i = in_i;
assign in_5_10_r = in_r;
assign in_5_10_i = in_i;
assign in_5_11_r = in_r;
assign in_5_11_i = in_i;
assign in_5_12_r = in_r;
assign in_5_12_i = in_i;
assign in_5_13_r = in_r;
assign in_5_13_i = in_i;
assign in_5_14_r = in_r;
assign in_5_14_i = in_i;
assign in_5_15_r = in_r;
assign in_5_15_i = in_i;
assign in_5_16_r = in_r;
assign in_5_16_i = in_i;
assign in_6_1_r = in_r;
assign in_6_1_i = in_i;
assign in_6_2_r = in_r;
assign in_6_2_i = in_i;
assign in_6_3_r = in_r;
assign in_6_3_i = in_i;
assign in_6_4_r = in_r;
assign in_6_4_i = in_i;
assign in_6_5_r = in_r;
assign in_6_5_i = in_i;
assign in_6_6_r = in_r;
assign in_6_6_i = in_i;
assign in_6_7_r = in_r;
assign in_6_7_i = in_i;
assign in_6_8_r = in_r;
assign in_6_8_i = in_i;
assign in_6_9_r = in_r;
assign in_6_9_i = in_i;
assign in_6_10_r = in_r;
assign in_6_10_i = in_i;
assign in_6_11_r = in_r;
assign in_6_11_i = in_i;
assign in_6_12_r = in_r;
assign in_6_12_i = in_i;
assign in_6_13_r = in_r;
assign in_6_13_i = in_i;
assign in_6_14_r = in_r;
assign in_6_14_i = in_i;
assign in_6_15_r = in_r;
assign in_6_15_i = in_i;
assign in_6_16_r = in_r;
assign in_6_16_i = in_i;
assign in_7_1_r = in_r;
assign in_7_1_i = in_i;
assign in_7_2_r = in_r;
assign in_7_2_i = in_i;
assign in_7_3_r = in_r;
assign in_7_3_i = in_i;
assign in_7_4_r = in_r;
assign in_7_4_i = in_i;
assign in_7_5_r = in_r;
assign in_7_5_i = in_i;
assign in_7_6_r = in_r;
assign in_7_6_i = in_i;
assign in_7_7_r = in_r;
assign in_7_7_i = in_i;
assign in_7_8_r = in_r;
assign in_7_8_i = in_i;
assign in_7_9_r = in_r;
assign in_7_9_i = in_i;
assign in_7_10_r = in_r;
assign in_7_10_i = in_i;
assign in_7_11_r = in_r;
assign in_7_11_i = in_i;
assign in_7_12_r = in_r;
assign in_7_12_i = in_i;
assign in_7_13_r = in_r;
assign in_7_13_i = in_i;
assign in_7_14_r = in_r;
assign in_7_14_i = in_i;
assign in_7_15_r = in_r;
assign in_7_15_i = in_i;
assign in_7_16_r = in_r;
assign in_7_16_i = in_i;
assign in_8_1_r = in_r;
assign in_8_1_i = in_i;
assign in_8_2_r = in_r;
assign in_8_2_i = in_i;
assign in_8_3_r = in_r;
assign in_8_3_i = in_i;
assign in_8_4_r = in_r;
assign in_8_4_i = in_i;
assign in_8_5_r = in_r;
assign in_8_5_i = in_i;
assign in_8_6_r = in_r;
assign in_8_6_i = in_i;
assign in_8_7_r = in_r;
assign in_8_7_i = in_i;
assign in_8_8_r = in_r;
assign in_8_8_i = in_i;
assign in_8_9_r = in_r;
assign in_8_9_i = in_i;
assign in_8_10_r = in_r;
assign in_8_10_i = in_i;
assign in_8_11_r = in_r;
assign in_8_11_i = in_i;
assign in_8_12_r = in_r;
assign in_8_12_i = in_i;
assign in_8_13_r = in_r;
assign in_8_13_i = in_i;
assign in_8_14_r = in_r;
assign in_8_14_i = in_i;
assign in_8_15_r = in_r;
assign in_8_15_i = in_i;
assign in_8_16_r = in_r;
assign in_8_16_i = in_i;
assign in_9_1_r = in_r;
assign in_9_1_i = in_i;
assign in_9_2_r = in_r;
assign in_9_2_i = in_i;
assign in_9_3_r = in_r;
assign in_9_3_i = in_i;
assign in_9_4_r = in_r;
assign in_9_4_i = in_i;
assign in_9_5_r = in_r;
assign in_9_5_i = in_i;
assign in_9_6_r = in_r;
assign in_9_6_i = in_i;
assign in_9_7_r = in_r;
assign in_9_7_i = in_i;
assign in_9_8_r = in_r;
assign in_9_8_i = in_i;
assign in_9_9_r = in_r;
assign in_9_9_i = in_i;
assign in_9_10_r = in_r;
assign in_9_10_i = in_i;
assign in_9_11_r = in_r;
assign in_9_11_i = in_i;
assign in_9_12_r = in_r;
assign in_9_12_i = in_i;
assign in_9_13_r = in_r;
assign in_9_13_i = in_i;
assign in_9_14_r = in_r;
assign in_9_14_i = in_i;
assign in_9_15_r = in_r;
assign in_9_15_i = in_i;
assign in_9_16_r = in_r;
assign in_9_16_i = in_i;
assign in_10_1_r = in_r;
assign in_10_1_i = in_i;
assign in_10_2_r = in_r;
assign in_10_2_i = in_i;
assign in_10_3_r = in_r;
assign in_10_3_i = in_i;
assign in_10_4_r = in_r;
assign in_10_4_i = in_i;
assign in_10_5_r = in_r;
assign in_10_5_i = in_i;
assign in_10_6_r = in_r;
assign in_10_6_i = in_i;
assign in_10_7_r = in_r;
assign in_10_7_i = in_i;
assign in_10_8_r = in_r;
assign in_10_8_i = in_i;
assign in_10_9_r = in_r;
assign in_10_9_i = in_i;
assign in_10_10_r = in_r;
assign in_10_10_i = in_i;
assign in_10_11_r = in_r;
assign in_10_11_i = in_i;
assign in_10_12_r = in_r;
assign in_10_12_i = in_i;
assign in_10_13_r = in_r;
assign in_10_13_i = in_i;
assign in_10_14_r = in_r;
assign in_10_14_i = in_i;
assign in_10_15_r = in_r;
assign in_10_15_i = in_i;
assign in_10_16_r = in_r;
assign in_10_16_i = in_i;
assign in_11_1_r = in_r;
assign in_11_1_i = in_i;
assign in_11_2_r = in_r;
assign in_11_2_i = in_i;
assign in_11_3_r = in_r;
assign in_11_3_i = in_i;
assign in_11_4_r = in_r;
assign in_11_4_i = in_i;
assign in_11_5_r = in_r;
assign in_11_5_i = in_i;
assign in_11_6_r = in_r;
assign in_11_6_i = in_i;
assign in_11_7_r = in_r;
assign in_11_7_i = in_i;
assign in_11_8_r = in_r;
assign in_11_8_i = in_i;
assign in_11_9_r = in_r;
assign in_11_9_i = in_i;
assign in_11_10_r = in_r;
assign in_11_10_i = in_i;
assign in_11_11_r = in_r;
assign in_11_11_i = in_i;
assign in_11_12_r = in_r;
assign in_11_12_i = in_i;
assign in_11_13_r = in_r;
assign in_11_13_i = in_i;
assign in_11_14_r = in_r;
assign in_11_14_i = in_i;
assign in_11_15_r = in_r;
assign in_11_15_i = in_i;
assign in_11_16_r = in_r;
assign in_11_16_i = in_i;
assign in_12_1_r = in_r;
assign in_12_1_i = in_i;
assign in_12_2_r = in_r;
assign in_12_2_i = in_i;
assign in_12_3_r = in_r;
assign in_12_3_i = in_i;
assign in_12_4_r = in_r;
assign in_12_4_i = in_i;
assign in_12_5_r = in_r;
assign in_12_5_i = in_i;
assign in_12_6_r = in_r;
assign in_12_6_i = in_i;
assign in_12_7_r = in_r;
assign in_12_7_i = in_i;
assign in_12_8_r = in_r;
assign in_12_8_i = in_i;
assign in_12_9_r = in_r;
assign in_12_9_i = in_i;
assign in_12_10_r = in_r;
assign in_12_10_i = in_i;
assign in_12_11_r = in_r;
assign in_12_11_i = in_i;
assign in_12_12_r = in_r;
assign in_12_12_i = in_i;
assign in_12_13_r = in_r;
assign in_12_13_i = in_i;
assign in_12_14_r = in_r;
assign in_12_14_i = in_i;
assign in_12_15_r = in_r;
assign in_12_15_i = in_i;
assign in_12_16_r = in_r;
assign in_12_16_i = in_i;
assign in_13_1_r = in_r;
assign in_13_1_i = in_i;
assign in_13_2_r = in_r;
assign in_13_2_i = in_i;
assign in_13_3_r = in_r;
assign in_13_3_i = in_i;
assign in_13_4_r = in_r;
assign in_13_4_i = in_i;
assign in_13_5_r = in_r;
assign in_13_5_i = in_i;
assign in_13_6_r = in_r;
assign in_13_6_i = in_i;
assign in_13_7_r = in_r;
assign in_13_7_i = in_i;
assign in_13_8_r = in_r;
assign in_13_8_i = in_i;
assign in_13_9_r = in_r;
assign in_13_9_i = in_i;
assign in_13_10_r = in_r;
assign in_13_10_i = in_i;
assign in_13_11_r = in_r;
assign in_13_11_i = in_i;
assign in_13_12_r = in_r;
assign in_13_12_i = in_i;
assign in_13_13_r = in_r;
assign in_13_13_i = in_i;
assign in_13_14_r = in_r;
assign in_13_14_i = in_i;
assign in_13_15_r = in_r;
assign in_13_15_i = in_i;
assign in_13_16_r = in_r;
assign in_13_16_i = in_i;
assign in_14_1_r = in_r;
assign in_14_1_i = in_i;
assign in_14_2_r = in_r;
assign in_14_2_i = in_i;
assign in_14_3_r = in_r;
assign in_14_3_i = in_i;
assign in_14_4_r = in_r;
assign in_14_4_i = in_i;
assign in_14_5_r = in_r;
assign in_14_5_i = in_i;
assign in_14_6_r = in_r;
assign in_14_6_i = in_i;
assign in_14_7_r = in_r;
assign in_14_7_i = in_i;
assign in_14_8_r = in_r;
assign in_14_8_i = in_i;
assign in_14_9_r = in_r;
assign in_14_9_i = in_i;
assign in_14_10_r = in_r;
assign in_14_10_i = in_i;
assign in_14_11_r = in_r;
assign in_14_11_i = in_i;
assign in_14_12_r = in_r;
assign in_14_12_i = in_i;
assign in_14_13_r = in_r;
assign in_14_13_i = in_i;
assign in_14_14_r = in_r;
assign in_14_14_i = in_i;
assign in_14_15_r = in_r;
assign in_14_15_i = in_i;
assign in_14_16_r = in_r;
assign in_14_16_i = in_i;
assign in_15_1_r = in_r;
assign in_15_1_i = in_i;
assign in_15_2_r = in_r;
assign in_15_2_i = in_i;
assign in_15_3_r = in_r;
assign in_15_3_i = in_i;
assign in_15_4_r = in_r;
assign in_15_4_i = in_i;
assign in_15_5_r = in_r;
assign in_15_5_i = in_i;
assign in_15_6_r = in_r;
assign in_15_6_i = in_i;
assign in_15_7_r = in_r;
assign in_15_7_i = in_i;
assign in_15_8_r = in_r;
assign in_15_8_i = in_i;
assign in_15_9_r = in_r;
assign in_15_9_i = in_i;
assign in_15_10_r = in_r;
assign in_15_10_i = in_i;
assign in_15_11_r = in_r;
assign in_15_11_i = in_i;
assign in_15_12_r = in_r;
assign in_15_12_i = in_i;
assign in_15_13_r = in_r;
assign in_15_13_i = in_i;
assign in_15_14_r = in_r;
assign in_15_14_i = in_i;
assign in_15_15_r = in_r;
assign in_15_15_i = in_i;
assign in_15_16_r = in_r;
assign in_15_16_i = in_i;
assign in_16_1_r = in_r;
assign in_16_1_i = in_i;
assign in_16_2_r = in_r;
assign in_16_2_i = in_i;
assign in_16_3_r = in_r;
assign in_16_3_i = in_i;
assign in_16_4_r = in_r;
assign in_16_4_i = in_i;
assign in_16_5_r = in_r;
assign in_16_5_i = in_i;
assign in_16_6_r = in_r;
assign in_16_6_i = in_i;
assign in_16_7_r = in_r;
assign in_16_7_i = in_i;
assign in_16_8_r = in_r;
assign in_16_8_i = in_i;
assign in_16_9_r = in_r;
assign in_16_9_i = in_i;
assign in_16_10_r = in_r;
assign in_16_10_i = in_i;
assign in_16_11_r = in_r;
assign in_16_11_i = in_i;
assign in_16_12_r = in_r;
assign in_16_12_i = in_i;
assign in_16_13_r = in_r;
assign in_16_13_i = in_i;
assign in_16_14_r = in_r;
assign in_16_14_i = in_i;
assign in_16_15_r = in_r;
assign in_16_15_i = in_i;
assign in_16_16_r = in_r;
assign in_16_16_i = in_i;

assign out_1_1_r = temp_b4_1_1_r;
assign out_1_1_i = temp_b4_1_1_i;
assign out_1_2_r = temp_b4_1_2_r;
assign out_1_2_i = temp_b4_1_2_i;
assign out_1_3_r = temp_b4_1_3_r;
assign out_1_3_i = temp_b4_1_3_i;
assign out_1_4_r = temp_b4_1_4_r;
assign out_1_4_i = temp_b4_1_4_i;
assign out_1_5_r = temp_b4_1_5_r;
assign out_1_5_i = temp_b4_1_5_i;
assign out_1_6_r = temp_b4_1_6_r;
assign out_1_6_i = temp_b4_1_6_i;
assign out_1_7_r = temp_b4_1_7_r;
assign out_1_7_i = temp_b4_1_7_i;
assign out_1_8_r = temp_b4_1_8_r;
assign out_1_8_i = temp_b4_1_8_i;
assign out_1_9_r = temp_b4_1_9_r;
assign out_1_9_i = temp_b4_1_9_i;
assign out_1_10_r = temp_b4_1_10_r;
assign out_1_10_i = temp_b4_1_10_i;
assign out_1_11_r = temp_b4_1_11_r;
assign out_1_11_i = temp_b4_1_11_i;
assign out_1_12_r = temp_b4_1_12_r;
assign out_1_12_i = temp_b4_1_12_i;
assign out_1_13_r = temp_b4_1_13_r;
assign out_1_13_i = temp_b4_1_13_i;
assign out_1_14_r = temp_b4_1_14_r;
assign out_1_14_i = temp_b4_1_14_i;
assign out_1_15_r = temp_b4_1_15_r;
assign out_1_15_i = temp_b4_1_15_i;
assign out_1_16_r = temp_b4_1_16_r;
assign out_1_16_i = temp_b4_1_16_i;
assign out_2_1_r = temp_b4_2_1_r;
assign out_2_1_i = temp_b4_2_1_i;
assign out_2_2_r = temp_b4_2_2_r;
assign out_2_2_i = temp_b4_2_2_i;
assign out_2_3_r = temp_b4_2_3_r;
assign out_2_3_i = temp_b4_2_3_i;
assign out_2_4_r = temp_b4_2_4_r;
assign out_2_4_i = temp_b4_2_4_i;
assign out_2_5_r = temp_b4_2_5_r;
assign out_2_5_i = temp_b4_2_5_i;
assign out_2_6_r = temp_b4_2_6_r;
assign out_2_6_i = temp_b4_2_6_i;
assign out_2_7_r = temp_b4_2_7_r;
assign out_2_7_i = temp_b4_2_7_i;
assign out_2_8_r = temp_b4_2_8_r;
assign out_2_8_i = temp_b4_2_8_i;
assign out_2_9_r = temp_b4_2_9_r;
assign out_2_9_i = temp_b4_2_9_i;
assign out_2_10_r = temp_b4_2_10_r;
assign out_2_10_i = temp_b4_2_10_i;
assign out_2_11_r = temp_b4_2_11_r;
assign out_2_11_i = temp_b4_2_11_i;
assign out_2_12_r = temp_b4_2_12_r;
assign out_2_12_i = temp_b4_2_12_i;
assign out_2_13_r = temp_b4_2_13_r;
assign out_2_13_i = temp_b4_2_13_i;
assign out_2_14_r = temp_b4_2_14_r;
assign out_2_14_i = temp_b4_2_14_i;
assign out_2_15_r = temp_b4_2_15_r;
assign out_2_15_i = temp_b4_2_15_i;
assign out_2_16_r = temp_b4_2_16_r;
assign out_2_16_i = temp_b4_2_16_i;
assign out_3_1_r = temp_b4_3_1_r;
assign out_3_1_i = temp_b4_3_1_i;
assign out_3_2_r = temp_b4_3_2_r;
assign out_3_2_i = temp_b4_3_2_i;
assign out_3_3_r = temp_b4_3_3_r;
assign out_3_3_i = temp_b4_3_3_i;
assign out_3_4_r = temp_b4_3_4_r;
assign out_3_4_i = temp_b4_3_4_i;
assign out_3_5_r = temp_b4_3_5_r;
assign out_3_5_i = temp_b4_3_5_i;
assign out_3_6_r = temp_b4_3_6_r;
assign out_3_6_i = temp_b4_3_6_i;
assign out_3_7_r = temp_b4_3_7_r;
assign out_3_7_i = temp_b4_3_7_i;
assign out_3_8_r = temp_b4_3_8_r;
assign out_3_8_i = temp_b4_3_8_i;
assign out_3_9_r = temp_b4_3_9_r;
assign out_3_9_i = temp_b4_3_9_i;
assign out_3_10_r = temp_b4_3_10_r;
assign out_3_10_i = temp_b4_3_10_i;
assign out_3_11_r = temp_b4_3_11_r;
assign out_3_11_i = temp_b4_3_11_i;
assign out_3_12_r = temp_b4_3_12_r;
assign out_3_12_i = temp_b4_3_12_i;
assign out_3_13_r = temp_b4_3_13_r;
assign out_3_13_i = temp_b4_3_13_i;
assign out_3_14_r = temp_b4_3_14_r;
assign out_3_14_i = temp_b4_3_14_i;
assign out_3_15_r = temp_b4_3_15_r;
assign out_3_15_i = temp_b4_3_15_i;
assign out_3_16_r = temp_b4_3_16_r;
assign out_3_16_i = temp_b4_3_16_i;
assign out_4_1_r = temp_b4_4_1_r;
assign out_4_1_i = temp_b4_4_1_i;
assign out_4_2_r = temp_b4_4_2_r;
assign out_4_2_i = temp_b4_4_2_i;
assign out_4_3_r = temp_b4_4_3_r;
assign out_4_3_i = temp_b4_4_3_i;
assign out_4_4_r = temp_b4_4_4_r;
assign out_4_4_i = temp_b4_4_4_i;
assign out_4_5_r = temp_b4_4_5_r;
assign out_4_5_i = temp_b4_4_5_i;
assign out_4_6_r = temp_b4_4_6_r;
assign out_4_6_i = temp_b4_4_6_i;
assign out_4_7_r = temp_b4_4_7_r;
assign out_4_7_i = temp_b4_4_7_i;
assign out_4_8_r = temp_b4_4_8_r;
assign out_4_8_i = temp_b4_4_8_i;
assign out_4_9_r = temp_b4_4_9_r;
assign out_4_9_i = temp_b4_4_9_i;
assign out_4_10_r = temp_b4_4_10_r;
assign out_4_10_i = temp_b4_4_10_i;
assign out_4_11_r = temp_b4_4_11_r;
assign out_4_11_i = temp_b4_4_11_i;
assign out_4_12_r = temp_b4_4_12_r;
assign out_4_12_i = temp_b4_4_12_i;
assign out_4_13_r = temp_b4_4_13_r;
assign out_4_13_i = temp_b4_4_13_i;
assign out_4_14_r = temp_b4_4_14_r;
assign out_4_14_i = temp_b4_4_14_i;
assign out_4_15_r = temp_b4_4_15_r;
assign out_4_15_i = temp_b4_4_15_i;
assign out_4_16_r = temp_b4_4_16_r;
assign out_4_16_i = temp_b4_4_16_i;
assign out_5_1_r = temp_b4_5_1_r;
assign out_5_1_i = temp_b4_5_1_i;
assign out_5_2_r = temp_b4_5_2_r;
assign out_5_2_i = temp_b4_5_2_i;
assign out_5_3_r = temp_b4_5_3_r;
assign out_5_3_i = temp_b4_5_3_i;
assign out_5_4_r = temp_b4_5_4_r;
assign out_5_4_i = temp_b4_5_4_i;
assign out_5_5_r = temp_b4_5_5_r;
assign out_5_5_i = temp_b4_5_5_i;
assign out_5_6_r = temp_b4_5_6_r;
assign out_5_6_i = temp_b4_5_6_i;
assign out_5_7_r = temp_b4_5_7_r;
assign out_5_7_i = temp_b4_5_7_i;
assign out_5_8_r = temp_b4_5_8_r;
assign out_5_8_i = temp_b4_5_8_i;
assign out_5_9_r = temp_b4_5_9_r;
assign out_5_9_i = temp_b4_5_9_i;
assign out_5_10_r = temp_b4_5_10_r;
assign out_5_10_i = temp_b4_5_10_i;
assign out_5_11_r = temp_b4_5_11_r;
assign out_5_11_i = temp_b4_5_11_i;
assign out_5_12_r = temp_b4_5_12_r;
assign out_5_12_i = temp_b4_5_12_i;
assign out_5_13_r = temp_b4_5_13_r;
assign out_5_13_i = temp_b4_5_13_i;
assign out_5_14_r = temp_b4_5_14_r;
assign out_5_14_i = temp_b4_5_14_i;
assign out_5_15_r = temp_b4_5_15_r;
assign out_5_15_i = temp_b4_5_15_i;
assign out_5_16_r = temp_b4_5_16_r;
assign out_5_16_i = temp_b4_5_16_i;
assign out_6_1_r = temp_b4_6_1_r;
assign out_6_1_i = temp_b4_6_1_i;
assign out_6_2_r = temp_b4_6_2_r;
assign out_6_2_i = temp_b4_6_2_i;
assign out_6_3_r = temp_b4_6_3_r;
assign out_6_3_i = temp_b4_6_3_i;
assign out_6_4_r = temp_b4_6_4_r;
assign out_6_4_i = temp_b4_6_4_i;
assign out_6_5_r = temp_b4_6_5_r;
assign out_6_5_i = temp_b4_6_5_i;
assign out_6_6_r = temp_b4_6_6_r;
assign out_6_6_i = temp_b4_6_6_i;
assign out_6_7_r = temp_b4_6_7_r;
assign out_6_7_i = temp_b4_6_7_i;
assign out_6_8_r = temp_b4_6_8_r;
assign out_6_8_i = temp_b4_6_8_i;
assign out_6_9_r = temp_b4_6_9_r;
assign out_6_9_i = temp_b4_6_9_i;
assign out_6_10_r = temp_b4_6_10_r;
assign out_6_10_i = temp_b4_6_10_i;
assign out_6_11_r = temp_b4_6_11_r;
assign out_6_11_i = temp_b4_6_11_i;
assign out_6_12_r = temp_b4_6_12_r;
assign out_6_12_i = temp_b4_6_12_i;
assign out_6_13_r = temp_b4_6_13_r;
assign out_6_13_i = temp_b4_6_13_i;
assign out_6_14_r = temp_b4_6_14_r;
assign out_6_14_i = temp_b4_6_14_i;
assign out_6_15_r = temp_b4_6_15_r;
assign out_6_15_i = temp_b4_6_15_i;
assign out_6_16_r = temp_b4_6_16_r;
assign out_6_16_i = temp_b4_6_16_i;
assign out_7_1_r = temp_b4_7_1_r;
assign out_7_1_i = temp_b4_7_1_i;
assign out_7_2_r = temp_b4_7_2_r;
assign out_7_2_i = temp_b4_7_2_i;
assign out_7_3_r = temp_b4_7_3_r;
assign out_7_3_i = temp_b4_7_3_i;
assign out_7_4_r = temp_b4_7_4_r;
assign out_7_4_i = temp_b4_7_4_i;
assign out_7_5_r = temp_b4_7_5_r;
assign out_7_5_i = temp_b4_7_5_i;
assign out_7_6_r = temp_b4_7_6_r;
assign out_7_6_i = temp_b4_7_6_i;
assign out_7_7_r = temp_b4_7_7_r;
assign out_7_7_i = temp_b4_7_7_i;
assign out_7_8_r = temp_b4_7_8_r;
assign out_7_8_i = temp_b4_7_8_i;
assign out_7_9_r = temp_b4_7_9_r;
assign out_7_9_i = temp_b4_7_9_i;
assign out_7_10_r = temp_b4_7_10_r;
assign out_7_10_i = temp_b4_7_10_i;
assign out_7_11_r = temp_b4_7_11_r;
assign out_7_11_i = temp_b4_7_11_i;
assign out_7_12_r = temp_b4_7_12_r;
assign out_7_12_i = temp_b4_7_12_i;
assign out_7_13_r = temp_b4_7_13_r;
assign out_7_13_i = temp_b4_7_13_i;
assign out_7_14_r = temp_b4_7_14_r;
assign out_7_14_i = temp_b4_7_14_i;
assign out_7_15_r = temp_b4_7_15_r;
assign out_7_15_i = temp_b4_7_15_i;
assign out_7_16_r = temp_b4_7_16_r;
assign out_7_16_i = temp_b4_7_16_i;
assign out_8_1_r = temp_b4_8_1_r;
assign out_8_1_i = temp_b4_8_1_i;
assign out_8_2_r = temp_b4_8_2_r;
assign out_8_2_i = temp_b4_8_2_i;
assign out_8_3_r = temp_b4_8_3_r;
assign out_8_3_i = temp_b4_8_3_i;
assign out_8_4_r = temp_b4_8_4_r;
assign out_8_4_i = temp_b4_8_4_i;
assign out_8_5_r = temp_b4_8_5_r;
assign out_8_5_i = temp_b4_8_5_i;
assign out_8_6_r = temp_b4_8_6_r;
assign out_8_6_i = temp_b4_8_6_i;
assign out_8_7_r = temp_b4_8_7_r;
assign out_8_7_i = temp_b4_8_7_i;
assign out_8_8_r = temp_b4_8_8_r;
assign out_8_8_i = temp_b4_8_8_i;
assign out_8_9_r = temp_b4_8_9_r;
assign out_8_9_i = temp_b4_8_9_i;
assign out_8_10_r = temp_b4_8_10_r;
assign out_8_10_i = temp_b4_8_10_i;
assign out_8_11_r = temp_b4_8_11_r;
assign out_8_11_i = temp_b4_8_11_i;
assign out_8_12_r = temp_b4_8_12_r;
assign out_8_12_i = temp_b4_8_12_i;
assign out_8_13_r = temp_b4_8_13_r;
assign out_8_13_i = temp_b4_8_13_i;
assign out_8_14_r = temp_b4_8_14_r;
assign out_8_14_i = temp_b4_8_14_i;
assign out_8_15_r = temp_b4_8_15_r;
assign out_8_15_i = temp_b4_8_15_i;
assign out_8_16_r = temp_b4_8_16_r;
assign out_8_16_i = temp_b4_8_16_i;
assign out_9_1_r = temp_b4_9_1_r;
assign out_9_1_i = temp_b4_9_1_i;
assign out_9_2_r = temp_b4_9_2_r;
assign out_9_2_i = temp_b4_9_2_i;
assign out_9_3_r = temp_b4_9_3_r;
assign out_9_3_i = temp_b4_9_3_i;
assign out_9_4_r = temp_b4_9_4_r;
assign out_9_4_i = temp_b4_9_4_i;
assign out_9_5_r = temp_b4_9_5_r;
assign out_9_5_i = temp_b4_9_5_i;
assign out_9_6_r = temp_b4_9_6_r;
assign out_9_6_i = temp_b4_9_6_i;
assign out_9_7_r = temp_b4_9_7_r;
assign out_9_7_i = temp_b4_9_7_i;
assign out_9_8_r = temp_b4_9_8_r;
assign out_9_8_i = temp_b4_9_8_i;
assign out_9_9_r = temp_b4_9_9_r;
assign out_9_9_i = temp_b4_9_9_i;
assign out_9_10_r = temp_b4_9_10_r;
assign out_9_10_i = temp_b4_9_10_i;
assign out_9_11_r = temp_b4_9_11_r;
assign out_9_11_i = temp_b4_9_11_i;
assign out_9_12_r = temp_b4_9_12_r;
assign out_9_12_i = temp_b4_9_12_i;
assign out_9_13_r = temp_b4_9_13_r;
assign out_9_13_i = temp_b4_9_13_i;
assign out_9_14_r = temp_b4_9_14_r;
assign out_9_14_i = temp_b4_9_14_i;
assign out_9_15_r = temp_b4_9_15_r;
assign out_9_15_i = temp_b4_9_15_i;
assign out_9_16_r = temp_b4_9_16_r;
assign out_9_16_i = temp_b4_9_16_i;
assign out_10_1_r = temp_b4_10_1_r;
assign out_10_1_i = temp_b4_10_1_i;
assign out_10_2_r = temp_b4_10_2_r;
assign out_10_2_i = temp_b4_10_2_i;
assign out_10_3_r = temp_b4_10_3_r;
assign out_10_3_i = temp_b4_10_3_i;
assign out_10_4_r = temp_b4_10_4_r;
assign out_10_4_i = temp_b4_10_4_i;
assign out_10_5_r = temp_b4_10_5_r;
assign out_10_5_i = temp_b4_10_5_i;
assign out_10_6_r = temp_b4_10_6_r;
assign out_10_6_i = temp_b4_10_6_i;
assign out_10_7_r = temp_b4_10_7_r;
assign out_10_7_i = temp_b4_10_7_i;
assign out_10_8_r = temp_b4_10_8_r;
assign out_10_8_i = temp_b4_10_8_i;
assign out_10_9_r = temp_b4_10_9_r;
assign out_10_9_i = temp_b4_10_9_i;
assign out_10_10_r = temp_b4_10_10_r;
assign out_10_10_i = temp_b4_10_10_i;
assign out_10_11_r = temp_b4_10_11_r;
assign out_10_11_i = temp_b4_10_11_i;
assign out_10_12_r = temp_b4_10_12_r;
assign out_10_12_i = temp_b4_10_12_i;
assign out_10_13_r = temp_b4_10_13_r;
assign out_10_13_i = temp_b4_10_13_i;
assign out_10_14_r = temp_b4_10_14_r;
assign out_10_14_i = temp_b4_10_14_i;
assign out_10_15_r = temp_b4_10_15_r;
assign out_10_15_i = temp_b4_10_15_i;
assign out_10_16_r = temp_b4_10_16_r;
assign out_10_16_i = temp_b4_10_16_i;
assign out_11_1_r = temp_b4_11_1_r;
assign out_11_1_i = temp_b4_11_1_i;
assign out_11_2_r = temp_b4_11_2_r;
assign out_11_2_i = temp_b4_11_2_i;
assign out_11_3_r = temp_b4_11_3_r;
assign out_11_3_i = temp_b4_11_3_i;
assign out_11_4_r = temp_b4_11_4_r;
assign out_11_4_i = temp_b4_11_4_i;
assign out_11_5_r = temp_b4_11_5_r;
assign out_11_5_i = temp_b4_11_5_i;
assign out_11_6_r = temp_b4_11_6_r;
assign out_11_6_i = temp_b4_11_6_i;
assign out_11_7_r = temp_b4_11_7_r;
assign out_11_7_i = temp_b4_11_7_i;
assign out_11_8_r = temp_b4_11_8_r;
assign out_11_8_i = temp_b4_11_8_i;
assign out_11_9_r = temp_b4_11_9_r;
assign out_11_9_i = temp_b4_11_9_i;
assign out_11_10_r = temp_b4_11_10_r;
assign out_11_10_i = temp_b4_11_10_i;
assign out_11_11_r = temp_b4_11_11_r;
assign out_11_11_i = temp_b4_11_11_i;
assign out_11_12_r = temp_b4_11_12_r;
assign out_11_12_i = temp_b4_11_12_i;
assign out_11_13_r = temp_b4_11_13_r;
assign out_11_13_i = temp_b4_11_13_i;
assign out_11_14_r = temp_b4_11_14_r;
assign out_11_14_i = temp_b4_11_14_i;
assign out_11_15_r = temp_b4_11_15_r;
assign out_11_15_i = temp_b4_11_15_i;
assign out_11_16_r = temp_b4_11_16_r;
assign out_11_16_i = temp_b4_11_16_i;
assign out_12_1_r = temp_b4_12_1_r;
assign out_12_1_i = temp_b4_12_1_i;
assign out_12_2_r = temp_b4_12_2_r;
assign out_12_2_i = temp_b4_12_2_i;
assign out_12_3_r = temp_b4_12_3_r;
assign out_12_3_i = temp_b4_12_3_i;
assign out_12_4_r = temp_b4_12_4_r;
assign out_12_4_i = temp_b4_12_4_i;
assign out_12_5_r = temp_b4_12_5_r;
assign out_12_5_i = temp_b4_12_5_i;
assign out_12_6_r = temp_b4_12_6_r;
assign out_12_6_i = temp_b4_12_6_i;
assign out_12_7_r = temp_b4_12_7_r;
assign out_12_7_i = temp_b4_12_7_i;
assign out_12_8_r = temp_b4_12_8_r;
assign out_12_8_i = temp_b4_12_8_i;
assign out_12_9_r = temp_b4_12_9_r;
assign out_12_9_i = temp_b4_12_9_i;
assign out_12_10_r = temp_b4_12_10_r;
assign out_12_10_i = temp_b4_12_10_i;
assign out_12_11_r = temp_b4_12_11_r;
assign out_12_11_i = temp_b4_12_11_i;
assign out_12_12_r = temp_b4_12_12_r;
assign out_12_12_i = temp_b4_12_12_i;
assign out_12_13_r = temp_b4_12_13_r;
assign out_12_13_i = temp_b4_12_13_i;
assign out_12_14_r = temp_b4_12_14_r;
assign out_12_14_i = temp_b4_12_14_i;
assign out_12_15_r = temp_b4_12_15_r;
assign out_12_15_i = temp_b4_12_15_i;
assign out_12_16_r = temp_b4_12_16_r;
assign out_12_16_i = temp_b4_12_16_i;
assign out_13_1_r = temp_b4_13_1_r;
assign out_13_1_i = temp_b4_13_1_i;
assign out_13_2_r = temp_b4_13_2_r;
assign out_13_2_i = temp_b4_13_2_i;
assign out_13_3_r = temp_b4_13_3_r;
assign out_13_3_i = temp_b4_13_3_i;
assign out_13_4_r = temp_b4_13_4_r;
assign out_13_4_i = temp_b4_13_4_i;
assign out_13_5_r = temp_b4_13_5_r;
assign out_13_5_i = temp_b4_13_5_i;
assign out_13_6_r = temp_b4_13_6_r;
assign out_13_6_i = temp_b4_13_6_i;
assign out_13_7_r = temp_b4_13_7_r;
assign out_13_7_i = temp_b4_13_7_i;
assign out_13_8_r = temp_b4_13_8_r;
assign out_13_8_i = temp_b4_13_8_i;
assign out_13_9_r = temp_b4_13_9_r;
assign out_13_9_i = temp_b4_13_9_i;
assign out_13_10_r = temp_b4_13_10_r;
assign out_13_10_i = temp_b4_13_10_i;
assign out_13_11_r = temp_b4_13_11_r;
assign out_13_11_i = temp_b4_13_11_i;
assign out_13_12_r = temp_b4_13_12_r;
assign out_13_12_i = temp_b4_13_12_i;
assign out_13_13_r = temp_b4_13_13_r;
assign out_13_13_i = temp_b4_13_13_i;
assign out_13_14_r = temp_b4_13_14_r;
assign out_13_14_i = temp_b4_13_14_i;
assign out_13_15_r = temp_b4_13_15_r;
assign out_13_15_i = temp_b4_13_15_i;
assign out_13_16_r = temp_b4_13_16_r;
assign out_13_16_i = temp_b4_13_16_i;
assign out_14_1_r = temp_b4_14_1_r;
assign out_14_1_i = temp_b4_14_1_i;
assign out_14_2_r = temp_b4_14_2_r;
assign out_14_2_i = temp_b4_14_2_i;
assign out_14_3_r = temp_b4_14_3_r;
assign out_14_3_i = temp_b4_14_3_i;
assign out_14_4_r = temp_b4_14_4_r;
assign out_14_4_i = temp_b4_14_4_i;
assign out_14_5_r = temp_b4_14_5_r;
assign out_14_5_i = temp_b4_14_5_i;
assign out_14_6_r = temp_b4_14_6_r;
assign out_14_6_i = temp_b4_14_6_i;
assign out_14_7_r = temp_b4_14_7_r;
assign out_14_7_i = temp_b4_14_7_i;
assign out_14_8_r = temp_b4_14_8_r;
assign out_14_8_i = temp_b4_14_8_i;
assign out_14_9_r = temp_b4_14_9_r;
assign out_14_9_i = temp_b4_14_9_i;
assign out_14_10_r = temp_b4_14_10_r;
assign out_14_10_i = temp_b4_14_10_i;
assign out_14_11_r = temp_b4_14_11_r;
assign out_14_11_i = temp_b4_14_11_i;
assign out_14_12_r = temp_b4_14_12_r;
assign out_14_12_i = temp_b4_14_12_i;
assign out_14_13_r = temp_b4_14_13_r;
assign out_14_13_i = temp_b4_14_13_i;
assign out_14_14_r = temp_b4_14_14_r;
assign out_14_14_i = temp_b4_14_14_i;
assign out_14_15_r = temp_b4_14_15_r;
assign out_14_15_i = temp_b4_14_15_i;
assign out_14_16_r = temp_b4_14_16_r;
assign out_14_16_i = temp_b4_14_16_i;
assign out_15_1_r = temp_b4_15_1_r;
assign out_15_1_i = temp_b4_15_1_i;
assign out_15_2_r = temp_b4_15_2_r;
assign out_15_2_i = temp_b4_15_2_i;
assign out_15_3_r = temp_b4_15_3_r;
assign out_15_3_i = temp_b4_15_3_i;
assign out_15_4_r = temp_b4_15_4_r;
assign out_15_4_i = temp_b4_15_4_i;
assign out_15_5_r = temp_b4_15_5_r;
assign out_15_5_i = temp_b4_15_5_i;
assign out_15_6_r = temp_b4_15_6_r;
assign out_15_6_i = temp_b4_15_6_i;
assign out_15_7_r = temp_b4_15_7_r;
assign out_15_7_i = temp_b4_15_7_i;
assign out_15_8_r = temp_b4_15_8_r;
assign out_15_8_i = temp_b4_15_8_i;
assign out_15_9_r = temp_b4_15_9_r;
assign out_15_9_i = temp_b4_15_9_i;
assign out_15_10_r = temp_b4_15_10_r;
assign out_15_10_i = temp_b4_15_10_i;
assign out_15_11_r = temp_b4_15_11_r;
assign out_15_11_i = temp_b4_15_11_i;
assign out_15_12_r = temp_b4_15_12_r;
assign out_15_12_i = temp_b4_15_12_i;
assign out_15_13_r = temp_b4_15_13_r;
assign out_15_13_i = temp_b4_15_13_i;
assign out_15_14_r = temp_b4_15_14_r;
assign out_15_14_i = temp_b4_15_14_i;
assign out_15_15_r = temp_b4_15_15_r;
assign out_15_15_i = temp_b4_15_15_i;
assign out_15_16_r = temp_b4_15_16_r;
assign out_15_16_i = temp_b4_15_16_i;
assign out_16_1_r = temp_b4_16_1_r;
assign out_16_1_i = temp_b4_16_1_i;
assign out_16_2_r = temp_b4_16_2_r;
assign out_16_2_i = temp_b4_16_2_i;
assign out_16_3_r = temp_b4_16_3_r;
assign out_16_3_i = temp_b4_16_3_i;
assign out_16_4_r = temp_b4_16_4_r;
assign out_16_4_i = temp_b4_16_4_i;
assign out_16_5_r = temp_b4_16_5_r;
assign out_16_5_i = temp_b4_16_5_i;
assign out_16_6_r = temp_b4_16_6_r;
assign out_16_6_i = temp_b4_16_6_i;
assign out_16_7_r = temp_b4_16_7_r;
assign out_16_7_i = temp_b4_16_7_i;
assign out_16_8_r = temp_b4_16_8_r;
assign out_16_8_i = temp_b4_16_8_i;
assign out_16_9_r = temp_b4_16_9_r;
assign out_16_9_i = temp_b4_16_9_i;
assign out_16_10_r = temp_b4_16_10_r;
assign out_16_10_i = temp_b4_16_10_i;
assign out_16_11_r = temp_b4_16_11_r;
assign out_16_11_i = temp_b4_16_11_i;
assign out_16_12_r = temp_b4_16_12_r;
assign out_16_12_i = temp_b4_16_12_i;
assign out_16_13_r = temp_b4_16_13_r;
assign out_16_13_i = temp_b4_16_13_i;
assign out_16_14_r = temp_b4_16_14_r;
assign out_16_14_i = temp_b4_16_14_i;
assign out_16_15_r = temp_b4_16_15_r;
assign out_16_15_i = temp_b4_16_15_i;
assign out_16_16_r = temp_b4_16_16_r;
assign out_16_16_i = temp_b4_16_16_i;

assign out_r = out_1_1_r;
assign out_i = out_1_1_i;



endmodule
