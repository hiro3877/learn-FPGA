`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/08/20 20:43:41
// Design Name: 
// Module Name: top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
/////////////////////////////////////////////////////////////////////////////////

`include "./nettype.h"
`include "./std_define.h"

module top(
input wire		clk,

input wire signed [`InBus]		in_1_1_r,
input wire signed [`InBus]		in_1_1_i,
input wire signed [`InBus]		in_1_2_r,
input wire signed [`InBus]		in_1_2_i,
input wire signed [`InBus]		in_1_3_r,
input wire signed [`InBus]		in_1_3_i,
input wire signed [`InBus]		in_1_4_r,
input wire signed [`InBus]		in_1_4_i,
input wire signed [`InBus]		in_1_5_r,
input wire signed [`InBus]		in_1_5_i,
input wire signed [`InBus]		in_1_6_r,
input wire signed [`InBus]		in_1_6_i,
input wire signed [`InBus]		in_1_7_r,
input wire signed [`InBus]		in_1_7_i,
input wire signed [`InBus]		in_1_8_r,
input wire signed [`InBus]		in_1_8_i,
input wire signed [`InBus]		in_2_1_r,
input wire signed [`InBus]		in_2_1_i,
input wire signed [`InBus]		in_2_2_r,
input wire signed [`InBus]		in_2_2_i,
input wire signed [`InBus]		in_2_3_r,
input wire signed [`InBus]		in_2_3_i,
input wire signed [`InBus]		in_2_4_r,
input wire signed [`InBus]		in_2_4_i,
input wire signed [`InBus]		in_2_5_r,
input wire signed [`InBus]		in_2_5_i,
input wire signed [`InBus]		in_2_6_r,
input wire signed [`InBus]		in_2_6_i,
input wire signed [`InBus]		in_2_7_r,
input wire signed [`InBus]		in_2_7_i,
input wire signed [`InBus]		in_2_8_r,
input wire signed [`InBus]		in_2_8_i,
input wire signed [`InBus]		in_3_1_r,
input wire signed [`InBus]		in_3_1_i,
input wire signed [`InBus]		in_3_2_r,
input wire signed [`InBus]		in_3_2_i,
input wire signed [`InBus]		in_3_3_r,
input wire signed [`InBus]		in_3_3_i,
input wire signed [`InBus]		in_3_4_r,
input wire signed [`InBus]		in_3_4_i,
input wire signed [`InBus]		in_3_5_r,
input wire signed [`InBus]		in_3_5_i,
input wire signed [`InBus]		in_3_6_r,
input wire signed [`InBus]		in_3_6_i,
input wire signed [`InBus]		in_3_7_r,
input wire signed [`InBus]		in_3_7_i,
input wire signed [`InBus]		in_3_8_r,
input wire signed [`InBus]		in_3_8_i,
input wire signed [`InBus]		in_4_1_r,
input wire signed [`InBus]		in_4_1_i,
input wire signed [`InBus]		in_4_2_r,
input wire signed [`InBus]		in_4_2_i,
input wire signed [`InBus]		in_4_3_r,
input wire signed [`InBus]		in_4_3_i,
input wire signed [`InBus]		in_4_4_r,
input wire signed [`InBus]		in_4_4_i,
input wire signed [`InBus]		in_4_5_r,
input wire signed [`InBus]		in_4_5_i,
input wire signed [`InBus]		in_4_6_r,
input wire signed [`InBus]		in_4_6_i,
input wire signed [`InBus]		in_4_7_r,
input wire signed [`InBus]		in_4_7_i,
input wire signed [`InBus]		in_4_8_r,
input wire signed [`InBus]		in_4_8_i,
input wire signed [`InBus]		in_5_1_r,
input wire signed [`InBus]		in_5_1_i,
input wire signed [`InBus]		in_5_2_r,
input wire signed [`InBus]		in_5_2_i,
input wire signed [`InBus]		in_5_3_r,
input wire signed [`InBus]		in_5_3_i,
input wire signed [`InBus]		in_5_4_r,
input wire signed [`InBus]		in_5_4_i,
input wire signed [`InBus]		in_5_5_r,
input wire signed [`InBus]		in_5_5_i,
input wire signed [`InBus]		in_5_6_r,
input wire signed [`InBus]		in_5_6_i,
input wire signed [`InBus]		in_5_7_r,
input wire signed [`InBus]		in_5_7_i,
input wire signed [`InBus]		in_5_8_r,
input wire signed [`InBus]		in_5_8_i,
input wire signed [`InBus]		in_6_1_r,
input wire signed [`InBus]		in_6_1_i,
input wire signed [`InBus]		in_6_2_r,
input wire signed [`InBus]		in_6_2_i,
input wire signed [`InBus]		in_6_3_r,
input wire signed [`InBus]		in_6_3_i,
input wire signed [`InBus]		in_6_4_r,
input wire signed [`InBus]		in_6_4_i,
input wire signed [`InBus]		in_6_5_r,
input wire signed [`InBus]		in_6_5_i,
input wire signed [`InBus]		in_6_6_r,
input wire signed [`InBus]		in_6_6_i,
input wire signed [`InBus]		in_6_7_r,
input wire signed [`InBus]		in_6_7_i,
input wire signed [`InBus]		in_6_8_r,
input wire signed [`InBus]		in_6_8_i,
input wire signed [`InBus]		in_7_1_r,
input wire signed [`InBus]		in_7_1_i,
input wire signed [`InBus]		in_7_2_r,
input wire signed [`InBus]		in_7_2_i,
input wire signed [`InBus]		in_7_3_r,
input wire signed [`InBus]		in_7_3_i,
input wire signed [`InBus]		in_7_4_r,
input wire signed [`InBus]		in_7_4_i,
input wire signed [`InBus]		in_7_5_r,
input wire signed [`InBus]		in_7_5_i,
input wire signed [`InBus]		in_7_6_r,
input wire signed [`InBus]		in_7_6_i,
input wire signed [`InBus]		in_7_7_r,
input wire signed [`InBus]		in_7_7_i,
input wire signed [`InBus]		in_7_8_r,
input wire signed [`InBus]		in_7_8_i,
input wire signed [`InBus]		in_8_1_r,
input wire signed [`InBus]		in_8_1_i,
input wire signed [`InBus]		in_8_2_r,
input wire signed [`InBus]		in_8_2_i,
input wire signed [`InBus]		in_8_3_r,
input wire signed [`InBus]		in_8_3_i,
input wire signed [`InBus]		in_8_4_r,
input wire signed [`InBus]		in_8_4_i,
input wire signed [`InBus]		in_8_5_r,
input wire signed [`InBus]		in_8_5_i,
input wire signed [`InBus]		in_8_6_r,
input wire signed [`InBus]		in_8_6_i,
input wire signed [`InBus]		in_8_7_r,
input wire signed [`InBus]		in_8_7_i,
input wire signed [`InBus]		in_8_8_r,
input wire signed [`InBus]		in_8_8_i,

output wire signed [`OutBus]		out_1_1_r,
output wire signed [`OutBus]		out_1_1_i,
output wire signed [`OutBus]		out_1_2_r,
output wire signed [`OutBus]		out_1_2_i,
output wire signed [`OutBus]		out_1_3_r,
output wire signed [`OutBus]		out_1_3_i,
output wire signed [`OutBus]		out_1_4_r,
output wire signed [`OutBus]		out_1_4_i,
output wire signed [`OutBus]		out_1_5_r,
output wire signed [`OutBus]		out_1_5_i,
output wire signed [`OutBus]		out_1_6_r,
output wire signed [`OutBus]		out_1_6_i,
output wire signed [`OutBus]		out_1_7_r,
output wire signed [`OutBus]		out_1_7_i,
output wire signed [`OutBus]		out_1_8_r,
output wire signed [`OutBus]		out_1_8_i,
output wire signed [`OutBus]		out_2_1_r,
output wire signed [`OutBus]		out_2_1_i,
output wire signed [`OutBus]		out_2_2_r,
output wire signed [`OutBus]		out_2_2_i,
output wire signed [`OutBus]		out_2_3_r,
output wire signed [`OutBus]		out_2_3_i,
output wire signed [`OutBus]		out_2_4_r,
output wire signed [`OutBus]		out_2_4_i,
output wire signed [`OutBus]		out_2_5_r,
output wire signed [`OutBus]		out_2_5_i,
output wire signed [`OutBus]		out_2_6_r,
output wire signed [`OutBus]		out_2_6_i,
output wire signed [`OutBus]		out_2_7_r,
output wire signed [`OutBus]		out_2_7_i,
output wire signed [`OutBus]		out_2_8_r,
output wire signed [`OutBus]		out_2_8_i,
output wire signed [`OutBus]		out_3_1_r,
output wire signed [`OutBus]		out_3_1_i,
output wire signed [`OutBus]		out_3_2_r,
output wire signed [`OutBus]		out_3_2_i,
output wire signed [`OutBus]		out_3_3_r,
output wire signed [`OutBus]		out_3_3_i,
output wire signed [`OutBus]		out_3_4_r,
output wire signed [`OutBus]		out_3_4_i,
output wire signed [`OutBus]		out_3_5_r,
output wire signed [`OutBus]		out_3_5_i,
output wire signed [`OutBus]		out_3_6_r,
output wire signed [`OutBus]		out_3_6_i,
output wire signed [`OutBus]		out_3_7_r,
output wire signed [`OutBus]		out_3_7_i,
output wire signed [`OutBus]		out_3_8_r,
output wire signed [`OutBus]		out_3_8_i,
output wire signed [`OutBus]		out_4_1_r,
output wire signed [`OutBus]		out_4_1_i,
output wire signed [`OutBus]		out_4_2_r,
output wire signed [`OutBus]		out_4_2_i,
output wire signed [`OutBus]		out_4_3_r,
output wire signed [`OutBus]		out_4_3_i,
output wire signed [`OutBus]		out_4_4_r,
output wire signed [`OutBus]		out_4_4_i,
output wire signed [`OutBus]		out_4_5_r,
output wire signed [`OutBus]		out_4_5_i,
output wire signed [`OutBus]		out_4_6_r,
output wire signed [`OutBus]		out_4_6_i,
output wire signed [`OutBus]		out_4_7_r,
output wire signed [`OutBus]		out_4_7_i,
output wire signed [`OutBus]		out_4_8_r,
output wire signed [`OutBus]		out_4_8_i,
output wire signed [`OutBus]		out_5_1_r,
output wire signed [`OutBus]		out_5_1_i,
output wire signed [`OutBus]		out_5_2_r,
output wire signed [`OutBus]		out_5_2_i,
output wire signed [`OutBus]		out_5_3_r,
output wire signed [`OutBus]		out_5_3_i,
output wire signed [`OutBus]		out_5_4_r,
output wire signed [`OutBus]		out_5_4_i,
output wire signed [`OutBus]		out_5_5_r,
output wire signed [`OutBus]		out_5_5_i,
output wire signed [`OutBus]		out_5_6_r,
output wire signed [`OutBus]		out_5_6_i,
output wire signed [`OutBus]		out_5_7_r,
output wire signed [`OutBus]		out_5_7_i,
output wire signed [`OutBus]		out_5_8_r,
output wire signed [`OutBus]		out_5_8_i,
output wire signed [`OutBus]		out_6_1_r,
output wire signed [`OutBus]		out_6_1_i,
output wire signed [`OutBus]		out_6_2_r,
output wire signed [`OutBus]		out_6_2_i,
output wire signed [`OutBus]		out_6_3_r,
output wire signed [`OutBus]		out_6_3_i,
output wire signed [`OutBus]		out_6_4_r,
output wire signed [`OutBus]		out_6_4_i,
output wire signed [`OutBus]		out_6_5_r,
output wire signed [`OutBus]		out_6_5_i,
output wire signed [`OutBus]		out_6_6_r,
output wire signed [`OutBus]		out_6_6_i,
output wire signed [`OutBus]		out_6_7_r,
output wire signed [`OutBus]		out_6_7_i,
output wire signed [`OutBus]		out_6_8_r,
output wire signed [`OutBus]		out_6_8_i,
output wire signed [`OutBus]		out_7_1_r,
output wire signed [`OutBus]		out_7_1_i,
output wire signed [`OutBus]		out_7_2_r,
output wire signed [`OutBus]		out_7_2_i,
output wire signed [`OutBus]		out_7_3_r,
output wire signed [`OutBus]		out_7_3_i,
output wire signed [`OutBus]		out_7_4_r,
output wire signed [`OutBus]		out_7_4_i,
output wire signed [`OutBus]		out_7_5_r,
output wire signed [`OutBus]		out_7_5_i,
output wire signed [`OutBus]		out_7_6_r,
output wire signed [`OutBus]		out_7_6_i,
output wire signed [`OutBus]		out_7_7_r,
output wire signed [`OutBus]		out_7_7_i,
output wire signed [`OutBus]		out_7_8_r,
output wire signed [`OutBus]		out_7_8_i,
output wire signed [`OutBus]		out_8_1_r,
output wire signed [`OutBus]		out_8_1_i,
output wire signed [`OutBus]		out_8_2_r,
output wire signed [`OutBus]		out_8_2_i,
output wire signed [`OutBus]		out_8_3_r,
output wire signed [`OutBus]		out_8_3_i,
output wire signed [`OutBus]		out_8_4_r,
output wire signed [`OutBus]		out_8_4_i,
output wire signed [`OutBus]		out_8_5_r,
output wire signed [`OutBus]		out_8_5_i,
output wire signed [`OutBus]		out_8_6_r,
output wire signed [`OutBus]		out_8_6_i,
output wire signed [`OutBus]		out_8_7_r,
output wire signed [`OutBus]		out_8_7_i,
output wire signed [`OutBus]		out_8_8_r,
output wire signed [`OutBus]		out_8_8_i

);

wire signed [`CalcTempBus]          temp_m1_1_1_r;
wire signed [`CalcTempBus]          temp_m1_1_1_i;
wire signed [`CalcTempBus]          temp_m1_1_2_r;
wire signed [`CalcTempBus]          temp_m1_1_2_i;
wire signed [`CalcTempBus]          temp_m1_1_3_r;
wire signed [`CalcTempBus]          temp_m1_1_3_i;
wire signed [`CalcTempBus]          temp_m1_1_4_r;
wire signed [`CalcTempBus]          temp_m1_1_4_i;
wire signed [`CalcTempBus]          temp_m1_1_5_r;
wire signed [`CalcTempBus]          temp_m1_1_5_i;
wire signed [`CalcTempBus]          temp_m1_1_6_r;
wire signed [`CalcTempBus]          temp_m1_1_6_i;
wire signed [`CalcTempBus]          temp_m1_1_7_r;
wire signed [`CalcTempBus]          temp_m1_1_7_i;
wire signed [`CalcTempBus]          temp_m1_1_8_r;
wire signed [`CalcTempBus]          temp_m1_1_8_i;
wire signed [`CalcTempBus]          temp_m1_2_1_r;
wire signed [`CalcTempBus]          temp_m1_2_1_i;
wire signed [`CalcTempBus]          temp_m1_2_2_r;
wire signed [`CalcTempBus]          temp_m1_2_2_i;
wire signed [`CalcTempBus]          temp_m1_2_3_r;
wire signed [`CalcTempBus]          temp_m1_2_3_i;
wire signed [`CalcTempBus]          temp_m1_2_4_r;
wire signed [`CalcTempBus]          temp_m1_2_4_i;
wire signed [`CalcTempBus]          temp_m1_2_5_r;
wire signed [`CalcTempBus]          temp_m1_2_5_i;
wire signed [`CalcTempBus]          temp_m1_2_6_r;
wire signed [`CalcTempBus]          temp_m1_2_6_i;
wire signed [`CalcTempBus]          temp_m1_2_7_r;
wire signed [`CalcTempBus]          temp_m1_2_7_i;
wire signed [`CalcTempBus]          temp_m1_2_8_r;
wire signed [`CalcTempBus]          temp_m1_2_8_i;
wire signed [`CalcTempBus]          temp_m1_3_1_r;
wire signed [`CalcTempBus]          temp_m1_3_1_i;
wire signed [`CalcTempBus]          temp_m1_3_2_r;
wire signed [`CalcTempBus]          temp_m1_3_2_i;
wire signed [`CalcTempBus]          temp_m1_3_3_r;
wire signed [`CalcTempBus]          temp_m1_3_3_i;
wire signed [`CalcTempBus]          temp_m1_3_4_r;
wire signed [`CalcTempBus]          temp_m1_3_4_i;
wire signed [`CalcTempBus]          temp_m1_3_5_r;
wire signed [`CalcTempBus]          temp_m1_3_5_i;
wire signed [`CalcTempBus]          temp_m1_3_6_r;
wire signed [`CalcTempBus]          temp_m1_3_6_i;
wire signed [`CalcTempBus]          temp_m1_3_7_r;
wire signed [`CalcTempBus]          temp_m1_3_7_i;
wire signed [`CalcTempBus]          temp_m1_3_8_r;
wire signed [`CalcTempBus]          temp_m1_3_8_i;
wire signed [`CalcTempBus]          temp_m1_4_1_r;
wire signed [`CalcTempBus]          temp_m1_4_1_i;
wire signed [`CalcTempBus]          temp_m1_4_2_r;
wire signed [`CalcTempBus]          temp_m1_4_2_i;
wire signed [`CalcTempBus]          temp_m1_4_3_r;
wire signed [`CalcTempBus]          temp_m1_4_3_i;
wire signed [`CalcTempBus]          temp_m1_4_4_r;
wire signed [`CalcTempBus]          temp_m1_4_4_i;
wire signed [`CalcTempBus]          temp_m1_4_5_r;
wire signed [`CalcTempBus]          temp_m1_4_5_i;
wire signed [`CalcTempBus]          temp_m1_4_6_r;
wire signed [`CalcTempBus]          temp_m1_4_6_i;
wire signed [`CalcTempBus]          temp_m1_4_7_r;
wire signed [`CalcTempBus]          temp_m1_4_7_i;
wire signed [`CalcTempBus]          temp_m1_4_8_r;
wire signed [`CalcTempBus]          temp_m1_4_8_i;
wire signed [`CalcTempBus]          temp_m1_5_1_r;
wire signed [`CalcTempBus]          temp_m1_5_1_i;
wire signed [`CalcTempBus]          temp_m1_5_2_r;
wire signed [`CalcTempBus]          temp_m1_5_2_i;
wire signed [`CalcTempBus]          temp_m1_5_3_r;
wire signed [`CalcTempBus]          temp_m1_5_3_i;
wire signed [`CalcTempBus]          temp_m1_5_4_r;
wire signed [`CalcTempBus]          temp_m1_5_4_i;
wire signed [`CalcTempBus]          temp_m1_5_5_r;
wire signed [`CalcTempBus]          temp_m1_5_5_i;
wire signed [`CalcTempBus]          temp_m1_5_6_r;
wire signed [`CalcTempBus]          temp_m1_5_6_i;
wire signed [`CalcTempBus]          temp_m1_5_7_r;
wire signed [`CalcTempBus]          temp_m1_5_7_i;
wire signed [`CalcTempBus]          temp_m1_5_8_r;
wire signed [`CalcTempBus]          temp_m1_5_8_i;
wire signed [`CalcTempBus]          temp_m1_6_1_r;
wire signed [`CalcTempBus]          temp_m1_6_1_i;
wire signed [`CalcTempBus]          temp_m1_6_2_r;
wire signed [`CalcTempBus]          temp_m1_6_2_i;
wire signed [`CalcTempBus]          temp_m1_6_3_r;
wire signed [`CalcTempBus]          temp_m1_6_3_i;
wire signed [`CalcTempBus]          temp_m1_6_4_r;
wire signed [`CalcTempBus]          temp_m1_6_4_i;
wire signed [`CalcTempBus]          temp_m1_6_5_r;
wire signed [`CalcTempBus]          temp_m1_6_5_i;
wire signed [`CalcTempBus]          temp_m1_6_6_r;
wire signed [`CalcTempBus]          temp_m1_6_6_i;
wire signed [`CalcTempBus]          temp_m1_6_7_r;
wire signed [`CalcTempBus]          temp_m1_6_7_i;
wire signed [`CalcTempBus]          temp_m1_6_8_r;
wire signed [`CalcTempBus]          temp_m1_6_8_i;
wire signed [`CalcTempBus]          temp_m1_7_1_r;
wire signed [`CalcTempBus]          temp_m1_7_1_i;
wire signed [`CalcTempBus]          temp_m1_7_2_r;
wire signed [`CalcTempBus]          temp_m1_7_2_i;
wire signed [`CalcTempBus]          temp_m1_7_3_r;
wire signed [`CalcTempBus]          temp_m1_7_3_i;
wire signed [`CalcTempBus]          temp_m1_7_4_r;
wire signed [`CalcTempBus]          temp_m1_7_4_i;
wire signed [`CalcTempBus]          temp_m1_7_5_r;
wire signed [`CalcTempBus]          temp_m1_7_5_i;
wire signed [`CalcTempBus]          temp_m1_7_6_r;
wire signed [`CalcTempBus]          temp_m1_7_6_i;
wire signed [`CalcTempBus]          temp_m1_7_7_r;
wire signed [`CalcTempBus]          temp_m1_7_7_i;
wire signed [`CalcTempBus]          temp_m1_7_8_r;
wire signed [`CalcTempBus]          temp_m1_7_8_i;
wire signed [`CalcTempBus]          temp_m1_8_1_r;
wire signed [`CalcTempBus]          temp_m1_8_1_i;
wire signed [`CalcTempBus]          temp_m1_8_2_r;
wire signed [`CalcTempBus]          temp_m1_8_2_i;
wire signed [`CalcTempBus]          temp_m1_8_3_r;
wire signed [`CalcTempBus]          temp_m1_8_3_i;
wire signed [`CalcTempBus]          temp_m1_8_4_r;
wire signed [`CalcTempBus]          temp_m1_8_4_i;
wire signed [`CalcTempBus]          temp_m1_8_5_r;
wire signed [`CalcTempBus]          temp_m1_8_5_i;
wire signed [`CalcTempBus]          temp_m1_8_6_r;
wire signed [`CalcTempBus]          temp_m1_8_6_i;
wire signed [`CalcTempBus]          temp_m1_8_7_r;
wire signed [`CalcTempBus]          temp_m1_8_7_i;
wire signed [`CalcTempBus]          temp_m1_8_8_r;
wire signed [`CalcTempBus]          temp_m1_8_8_i;
wire signed [`CalcTempBus]          temp_m2_1_1_r;
wire signed [`CalcTempBus]          temp_m2_1_1_i;
wire signed [`CalcTempBus]          temp_m2_1_2_r;
wire signed [`CalcTempBus]          temp_m2_1_2_i;
wire signed [`CalcTempBus]          temp_m2_1_3_r;
wire signed [`CalcTempBus]          temp_m2_1_3_i;
wire signed [`CalcTempBus]          temp_m2_1_4_r;
wire signed [`CalcTempBus]          temp_m2_1_4_i;
wire signed [`CalcTempBus]          temp_m2_1_5_r;
wire signed [`CalcTempBus]          temp_m2_1_5_i;
wire signed [`CalcTempBus]          temp_m2_1_6_r;
wire signed [`CalcTempBus]          temp_m2_1_6_i;
wire signed [`CalcTempBus]          temp_m2_1_7_r;
wire signed [`CalcTempBus]          temp_m2_1_7_i;
wire signed [`CalcTempBus]          temp_m2_1_8_r;
wire signed [`CalcTempBus]          temp_m2_1_8_i;
wire signed [`CalcTempBus]          temp_m2_2_1_r;
wire signed [`CalcTempBus]          temp_m2_2_1_i;
wire signed [`CalcTempBus]          temp_m2_2_2_r;
wire signed [`CalcTempBus]          temp_m2_2_2_i;
wire signed [`CalcTempBus]          temp_m2_2_3_r;
wire signed [`CalcTempBus]          temp_m2_2_3_i;
wire signed [`CalcTempBus]          temp_m2_2_4_r;
wire signed [`CalcTempBus]          temp_m2_2_4_i;
wire signed [`CalcTempBus]          temp_m2_2_5_r;
wire signed [`CalcTempBus]          temp_m2_2_5_i;
wire signed [`CalcTempBus]          temp_m2_2_6_r;
wire signed [`CalcTempBus]          temp_m2_2_6_i;
wire signed [`CalcTempBus]          temp_m2_2_7_r;
wire signed [`CalcTempBus]          temp_m2_2_7_i;
wire signed [`CalcTempBus]          temp_m2_2_8_r;
wire signed [`CalcTempBus]          temp_m2_2_8_i;
wire signed [`CalcTempBus]          temp_m2_3_1_r;
wire signed [`CalcTempBus]          temp_m2_3_1_i;
wire signed [`CalcTempBus]          temp_m2_3_2_r;
wire signed [`CalcTempBus]          temp_m2_3_2_i;
wire signed [`CalcTempBus]          temp_m2_3_3_r;
wire signed [`CalcTempBus]          temp_m2_3_3_i;
wire signed [`CalcTempBus]          temp_m2_3_4_r;
wire signed [`CalcTempBus]          temp_m2_3_4_i;
wire signed [`CalcTempBus]          temp_m2_3_5_r;
wire signed [`CalcTempBus]          temp_m2_3_5_i;
wire signed [`CalcTempBus]          temp_m2_3_6_r;
wire signed [`CalcTempBus]          temp_m2_3_6_i;
wire signed [`CalcTempBus]          temp_m2_3_7_r;
wire signed [`CalcTempBus]          temp_m2_3_7_i;
wire signed [`CalcTempBus]          temp_m2_3_8_r;
wire signed [`CalcTempBus]          temp_m2_3_8_i;
wire signed [`CalcTempBus]          temp_m2_4_1_r;
wire signed [`CalcTempBus]          temp_m2_4_1_i;
wire signed [`CalcTempBus]          temp_m2_4_2_r;
wire signed [`CalcTempBus]          temp_m2_4_2_i;
wire signed [`CalcTempBus]          temp_m2_4_3_r;
wire signed [`CalcTempBus]          temp_m2_4_3_i;
wire signed [`CalcTempBus]          temp_m2_4_4_r;
wire signed [`CalcTempBus]          temp_m2_4_4_i;
wire signed [`CalcTempBus]          temp_m2_4_5_r;
wire signed [`CalcTempBus]          temp_m2_4_5_i;
wire signed [`CalcTempBus]          temp_m2_4_6_r;
wire signed [`CalcTempBus]          temp_m2_4_6_i;
wire signed [`CalcTempBus]          temp_m2_4_7_r;
wire signed [`CalcTempBus]          temp_m2_4_7_i;
wire signed [`CalcTempBus]          temp_m2_4_8_r;
wire signed [`CalcTempBus]          temp_m2_4_8_i;
wire signed [`CalcTempBus]          temp_m2_5_1_r;
wire signed [`CalcTempBus]          temp_m2_5_1_i;
wire signed [`CalcTempBus]          temp_m2_5_2_r;
wire signed [`CalcTempBus]          temp_m2_5_2_i;
wire signed [`CalcTempBus]          temp_m2_5_3_r;
wire signed [`CalcTempBus]          temp_m2_5_3_i;
wire signed [`CalcTempBus]          temp_m2_5_4_r;
wire signed [`CalcTempBus]          temp_m2_5_4_i;
wire signed [`CalcTempBus]          temp_m2_5_5_r;
wire signed [`CalcTempBus]          temp_m2_5_5_i;
wire signed [`CalcTempBus]          temp_m2_5_6_r;
wire signed [`CalcTempBus]          temp_m2_5_6_i;
wire signed [`CalcTempBus]          temp_m2_5_7_r;
wire signed [`CalcTempBus]          temp_m2_5_7_i;
wire signed [`CalcTempBus]          temp_m2_5_8_r;
wire signed [`CalcTempBus]          temp_m2_5_8_i;
wire signed [`CalcTempBus]          temp_m2_6_1_r;
wire signed [`CalcTempBus]          temp_m2_6_1_i;
wire signed [`CalcTempBus]          temp_m2_6_2_r;
wire signed [`CalcTempBus]          temp_m2_6_2_i;
wire signed [`CalcTempBus]          temp_m2_6_3_r;
wire signed [`CalcTempBus]          temp_m2_6_3_i;
wire signed [`CalcTempBus]          temp_m2_6_4_r;
wire signed [`CalcTempBus]          temp_m2_6_4_i;
wire signed [`CalcTempBus]          temp_m2_6_5_r;
wire signed [`CalcTempBus]          temp_m2_6_5_i;
wire signed [`CalcTempBus]          temp_m2_6_6_r;
wire signed [`CalcTempBus]          temp_m2_6_6_i;
wire signed [`CalcTempBus]          temp_m2_6_7_r;
wire signed [`CalcTempBus]          temp_m2_6_7_i;
wire signed [`CalcTempBus]          temp_m2_6_8_r;
wire signed [`CalcTempBus]          temp_m2_6_8_i;
wire signed [`CalcTempBus]          temp_m2_7_1_r;
wire signed [`CalcTempBus]          temp_m2_7_1_i;
wire signed [`CalcTempBus]          temp_m2_7_2_r;
wire signed [`CalcTempBus]          temp_m2_7_2_i;
wire signed [`CalcTempBus]          temp_m2_7_3_r;
wire signed [`CalcTempBus]          temp_m2_7_3_i;
wire signed [`CalcTempBus]          temp_m2_7_4_r;
wire signed [`CalcTempBus]          temp_m2_7_4_i;
wire signed [`CalcTempBus]          temp_m2_7_5_r;
wire signed [`CalcTempBus]          temp_m2_7_5_i;
wire signed [`CalcTempBus]          temp_m2_7_6_r;
wire signed [`CalcTempBus]          temp_m2_7_6_i;
wire signed [`CalcTempBus]          temp_m2_7_7_r;
wire signed [`CalcTempBus]          temp_m2_7_7_i;
wire signed [`CalcTempBus]          temp_m2_7_8_r;
wire signed [`CalcTempBus]          temp_m2_7_8_i;
wire signed [`CalcTempBus]          temp_m2_8_1_r;
wire signed [`CalcTempBus]          temp_m2_8_1_i;
wire signed [`CalcTempBus]          temp_m2_8_2_r;
wire signed [`CalcTempBus]          temp_m2_8_2_i;
wire signed [`CalcTempBus]          temp_m2_8_3_r;
wire signed [`CalcTempBus]          temp_m2_8_3_i;
wire signed [`CalcTempBus]          temp_m2_8_4_r;
wire signed [`CalcTempBus]          temp_m2_8_4_i;
wire signed [`CalcTempBus]          temp_m2_8_5_r;
wire signed [`CalcTempBus]          temp_m2_8_5_i;
wire signed [`CalcTempBus]          temp_m2_8_6_r;
wire signed [`CalcTempBus]          temp_m2_8_6_i;
wire signed [`CalcTempBus]          temp_m2_8_7_r;
wire signed [`CalcTempBus]          temp_m2_8_7_i;
wire signed [`CalcTempBus]          temp_m2_8_8_r;
wire signed [`CalcTempBus]          temp_m2_8_8_i;
wire signed [`CalcTempBus]          temp_m3_1_1_r;
wire signed [`CalcTempBus]          temp_m3_1_1_i;
wire signed [`CalcTempBus]          temp_m3_1_2_r;
wire signed [`CalcTempBus]          temp_m3_1_2_i;
wire signed [`CalcTempBus]          temp_m3_1_3_r;
wire signed [`CalcTempBus]          temp_m3_1_3_i;
wire signed [`CalcTempBus]          temp_m3_1_4_r;
wire signed [`CalcTempBus]          temp_m3_1_4_i;
wire signed [`CalcTempBus]          temp_m3_1_5_r;
wire signed [`CalcTempBus]          temp_m3_1_5_i;
wire signed [`CalcTempBus]          temp_m3_1_6_r;
wire signed [`CalcTempBus]          temp_m3_1_6_i;
wire signed [`CalcTempBus]          temp_m3_1_7_r;
wire signed [`CalcTempBus]          temp_m3_1_7_i;
wire signed [`CalcTempBus]          temp_m3_1_8_r;
wire signed [`CalcTempBus]          temp_m3_1_8_i;
wire signed [`CalcTempBus]          temp_m3_2_1_r;
wire signed [`CalcTempBus]          temp_m3_2_1_i;
wire signed [`CalcTempBus]          temp_m3_2_2_r;
wire signed [`CalcTempBus]          temp_m3_2_2_i;
wire signed [`CalcTempBus]          temp_m3_2_3_r;
wire signed [`CalcTempBus]          temp_m3_2_3_i;
wire signed [`CalcTempBus]          temp_m3_2_4_r;
wire signed [`CalcTempBus]          temp_m3_2_4_i;
wire signed [`CalcTempBus]          temp_m3_2_5_r;
wire signed [`CalcTempBus]          temp_m3_2_5_i;
wire signed [`CalcTempBus]          temp_m3_2_6_r;
wire signed [`CalcTempBus]          temp_m3_2_6_i;
wire signed [`CalcTempBus]          temp_m3_2_7_r;
wire signed [`CalcTempBus]          temp_m3_2_7_i;
wire signed [`CalcTempBus]          temp_m3_2_8_r;
wire signed [`CalcTempBus]          temp_m3_2_8_i;
wire signed [`CalcTempBus]          temp_m3_3_1_r;
wire signed [`CalcTempBus]          temp_m3_3_1_i;
wire signed [`CalcTempBus]          temp_m3_3_2_r;
wire signed [`CalcTempBus]          temp_m3_3_2_i;
wire signed [`CalcTempBus]          temp_m3_3_3_r;
wire signed [`CalcTempBus]          temp_m3_3_3_i;
wire signed [`CalcTempBus]          temp_m3_3_4_r;
wire signed [`CalcTempBus]          temp_m3_3_4_i;
wire signed [`CalcTempBus]          temp_m3_3_5_r;
wire signed [`CalcTempBus]          temp_m3_3_5_i;
wire signed [`CalcTempBus]          temp_m3_3_6_r;
wire signed [`CalcTempBus]          temp_m3_3_6_i;
wire signed [`CalcTempBus]          temp_m3_3_7_r;
wire signed [`CalcTempBus]          temp_m3_3_7_i;
wire signed [`CalcTempBus]          temp_m3_3_8_r;
wire signed [`CalcTempBus]          temp_m3_3_8_i;
wire signed [`CalcTempBus]          temp_m3_4_1_r;
wire signed [`CalcTempBus]          temp_m3_4_1_i;
wire signed [`CalcTempBus]          temp_m3_4_2_r;
wire signed [`CalcTempBus]          temp_m3_4_2_i;
wire signed [`CalcTempBus]          temp_m3_4_3_r;
wire signed [`CalcTempBus]          temp_m3_4_3_i;
wire signed [`CalcTempBus]          temp_m3_4_4_r;
wire signed [`CalcTempBus]          temp_m3_4_4_i;
wire signed [`CalcTempBus]          temp_m3_4_5_r;
wire signed [`CalcTempBus]          temp_m3_4_5_i;
wire signed [`CalcTempBus]          temp_m3_4_6_r;
wire signed [`CalcTempBus]          temp_m3_4_6_i;
wire signed [`CalcTempBus]          temp_m3_4_7_r;
wire signed [`CalcTempBus]          temp_m3_4_7_i;
wire signed [`CalcTempBus]          temp_m3_4_8_r;
wire signed [`CalcTempBus]          temp_m3_4_8_i;
wire signed [`CalcTempBus]          temp_m3_5_1_r;
wire signed [`CalcTempBus]          temp_m3_5_1_i;
wire signed [`CalcTempBus]          temp_m3_5_2_r;
wire signed [`CalcTempBus]          temp_m3_5_2_i;
wire signed [`CalcTempBus]          temp_m3_5_3_r;
wire signed [`CalcTempBus]          temp_m3_5_3_i;
wire signed [`CalcTempBus]          temp_m3_5_4_r;
wire signed [`CalcTempBus]          temp_m3_5_4_i;
wire signed [`CalcTempBus]          temp_m3_5_5_r;
wire signed [`CalcTempBus]          temp_m3_5_5_i;
wire signed [`CalcTempBus]          temp_m3_5_6_r;
wire signed [`CalcTempBus]          temp_m3_5_6_i;
wire signed [`CalcTempBus]          temp_m3_5_7_r;
wire signed [`CalcTempBus]          temp_m3_5_7_i;
wire signed [`CalcTempBus]          temp_m3_5_8_r;
wire signed [`CalcTempBus]          temp_m3_5_8_i;
wire signed [`CalcTempBus]          temp_m3_6_1_r;
wire signed [`CalcTempBus]          temp_m3_6_1_i;
wire signed [`CalcTempBus]          temp_m3_6_2_r;
wire signed [`CalcTempBus]          temp_m3_6_2_i;
wire signed [`CalcTempBus]          temp_m3_6_3_r;
wire signed [`CalcTempBus]          temp_m3_6_3_i;
wire signed [`CalcTempBus]          temp_m3_6_4_r;
wire signed [`CalcTempBus]          temp_m3_6_4_i;
wire signed [`CalcTempBus]          temp_m3_6_5_r;
wire signed [`CalcTempBus]          temp_m3_6_5_i;
wire signed [`CalcTempBus]          temp_m3_6_6_r;
wire signed [`CalcTempBus]          temp_m3_6_6_i;
wire signed [`CalcTempBus]          temp_m3_6_7_r;
wire signed [`CalcTempBus]          temp_m3_6_7_i;
wire signed [`CalcTempBus]          temp_m3_6_8_r;
wire signed [`CalcTempBus]          temp_m3_6_8_i;
wire signed [`CalcTempBus]          temp_m3_7_1_r;
wire signed [`CalcTempBus]          temp_m3_7_1_i;
wire signed [`CalcTempBus]          temp_m3_7_2_r;
wire signed [`CalcTempBus]          temp_m3_7_2_i;
wire signed [`CalcTempBus]          temp_m3_7_3_r;
wire signed [`CalcTempBus]          temp_m3_7_3_i;
wire signed [`CalcTempBus]          temp_m3_7_4_r;
wire signed [`CalcTempBus]          temp_m3_7_4_i;
wire signed [`CalcTempBus]          temp_m3_7_5_r;
wire signed [`CalcTempBus]          temp_m3_7_5_i;
wire signed [`CalcTempBus]          temp_m3_7_6_r;
wire signed [`CalcTempBus]          temp_m3_7_6_i;
wire signed [`CalcTempBus]          temp_m3_7_7_r;
wire signed [`CalcTempBus]          temp_m3_7_7_i;
wire signed [`CalcTempBus]          temp_m3_7_8_r;
wire signed [`CalcTempBus]          temp_m3_7_8_i;
wire signed [`CalcTempBus]          temp_m3_8_1_r;
wire signed [`CalcTempBus]          temp_m3_8_1_i;
wire signed [`CalcTempBus]          temp_m3_8_2_r;
wire signed [`CalcTempBus]          temp_m3_8_2_i;
wire signed [`CalcTempBus]          temp_m3_8_3_r;
wire signed [`CalcTempBus]          temp_m3_8_3_i;
wire signed [`CalcTempBus]          temp_m3_8_4_r;
wire signed [`CalcTempBus]          temp_m3_8_4_i;
wire signed [`CalcTempBus]          temp_m3_8_5_r;
wire signed [`CalcTempBus]          temp_m3_8_5_i;
wire signed [`CalcTempBus]          temp_m3_8_6_r;
wire signed [`CalcTempBus]          temp_m3_8_6_i;
wire signed [`CalcTempBus]          temp_m3_8_7_r;
wire signed [`CalcTempBus]          temp_m3_8_7_i;
wire signed [`CalcTempBus]          temp_m3_8_8_r;
wire signed [`CalcTempBus]          temp_m3_8_8_i;

wire signed [`CalcTempBus]          temp_b1_1_1_r;
wire signed [`CalcTempBus]          temp_b1_1_1_i;
wire signed [`CalcTempBus]          temp_b1_1_2_r;
wire signed [`CalcTempBus]          temp_b1_1_2_i;
wire signed [`CalcTempBus]          temp_b1_1_3_r;
wire signed [`CalcTempBus]          temp_b1_1_3_i;
wire signed [`CalcTempBus]          temp_b1_1_4_r;
wire signed [`CalcTempBus]          temp_b1_1_4_i;
wire signed [`CalcTempBus]          temp_b1_1_5_r;
wire signed [`CalcTempBus]          temp_b1_1_5_i;
wire signed [`CalcTempBus]          temp_b1_1_6_r;
wire signed [`CalcTempBus]          temp_b1_1_6_i;
wire signed [`CalcTempBus]          temp_b1_1_7_r;
wire signed [`CalcTempBus]          temp_b1_1_7_i;
wire signed [`CalcTempBus]          temp_b1_1_8_r;
wire signed [`CalcTempBus]          temp_b1_1_8_i;
wire signed [`CalcTempBus]          temp_b1_2_1_r;
wire signed [`CalcTempBus]          temp_b1_2_1_i;
wire signed [`CalcTempBus]          temp_b1_2_2_r;
wire signed [`CalcTempBus]          temp_b1_2_2_i;
wire signed [`CalcTempBus]          temp_b1_2_3_r;
wire signed [`CalcTempBus]          temp_b1_2_3_i;
wire signed [`CalcTempBus]          temp_b1_2_4_r;
wire signed [`CalcTempBus]          temp_b1_2_4_i;
wire signed [`CalcTempBus]          temp_b1_2_5_r;
wire signed [`CalcTempBus]          temp_b1_2_5_i;
wire signed [`CalcTempBus]          temp_b1_2_6_r;
wire signed [`CalcTempBus]          temp_b1_2_6_i;
wire signed [`CalcTempBus]          temp_b1_2_7_r;
wire signed [`CalcTempBus]          temp_b1_2_7_i;
wire signed [`CalcTempBus]          temp_b1_2_8_r;
wire signed [`CalcTempBus]          temp_b1_2_8_i;
wire signed [`CalcTempBus]          temp_b1_3_1_r;
wire signed [`CalcTempBus]          temp_b1_3_1_i;
wire signed [`CalcTempBus]          temp_b1_3_2_r;
wire signed [`CalcTempBus]          temp_b1_3_2_i;
wire signed [`CalcTempBus]          temp_b1_3_3_r;
wire signed [`CalcTempBus]          temp_b1_3_3_i;
wire signed [`CalcTempBus]          temp_b1_3_4_r;
wire signed [`CalcTempBus]          temp_b1_3_4_i;
wire signed [`CalcTempBus]          temp_b1_3_5_r;
wire signed [`CalcTempBus]          temp_b1_3_5_i;
wire signed [`CalcTempBus]          temp_b1_3_6_r;
wire signed [`CalcTempBus]          temp_b1_3_6_i;
wire signed [`CalcTempBus]          temp_b1_3_7_r;
wire signed [`CalcTempBus]          temp_b1_3_7_i;
wire signed [`CalcTempBus]          temp_b1_3_8_r;
wire signed [`CalcTempBus]          temp_b1_3_8_i;
wire signed [`CalcTempBus]          temp_b1_4_1_r;
wire signed [`CalcTempBus]          temp_b1_4_1_i;
wire signed [`CalcTempBus]          temp_b1_4_2_r;
wire signed [`CalcTempBus]          temp_b1_4_2_i;
wire signed [`CalcTempBus]          temp_b1_4_3_r;
wire signed [`CalcTempBus]          temp_b1_4_3_i;
wire signed [`CalcTempBus]          temp_b1_4_4_r;
wire signed [`CalcTempBus]          temp_b1_4_4_i;
wire signed [`CalcTempBus]          temp_b1_4_5_r;
wire signed [`CalcTempBus]          temp_b1_4_5_i;
wire signed [`CalcTempBus]          temp_b1_4_6_r;
wire signed [`CalcTempBus]          temp_b1_4_6_i;
wire signed [`CalcTempBus]          temp_b1_4_7_r;
wire signed [`CalcTempBus]          temp_b1_4_7_i;
wire signed [`CalcTempBus]          temp_b1_4_8_r;
wire signed [`CalcTempBus]          temp_b1_4_8_i;
wire signed [`CalcTempBus]          temp_b1_5_1_r;
wire signed [`CalcTempBus]          temp_b1_5_1_i;
wire signed [`CalcTempBus]          temp_b1_5_2_r;
wire signed [`CalcTempBus]          temp_b1_5_2_i;
wire signed [`CalcTempBus]          temp_b1_5_3_r;
wire signed [`CalcTempBus]          temp_b1_5_3_i;
wire signed [`CalcTempBus]          temp_b1_5_4_r;
wire signed [`CalcTempBus]          temp_b1_5_4_i;
wire signed [`CalcTempBus]          temp_b1_5_5_r;
wire signed [`CalcTempBus]          temp_b1_5_5_i;
wire signed [`CalcTempBus]          temp_b1_5_6_r;
wire signed [`CalcTempBus]          temp_b1_5_6_i;
wire signed [`CalcTempBus]          temp_b1_5_7_r;
wire signed [`CalcTempBus]          temp_b1_5_7_i;
wire signed [`CalcTempBus]          temp_b1_5_8_r;
wire signed [`CalcTempBus]          temp_b1_5_8_i;
wire signed [`CalcTempBus]          temp_b1_6_1_r;
wire signed [`CalcTempBus]          temp_b1_6_1_i;
wire signed [`CalcTempBus]          temp_b1_6_2_r;
wire signed [`CalcTempBus]          temp_b1_6_2_i;
wire signed [`CalcTempBus]          temp_b1_6_3_r;
wire signed [`CalcTempBus]          temp_b1_6_3_i;
wire signed [`CalcTempBus]          temp_b1_6_4_r;
wire signed [`CalcTempBus]          temp_b1_6_4_i;
wire signed [`CalcTempBus]          temp_b1_6_5_r;
wire signed [`CalcTempBus]          temp_b1_6_5_i;
wire signed [`CalcTempBus]          temp_b1_6_6_r;
wire signed [`CalcTempBus]          temp_b1_6_6_i;
wire signed [`CalcTempBus]          temp_b1_6_7_r;
wire signed [`CalcTempBus]          temp_b1_6_7_i;
wire signed [`CalcTempBus]          temp_b1_6_8_r;
wire signed [`CalcTempBus]          temp_b1_6_8_i;
wire signed [`CalcTempBus]          temp_b1_7_1_r;
wire signed [`CalcTempBus]          temp_b1_7_1_i;
wire signed [`CalcTempBus]          temp_b1_7_2_r;
wire signed [`CalcTempBus]          temp_b1_7_2_i;
wire signed [`CalcTempBus]          temp_b1_7_3_r;
wire signed [`CalcTempBus]          temp_b1_7_3_i;
wire signed [`CalcTempBus]          temp_b1_7_4_r;
wire signed [`CalcTempBus]          temp_b1_7_4_i;
wire signed [`CalcTempBus]          temp_b1_7_5_r;
wire signed [`CalcTempBus]          temp_b1_7_5_i;
wire signed [`CalcTempBus]          temp_b1_7_6_r;
wire signed [`CalcTempBus]          temp_b1_7_6_i;
wire signed [`CalcTempBus]          temp_b1_7_7_r;
wire signed [`CalcTempBus]          temp_b1_7_7_i;
wire signed [`CalcTempBus]          temp_b1_7_8_r;
wire signed [`CalcTempBus]          temp_b1_7_8_i;
wire signed [`CalcTempBus]          temp_b1_8_1_r;
wire signed [`CalcTempBus]          temp_b1_8_1_i;
wire signed [`CalcTempBus]          temp_b1_8_2_r;
wire signed [`CalcTempBus]          temp_b1_8_2_i;
wire signed [`CalcTempBus]          temp_b1_8_3_r;
wire signed [`CalcTempBus]          temp_b1_8_3_i;
wire signed [`CalcTempBus]          temp_b1_8_4_r;
wire signed [`CalcTempBus]          temp_b1_8_4_i;
wire signed [`CalcTempBus]          temp_b1_8_5_r;
wire signed [`CalcTempBus]          temp_b1_8_5_i;
wire signed [`CalcTempBus]          temp_b1_8_6_r;
wire signed [`CalcTempBus]          temp_b1_8_6_i;
wire signed [`CalcTempBus]          temp_b1_8_7_r;
wire signed [`CalcTempBus]          temp_b1_8_7_i;
wire signed [`CalcTempBus]          temp_b1_8_8_r;
wire signed [`CalcTempBus]          temp_b1_8_8_i;
wire signed [`CalcTempBus]          temp_b2_1_1_r;
wire signed [`CalcTempBus]          temp_b2_1_1_i;
wire signed [`CalcTempBus]          temp_b2_1_2_r;
wire signed [`CalcTempBus]          temp_b2_1_2_i;
wire signed [`CalcTempBus]          temp_b2_1_3_r;
wire signed [`CalcTempBus]          temp_b2_1_3_i;
wire signed [`CalcTempBus]          temp_b2_1_4_r;
wire signed [`CalcTempBus]          temp_b2_1_4_i;
wire signed [`CalcTempBus]          temp_b2_1_5_r;
wire signed [`CalcTempBus]          temp_b2_1_5_i;
wire signed [`CalcTempBus]          temp_b2_1_6_r;
wire signed [`CalcTempBus]          temp_b2_1_6_i;
wire signed [`CalcTempBus]          temp_b2_1_7_r;
wire signed [`CalcTempBus]          temp_b2_1_7_i;
wire signed [`CalcTempBus]          temp_b2_1_8_r;
wire signed [`CalcTempBus]          temp_b2_1_8_i;
wire signed [`CalcTempBus]          temp_b2_2_1_r;
wire signed [`CalcTempBus]          temp_b2_2_1_i;
wire signed [`CalcTempBus]          temp_b2_2_2_r;
wire signed [`CalcTempBus]          temp_b2_2_2_i;
wire signed [`CalcTempBus]          temp_b2_2_3_r;
wire signed [`CalcTempBus]          temp_b2_2_3_i;
wire signed [`CalcTempBus]          temp_b2_2_4_r;
wire signed [`CalcTempBus]          temp_b2_2_4_i;
wire signed [`CalcTempBus]          temp_b2_2_5_r;
wire signed [`CalcTempBus]          temp_b2_2_5_i;
wire signed [`CalcTempBus]          temp_b2_2_6_r;
wire signed [`CalcTempBus]          temp_b2_2_6_i;
wire signed [`CalcTempBus]          temp_b2_2_7_r;
wire signed [`CalcTempBus]          temp_b2_2_7_i;
wire signed [`CalcTempBus]          temp_b2_2_8_r;
wire signed [`CalcTempBus]          temp_b2_2_8_i;
wire signed [`CalcTempBus]          temp_b2_3_1_r;
wire signed [`CalcTempBus]          temp_b2_3_1_i;
wire signed [`CalcTempBus]          temp_b2_3_2_r;
wire signed [`CalcTempBus]          temp_b2_3_2_i;
wire signed [`CalcTempBus]          temp_b2_3_3_r;
wire signed [`CalcTempBus]          temp_b2_3_3_i;
wire signed [`CalcTempBus]          temp_b2_3_4_r;
wire signed [`CalcTempBus]          temp_b2_3_4_i;
wire signed [`CalcTempBus]          temp_b2_3_5_r;
wire signed [`CalcTempBus]          temp_b2_3_5_i;
wire signed [`CalcTempBus]          temp_b2_3_6_r;
wire signed [`CalcTempBus]          temp_b2_3_6_i;
wire signed [`CalcTempBus]          temp_b2_3_7_r;
wire signed [`CalcTempBus]          temp_b2_3_7_i;
wire signed [`CalcTempBus]          temp_b2_3_8_r;
wire signed [`CalcTempBus]          temp_b2_3_8_i;
wire signed [`CalcTempBus]          temp_b2_4_1_r;
wire signed [`CalcTempBus]          temp_b2_4_1_i;
wire signed [`CalcTempBus]          temp_b2_4_2_r;
wire signed [`CalcTempBus]          temp_b2_4_2_i;
wire signed [`CalcTempBus]          temp_b2_4_3_r;
wire signed [`CalcTempBus]          temp_b2_4_3_i;
wire signed [`CalcTempBus]          temp_b2_4_4_r;
wire signed [`CalcTempBus]          temp_b2_4_4_i;
wire signed [`CalcTempBus]          temp_b2_4_5_r;
wire signed [`CalcTempBus]          temp_b2_4_5_i;
wire signed [`CalcTempBus]          temp_b2_4_6_r;
wire signed [`CalcTempBus]          temp_b2_4_6_i;
wire signed [`CalcTempBus]          temp_b2_4_7_r;
wire signed [`CalcTempBus]          temp_b2_4_7_i;
wire signed [`CalcTempBus]          temp_b2_4_8_r;
wire signed [`CalcTempBus]          temp_b2_4_8_i;
wire signed [`CalcTempBus]          temp_b2_5_1_r;
wire signed [`CalcTempBus]          temp_b2_5_1_i;
wire signed [`CalcTempBus]          temp_b2_5_2_r;
wire signed [`CalcTempBus]          temp_b2_5_2_i;
wire signed [`CalcTempBus]          temp_b2_5_3_r;
wire signed [`CalcTempBus]          temp_b2_5_3_i;
wire signed [`CalcTempBus]          temp_b2_5_4_r;
wire signed [`CalcTempBus]          temp_b2_5_4_i;
wire signed [`CalcTempBus]          temp_b2_5_5_r;
wire signed [`CalcTempBus]          temp_b2_5_5_i;
wire signed [`CalcTempBus]          temp_b2_5_6_r;
wire signed [`CalcTempBus]          temp_b2_5_6_i;
wire signed [`CalcTempBus]          temp_b2_5_7_r;
wire signed [`CalcTempBus]          temp_b2_5_7_i;
wire signed [`CalcTempBus]          temp_b2_5_8_r;
wire signed [`CalcTempBus]          temp_b2_5_8_i;
wire signed [`CalcTempBus]          temp_b2_6_1_r;
wire signed [`CalcTempBus]          temp_b2_6_1_i;
wire signed [`CalcTempBus]          temp_b2_6_2_r;
wire signed [`CalcTempBus]          temp_b2_6_2_i;
wire signed [`CalcTempBus]          temp_b2_6_3_r;
wire signed [`CalcTempBus]          temp_b2_6_3_i;
wire signed [`CalcTempBus]          temp_b2_6_4_r;
wire signed [`CalcTempBus]          temp_b2_6_4_i;
wire signed [`CalcTempBus]          temp_b2_6_5_r;
wire signed [`CalcTempBus]          temp_b2_6_5_i;
wire signed [`CalcTempBus]          temp_b2_6_6_r;
wire signed [`CalcTempBus]          temp_b2_6_6_i;
wire signed [`CalcTempBus]          temp_b2_6_7_r;
wire signed [`CalcTempBus]          temp_b2_6_7_i;
wire signed [`CalcTempBus]          temp_b2_6_8_r;
wire signed [`CalcTempBus]          temp_b2_6_8_i;
wire signed [`CalcTempBus]          temp_b2_7_1_r;
wire signed [`CalcTempBus]          temp_b2_7_1_i;
wire signed [`CalcTempBus]          temp_b2_7_2_r;
wire signed [`CalcTempBus]          temp_b2_7_2_i;
wire signed [`CalcTempBus]          temp_b2_7_3_r;
wire signed [`CalcTempBus]          temp_b2_7_3_i;
wire signed [`CalcTempBus]          temp_b2_7_4_r;
wire signed [`CalcTempBus]          temp_b2_7_4_i;
wire signed [`CalcTempBus]          temp_b2_7_5_r;
wire signed [`CalcTempBus]          temp_b2_7_5_i;
wire signed [`CalcTempBus]          temp_b2_7_6_r;
wire signed [`CalcTempBus]          temp_b2_7_6_i;
wire signed [`CalcTempBus]          temp_b2_7_7_r;
wire signed [`CalcTempBus]          temp_b2_7_7_i;
wire signed [`CalcTempBus]          temp_b2_7_8_r;
wire signed [`CalcTempBus]          temp_b2_7_8_i;
wire signed [`CalcTempBus]          temp_b2_8_1_r;
wire signed [`CalcTempBus]          temp_b2_8_1_i;
wire signed [`CalcTempBus]          temp_b2_8_2_r;
wire signed [`CalcTempBus]          temp_b2_8_2_i;
wire signed [`CalcTempBus]          temp_b2_8_3_r;
wire signed [`CalcTempBus]          temp_b2_8_3_i;
wire signed [`CalcTempBus]          temp_b2_8_4_r;
wire signed [`CalcTempBus]          temp_b2_8_4_i;
wire signed [`CalcTempBus]          temp_b2_8_5_r;
wire signed [`CalcTempBus]          temp_b2_8_5_i;
wire signed [`CalcTempBus]          temp_b2_8_6_r;
wire signed [`CalcTempBus]          temp_b2_8_6_i;
wire signed [`CalcTempBus]          temp_b2_8_7_r;
wire signed [`CalcTempBus]          temp_b2_8_7_i;
wire signed [`CalcTempBus]          temp_b2_8_8_r;
wire signed [`CalcTempBus]          temp_b2_8_8_i;
wire signed [`CalcTempBus]          temp_b3_1_1_r;
wire signed [`CalcTempBus]          temp_b3_1_1_i;
wire signed [`CalcTempBus]          temp_b3_1_2_r;
wire signed [`CalcTempBus]          temp_b3_1_2_i;
wire signed [`CalcTempBus]          temp_b3_1_3_r;
wire signed [`CalcTempBus]          temp_b3_1_3_i;
wire signed [`CalcTempBus]          temp_b3_1_4_r;
wire signed [`CalcTempBus]          temp_b3_1_4_i;
wire signed [`CalcTempBus]          temp_b3_1_5_r;
wire signed [`CalcTempBus]          temp_b3_1_5_i;
wire signed [`CalcTempBus]          temp_b3_1_6_r;
wire signed [`CalcTempBus]          temp_b3_1_6_i;
wire signed [`CalcTempBus]          temp_b3_1_7_r;
wire signed [`CalcTempBus]          temp_b3_1_7_i;
wire signed [`CalcTempBus]          temp_b3_1_8_r;
wire signed [`CalcTempBus]          temp_b3_1_8_i;
wire signed [`CalcTempBus]          temp_b3_2_1_r;
wire signed [`CalcTempBus]          temp_b3_2_1_i;
wire signed [`CalcTempBus]          temp_b3_2_2_r;
wire signed [`CalcTempBus]          temp_b3_2_2_i;
wire signed [`CalcTempBus]          temp_b3_2_3_r;
wire signed [`CalcTempBus]          temp_b3_2_3_i;
wire signed [`CalcTempBus]          temp_b3_2_4_r;
wire signed [`CalcTempBus]          temp_b3_2_4_i;
wire signed [`CalcTempBus]          temp_b3_2_5_r;
wire signed [`CalcTempBus]          temp_b3_2_5_i;
wire signed [`CalcTempBus]          temp_b3_2_6_r;
wire signed [`CalcTempBus]          temp_b3_2_6_i;
wire signed [`CalcTempBus]          temp_b3_2_7_r;
wire signed [`CalcTempBus]          temp_b3_2_7_i;
wire signed [`CalcTempBus]          temp_b3_2_8_r;
wire signed [`CalcTempBus]          temp_b3_2_8_i;
wire signed [`CalcTempBus]          temp_b3_3_1_r;
wire signed [`CalcTempBus]          temp_b3_3_1_i;
wire signed [`CalcTempBus]          temp_b3_3_2_r;
wire signed [`CalcTempBus]          temp_b3_3_2_i;
wire signed [`CalcTempBus]          temp_b3_3_3_r;
wire signed [`CalcTempBus]          temp_b3_3_3_i;
wire signed [`CalcTempBus]          temp_b3_3_4_r;
wire signed [`CalcTempBus]          temp_b3_3_4_i;
wire signed [`CalcTempBus]          temp_b3_3_5_r;
wire signed [`CalcTempBus]          temp_b3_3_5_i;
wire signed [`CalcTempBus]          temp_b3_3_6_r;
wire signed [`CalcTempBus]          temp_b3_3_6_i;
wire signed [`CalcTempBus]          temp_b3_3_7_r;
wire signed [`CalcTempBus]          temp_b3_3_7_i;
wire signed [`CalcTempBus]          temp_b3_3_8_r;
wire signed [`CalcTempBus]          temp_b3_3_8_i;
wire signed [`CalcTempBus]          temp_b3_4_1_r;
wire signed [`CalcTempBus]          temp_b3_4_1_i;
wire signed [`CalcTempBus]          temp_b3_4_2_r;
wire signed [`CalcTempBus]          temp_b3_4_2_i;
wire signed [`CalcTempBus]          temp_b3_4_3_r;
wire signed [`CalcTempBus]          temp_b3_4_3_i;
wire signed [`CalcTempBus]          temp_b3_4_4_r;
wire signed [`CalcTempBus]          temp_b3_4_4_i;
wire signed [`CalcTempBus]          temp_b3_4_5_r;
wire signed [`CalcTempBus]          temp_b3_4_5_i;
wire signed [`CalcTempBus]          temp_b3_4_6_r;
wire signed [`CalcTempBus]          temp_b3_4_6_i;
wire signed [`CalcTempBus]          temp_b3_4_7_r;
wire signed [`CalcTempBus]          temp_b3_4_7_i;
wire signed [`CalcTempBus]          temp_b3_4_8_r;
wire signed [`CalcTempBus]          temp_b3_4_8_i;
wire signed [`CalcTempBus]          temp_b3_5_1_r;
wire signed [`CalcTempBus]          temp_b3_5_1_i;
wire signed [`CalcTempBus]          temp_b3_5_2_r;
wire signed [`CalcTempBus]          temp_b3_5_2_i;
wire signed [`CalcTempBus]          temp_b3_5_3_r;
wire signed [`CalcTempBus]          temp_b3_5_3_i;
wire signed [`CalcTempBus]          temp_b3_5_4_r;
wire signed [`CalcTempBus]          temp_b3_5_4_i;
wire signed [`CalcTempBus]          temp_b3_5_5_r;
wire signed [`CalcTempBus]          temp_b3_5_5_i;
wire signed [`CalcTempBus]          temp_b3_5_6_r;
wire signed [`CalcTempBus]          temp_b3_5_6_i;
wire signed [`CalcTempBus]          temp_b3_5_7_r;
wire signed [`CalcTempBus]          temp_b3_5_7_i;
wire signed [`CalcTempBus]          temp_b3_5_8_r;
wire signed [`CalcTempBus]          temp_b3_5_8_i;
wire signed [`CalcTempBus]          temp_b3_6_1_r;
wire signed [`CalcTempBus]          temp_b3_6_1_i;
wire signed [`CalcTempBus]          temp_b3_6_2_r;
wire signed [`CalcTempBus]          temp_b3_6_2_i;
wire signed [`CalcTempBus]          temp_b3_6_3_r;
wire signed [`CalcTempBus]          temp_b3_6_3_i;
wire signed [`CalcTempBus]          temp_b3_6_4_r;
wire signed [`CalcTempBus]          temp_b3_6_4_i;
wire signed [`CalcTempBus]          temp_b3_6_5_r;
wire signed [`CalcTempBus]          temp_b3_6_5_i;
wire signed [`CalcTempBus]          temp_b3_6_6_r;
wire signed [`CalcTempBus]          temp_b3_6_6_i;
wire signed [`CalcTempBus]          temp_b3_6_7_r;
wire signed [`CalcTempBus]          temp_b3_6_7_i;
wire signed [`CalcTempBus]          temp_b3_6_8_r;
wire signed [`CalcTempBus]          temp_b3_6_8_i;
wire signed [`CalcTempBus]          temp_b3_7_1_r;
wire signed [`CalcTempBus]          temp_b3_7_1_i;
wire signed [`CalcTempBus]          temp_b3_7_2_r;
wire signed [`CalcTempBus]          temp_b3_7_2_i;
wire signed [`CalcTempBus]          temp_b3_7_3_r;
wire signed [`CalcTempBus]          temp_b3_7_3_i;
wire signed [`CalcTempBus]          temp_b3_7_4_r;
wire signed [`CalcTempBus]          temp_b3_7_4_i;
wire signed [`CalcTempBus]          temp_b3_7_5_r;
wire signed [`CalcTempBus]          temp_b3_7_5_i;
wire signed [`CalcTempBus]          temp_b3_7_6_r;
wire signed [`CalcTempBus]          temp_b3_7_6_i;
wire signed [`CalcTempBus]          temp_b3_7_7_r;
wire signed [`CalcTempBus]          temp_b3_7_7_i;
wire signed [`CalcTempBus]          temp_b3_7_8_r;
wire signed [`CalcTempBus]          temp_b3_7_8_i;
wire signed [`CalcTempBus]          temp_b3_8_1_r;
wire signed [`CalcTempBus]          temp_b3_8_1_i;
wire signed [`CalcTempBus]          temp_b3_8_2_r;
wire signed [`CalcTempBus]          temp_b3_8_2_i;
wire signed [`CalcTempBus]          temp_b3_8_3_r;
wire signed [`CalcTempBus]          temp_b3_8_3_i;
wire signed [`CalcTempBus]          temp_b3_8_4_r;
wire signed [`CalcTempBus]          temp_b3_8_4_i;
wire signed [`CalcTempBus]          temp_b3_8_5_r;
wire signed [`CalcTempBus]          temp_b3_8_5_i;
wire signed [`CalcTempBus]          temp_b3_8_6_r;
wire signed [`CalcTempBus]          temp_b3_8_6_i;
wire signed [`CalcTempBus]          temp_b3_8_7_r;
wire signed [`CalcTempBus]          temp_b3_8_7_i;
wire signed [`CalcTempBus]          temp_b3_8_8_r;
wire signed [`CalcTempBus]          temp_b3_8_8_i;

/******************port map******************/
MULT MULT1 (clk,in_1_1_r,in_1_1_i,in_1_2_r,in_1_2_i,in_2_1_r,in_2_1_i,in_2_2_r,in_2_2_i,temp_m1_1_1_r,temp_m1_1_1_i,temp_m1_1_2_r,temp_m1_1_2_i,temp_m1_2_1_r,temp_m1_2_1_i,temp_m1_2_2_r,temp_m1_2_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly1 (clk,temp_m1_1_1_r,temp_m1_1_1_i,temp_m1_1_2_r,temp_m1_1_2_i,temp_m1_2_1_r,temp_m1_2_1_i,temp_m1_2_2_r,temp_m1_2_2_i,temp_b1_1_1_r,temp_b1_1_1_i,temp_b1_1_2_r,temp_b1_1_2_i,temp_b1_2_1_r,temp_b1_2_1_i,temp_b1_2_2_r,temp_b1_2_2_i);
MULT MULT2 (clk,in_1_3_r,in_1_3_i,in_1_4_r,in_1_4_i,in_2_3_r,in_2_3_i,in_2_4_r,in_2_4_i,temp_m1_1_3_r,temp_m1_1_3_i,temp_m1_1_4_r,temp_m1_1_4_i,temp_m1_2_3_r,temp_m1_2_3_i,temp_m1_2_4_r,temp_m1_2_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly2 (clk,temp_m1_1_3_r,temp_m1_1_3_i,temp_m1_1_4_r,temp_m1_1_4_i,temp_m1_2_3_r,temp_m1_2_3_i,temp_m1_2_4_r,temp_m1_2_4_i,temp_b1_1_3_r,temp_b1_1_3_i,temp_b1_1_4_r,temp_b1_1_4_i,temp_b1_2_3_r,temp_b1_2_3_i,temp_b1_2_4_r,temp_b1_2_4_i);
MULT MULT3 (clk,in_1_5_r,in_1_5_i,in_1_6_r,in_1_6_i,in_2_5_r,in_2_5_i,in_2_6_r,in_2_6_i,temp_m1_1_5_r,temp_m1_1_5_i,temp_m1_1_6_r,temp_m1_1_6_i,temp_m1_2_5_r,temp_m1_2_5_i,temp_m1_2_6_r,temp_m1_2_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly3 (clk,temp_m1_1_5_r,temp_m1_1_5_i,temp_m1_1_6_r,temp_m1_1_6_i,temp_m1_2_5_r,temp_m1_2_5_i,temp_m1_2_6_r,temp_m1_2_6_i,temp_b1_1_5_r,temp_b1_1_5_i,temp_b1_1_6_r,temp_b1_1_6_i,temp_b1_2_5_r,temp_b1_2_5_i,temp_b1_2_6_r,temp_b1_2_6_i);
MULT MULT4 (clk,in_1_7_r,in_1_7_i,in_1_8_r,in_1_8_i,in_2_7_r,in_2_7_i,in_2_8_r,in_2_8_i,temp_m1_1_7_r,temp_m1_1_7_i,temp_m1_1_8_r,temp_m1_1_8_i,temp_m1_2_7_r,temp_m1_2_7_i,temp_m1_2_8_r,temp_m1_2_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly4 (clk,temp_m1_1_7_r,temp_m1_1_7_i,temp_m1_1_8_r,temp_m1_1_8_i,temp_m1_2_7_r,temp_m1_2_7_i,temp_m1_2_8_r,temp_m1_2_8_i,temp_b1_1_7_r,temp_b1_1_7_i,temp_b1_1_8_r,temp_b1_1_8_i,temp_b1_2_7_r,temp_b1_2_7_i,temp_b1_2_8_r,temp_b1_2_8_i);
MULT MULT5 (clk,in_3_1_r,in_3_1_i,in_3_2_r,in_3_2_i,in_4_1_r,in_4_1_i,in_4_2_r,in_4_2_i,temp_m1_3_1_r,temp_m1_3_1_i,temp_m1_3_2_r,temp_m1_3_2_i,temp_m1_4_1_r,temp_m1_4_1_i,temp_m1_4_2_r,temp_m1_4_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly5 (clk,temp_m1_3_1_r,temp_m1_3_1_i,temp_m1_3_2_r,temp_m1_3_2_i,temp_m1_4_1_r,temp_m1_4_1_i,temp_m1_4_2_r,temp_m1_4_2_i,temp_b1_3_1_r,temp_b1_3_1_i,temp_b1_3_2_r,temp_b1_3_2_i,temp_b1_4_1_r,temp_b1_4_1_i,temp_b1_4_2_r,temp_b1_4_2_i);
MULT MULT6 (clk,in_3_3_r,in_3_3_i,in_3_4_r,in_3_4_i,in_4_3_r,in_4_3_i,in_4_4_r,in_4_4_i,temp_m1_3_3_r,temp_m1_3_3_i,temp_m1_3_4_r,temp_m1_3_4_i,temp_m1_4_3_r,temp_m1_4_3_i,temp_m1_4_4_r,temp_m1_4_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly6 (clk,temp_m1_3_3_r,temp_m1_3_3_i,temp_m1_3_4_r,temp_m1_3_4_i,temp_m1_4_3_r,temp_m1_4_3_i,temp_m1_4_4_r,temp_m1_4_4_i,temp_b1_3_3_r,temp_b1_3_3_i,temp_b1_3_4_r,temp_b1_3_4_i,temp_b1_4_3_r,temp_b1_4_3_i,temp_b1_4_4_r,temp_b1_4_4_i);
MULT MULT7 (clk,in_3_5_r,in_3_5_i,in_3_6_r,in_3_6_i,in_4_5_r,in_4_5_i,in_4_6_r,in_4_6_i,temp_m1_3_5_r,temp_m1_3_5_i,temp_m1_3_6_r,temp_m1_3_6_i,temp_m1_4_5_r,temp_m1_4_5_i,temp_m1_4_6_r,temp_m1_4_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly7 (clk,temp_m1_3_5_r,temp_m1_3_5_i,temp_m1_3_6_r,temp_m1_3_6_i,temp_m1_4_5_r,temp_m1_4_5_i,temp_m1_4_6_r,temp_m1_4_6_i,temp_b1_3_5_r,temp_b1_3_5_i,temp_b1_3_6_r,temp_b1_3_6_i,temp_b1_4_5_r,temp_b1_4_5_i,temp_b1_4_6_r,temp_b1_4_6_i);
MULT MULT8 (clk,in_3_7_r,in_3_7_i,in_3_8_r,in_3_8_i,in_4_7_r,in_4_7_i,in_4_8_r,in_4_8_i,temp_m1_3_7_r,temp_m1_3_7_i,temp_m1_3_8_r,temp_m1_3_8_i,temp_m1_4_7_r,temp_m1_4_7_i,temp_m1_4_8_r,temp_m1_4_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly8 (clk,temp_m1_3_7_r,temp_m1_3_7_i,temp_m1_3_8_r,temp_m1_3_8_i,temp_m1_4_7_r,temp_m1_4_7_i,temp_m1_4_8_r,temp_m1_4_8_i,temp_b1_3_7_r,temp_b1_3_7_i,temp_b1_3_8_r,temp_b1_3_8_i,temp_b1_4_7_r,temp_b1_4_7_i,temp_b1_4_8_r,temp_b1_4_8_i);
MULT MULT9 (clk,in_5_1_r,in_5_1_i,in_5_2_r,in_5_2_i,in_6_1_r,in_6_1_i,in_6_2_r,in_6_2_i,temp_m1_5_1_r,temp_m1_5_1_i,temp_m1_5_2_r,temp_m1_5_2_i,temp_m1_6_1_r,temp_m1_6_1_i,temp_m1_6_2_r,temp_m1_6_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly9 (clk,temp_m1_5_1_r,temp_m1_5_1_i,temp_m1_5_2_r,temp_m1_5_2_i,temp_m1_6_1_r,temp_m1_6_1_i,temp_m1_6_2_r,temp_m1_6_2_i,temp_b1_5_1_r,temp_b1_5_1_i,temp_b1_5_2_r,temp_b1_5_2_i,temp_b1_6_1_r,temp_b1_6_1_i,temp_b1_6_2_r,temp_b1_6_2_i);
MULT MULT10 (clk,in_5_3_r,in_5_3_i,in_5_4_r,in_5_4_i,in_6_3_r,in_6_3_i,in_6_4_r,in_6_4_i,temp_m1_5_3_r,temp_m1_5_3_i,temp_m1_5_4_r,temp_m1_5_4_i,temp_m1_6_3_r,temp_m1_6_3_i,temp_m1_6_4_r,temp_m1_6_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly10 (clk,temp_m1_5_3_r,temp_m1_5_3_i,temp_m1_5_4_r,temp_m1_5_4_i,temp_m1_6_3_r,temp_m1_6_3_i,temp_m1_6_4_r,temp_m1_6_4_i,temp_b1_5_3_r,temp_b1_5_3_i,temp_b1_5_4_r,temp_b1_5_4_i,temp_b1_6_3_r,temp_b1_6_3_i,temp_b1_6_4_r,temp_b1_6_4_i);
MULT MULT11 (clk,in_5_5_r,in_5_5_i,in_5_6_r,in_5_6_i,in_6_5_r,in_6_5_i,in_6_6_r,in_6_6_i,temp_m1_5_5_r,temp_m1_5_5_i,temp_m1_5_6_r,temp_m1_5_6_i,temp_m1_6_5_r,temp_m1_6_5_i,temp_m1_6_6_r,temp_m1_6_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly11 (clk,temp_m1_5_5_r,temp_m1_5_5_i,temp_m1_5_6_r,temp_m1_5_6_i,temp_m1_6_5_r,temp_m1_6_5_i,temp_m1_6_6_r,temp_m1_6_6_i,temp_b1_5_5_r,temp_b1_5_5_i,temp_b1_5_6_r,temp_b1_5_6_i,temp_b1_6_5_r,temp_b1_6_5_i,temp_b1_6_6_r,temp_b1_6_6_i);
MULT MULT12 (clk,in_5_7_r,in_5_7_i,in_5_8_r,in_5_8_i,in_6_7_r,in_6_7_i,in_6_8_r,in_6_8_i,temp_m1_5_7_r,temp_m1_5_7_i,temp_m1_5_8_r,temp_m1_5_8_i,temp_m1_6_7_r,temp_m1_6_7_i,temp_m1_6_8_r,temp_m1_6_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly12 (clk,temp_m1_5_7_r,temp_m1_5_7_i,temp_m1_5_8_r,temp_m1_5_8_i,temp_m1_6_7_r,temp_m1_6_7_i,temp_m1_6_8_r,temp_m1_6_8_i,temp_b1_5_7_r,temp_b1_5_7_i,temp_b1_5_8_r,temp_b1_5_8_i,temp_b1_6_7_r,temp_b1_6_7_i,temp_b1_6_8_r,temp_b1_6_8_i);
MULT MULT13 (clk,in_7_1_r,in_7_1_i,in_7_2_r,in_7_2_i,in_8_1_r,in_8_1_i,in_8_2_r,in_8_2_i,temp_m1_7_1_r,temp_m1_7_1_i,temp_m1_7_2_r,temp_m1_7_2_i,temp_m1_8_1_r,temp_m1_8_1_i,temp_m1_8_2_r,temp_m1_8_2_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly13 (clk,temp_m1_7_1_r,temp_m1_7_1_i,temp_m1_7_2_r,temp_m1_7_2_i,temp_m1_8_1_r,temp_m1_8_1_i,temp_m1_8_2_r,temp_m1_8_2_i,temp_b1_7_1_r,temp_b1_7_1_i,temp_b1_7_2_r,temp_b1_7_2_i,temp_b1_8_1_r,temp_b1_8_1_i,temp_b1_8_2_r,temp_b1_8_2_i);
MULT MULT14 (clk,in_7_3_r,in_7_3_i,in_7_4_r,in_7_4_i,in_8_3_r,in_8_3_i,in_8_4_r,in_8_4_i,temp_m1_7_3_r,temp_m1_7_3_i,temp_m1_7_4_r,temp_m1_7_4_i,temp_m1_8_3_r,temp_m1_8_3_i,temp_m1_8_4_r,temp_m1_8_4_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly14 (clk,temp_m1_7_3_r,temp_m1_7_3_i,temp_m1_7_4_r,temp_m1_7_4_i,temp_m1_8_3_r,temp_m1_8_3_i,temp_m1_8_4_r,temp_m1_8_4_i,temp_b1_7_3_r,temp_b1_7_3_i,temp_b1_7_4_r,temp_b1_7_4_i,temp_b1_8_3_r,temp_b1_8_3_i,temp_b1_8_4_r,temp_b1_8_4_i);
MULT MULT15 (clk,in_7_5_r,in_7_5_i,in_7_6_r,in_7_6_i,in_8_5_r,in_8_5_i,in_8_6_r,in_8_6_i,temp_m1_7_5_r,temp_m1_7_5_i,temp_m1_7_6_r,temp_m1_7_6_i,temp_m1_8_5_r,temp_m1_8_5_i,temp_m1_8_6_r,temp_m1_8_6_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly15 (clk,temp_m1_7_5_r,temp_m1_7_5_i,temp_m1_7_6_r,temp_m1_7_6_i,temp_m1_8_5_r,temp_m1_8_5_i,temp_m1_8_6_r,temp_m1_8_6_i,temp_b1_7_5_r,temp_b1_7_5_i,temp_b1_7_6_r,temp_b1_7_6_i,temp_b1_8_5_r,temp_b1_8_5_i,temp_b1_8_6_r,temp_b1_8_6_i);
MULT MULT16 (clk,in_7_7_r,in_7_7_i,in_7_8_r,in_7_8_i,in_8_7_r,in_8_7_i,in_8_8_r,in_8_8_i,temp_m1_7_7_r,temp_m1_7_7_i,temp_m1_7_8_r,temp_m1_7_8_i,temp_m1_8_7_r,temp_m1_8_7_i,temp_m1_8_8_r,temp_m1_8_8_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly16 (clk,temp_m1_7_7_r,temp_m1_7_7_i,temp_m1_7_8_r,temp_m1_7_8_i,temp_m1_8_7_r,temp_m1_8_7_i,temp_m1_8_8_r,temp_m1_8_8_i,temp_b1_7_7_r,temp_b1_7_7_i,temp_b1_7_8_r,temp_b1_7_8_i,temp_b1_8_7_r,temp_b1_8_7_i,temp_b1_8_8_r,temp_b1_8_8_i);
MULT MULT17 (clk,temp_b1_1_1_r,temp_b1_1_1_i,temp_b1_1_3_r,temp_b1_1_3_i,temp_b1_3_1_r,temp_b1_3_1_i,temp_b1_3_3_r,temp_b1_3_3_i,temp_m2_1_1_r,temp_m2_1_1_i,temp_m2_1_3_r,temp_m2_1_3_i,temp_m2_3_1_r,temp_m2_3_1_i,temp_m2_3_3_r,temp_m2_3_3_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly17 (clk,temp_m2_1_1_r,temp_m2_1_1_i,temp_m2_1_3_r,temp_m2_1_3_i,temp_m2_3_1_r,temp_m2_3_1_i,temp_m2_3_3_r,temp_m2_3_3_i,temp_b2_1_1_r,temp_b2_1_1_i,temp_b2_1_3_r,temp_b2_1_3_i,temp_b2_3_1_r,temp_b2_3_1_i,temp_b2_3_3_r,temp_b2_3_3_i);
MULT MULT18 (clk,temp_b1_1_2_r,temp_b1_1_2_i,temp_b1_1_4_r,temp_b1_1_4_i,temp_b1_3_2_r,temp_b1_3_2_i,temp_b1_3_4_r,temp_b1_3_4_i,temp_m2_1_2_r,temp_m2_1_2_i,temp_m2_1_4_r,temp_m2_1_4_i,temp_m2_3_2_r,temp_m2_3_2_i,temp_m2_3_4_r,temp_m2_3_4_i,`W2_real,`W2_imag,`W0_real,`W0_imag,`W2_real,`W2_imag);
butterfly butterfly18 (clk,temp_m2_1_2_r,temp_m2_1_2_i,temp_m2_1_4_r,temp_m2_1_4_i,temp_m2_3_2_r,temp_m2_3_2_i,temp_m2_3_4_r,temp_m2_3_4_i,temp_b2_1_2_r,temp_b2_1_2_i,temp_b2_1_4_r,temp_b2_1_4_i,temp_b2_3_2_r,temp_b2_3_2_i,temp_b2_3_4_r,temp_b2_3_4_i);
MULT MULT19 (clk,temp_b1_2_1_r,temp_b1_2_1_i,temp_b1_2_3_r,temp_b1_2_3_i,temp_b1_4_1_r,temp_b1_4_1_i,temp_b1_4_3_r,temp_b1_4_3_i,temp_m2_2_1_r,temp_m2_2_1_i,temp_m2_2_3_r,temp_m2_2_3_i,temp_m2_4_1_r,temp_m2_4_1_i,temp_m2_4_3_r,temp_m2_4_3_i,`W0_real,`W0_imag,`W2_real,`W2_imag,`W2_real,`W2_imag);
butterfly butterfly19 (clk,temp_m2_2_1_r,temp_m2_2_1_i,temp_m2_2_3_r,temp_m2_2_3_i,temp_m2_4_1_r,temp_m2_4_1_i,temp_m2_4_3_r,temp_m2_4_3_i,temp_b2_2_1_r,temp_b2_2_1_i,temp_b2_2_3_r,temp_b2_2_3_i,temp_b2_4_1_r,temp_b2_4_1_i,temp_b2_4_3_r,temp_b2_4_3_i);
MULT MULT20 (clk,temp_b1_2_2_r,temp_b1_2_2_i,temp_b1_2_4_r,temp_b1_2_4_i,temp_b1_4_2_r,temp_b1_4_2_i,temp_b1_4_4_r,temp_b1_4_4_i,temp_m2_2_2_r,temp_m2_2_2_i,temp_m2_2_4_r,temp_m2_2_4_i,temp_m2_4_2_r,temp_m2_4_2_i,temp_m2_4_4_r,temp_m2_4_4_i,`W2_real,`W2_imag,`W2_real,`W2_imag,`W4_real,`W4_imag);
butterfly butterfly20 (clk,temp_m2_2_2_r,temp_m2_2_2_i,temp_m2_2_4_r,temp_m2_2_4_i,temp_m2_4_2_r,temp_m2_4_2_i,temp_m2_4_4_r,temp_m2_4_4_i,temp_b2_2_2_r,temp_b2_2_2_i,temp_b2_2_4_r,temp_b2_2_4_i,temp_b2_4_2_r,temp_b2_4_2_i,temp_b2_4_4_r,temp_b2_4_4_i);
MULT MULT21 (clk,temp_b1_1_5_r,temp_b1_1_5_i,temp_b1_1_7_r,temp_b1_1_7_i,temp_b1_3_5_r,temp_b1_3_5_i,temp_b1_3_7_r,temp_b1_3_7_i,temp_m2_1_5_r,temp_m2_1_5_i,temp_m2_1_7_r,temp_m2_1_7_i,temp_m2_3_5_r,temp_m2_3_5_i,temp_m2_3_7_r,temp_m2_3_7_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly21 (clk,temp_m2_1_5_r,temp_m2_1_5_i,temp_m2_1_7_r,temp_m2_1_7_i,temp_m2_3_5_r,temp_m2_3_5_i,temp_m2_3_7_r,temp_m2_3_7_i,temp_b2_1_5_r,temp_b2_1_5_i,temp_b2_1_7_r,temp_b2_1_7_i,temp_b2_3_5_r,temp_b2_3_5_i,temp_b2_3_7_r,temp_b2_3_7_i);
MULT MULT22 (clk,temp_b1_1_6_r,temp_b1_1_6_i,temp_b1_1_8_r,temp_b1_1_8_i,temp_b1_3_6_r,temp_b1_3_6_i,temp_b1_3_8_r,temp_b1_3_8_i,temp_m2_1_6_r,temp_m2_1_6_i,temp_m2_1_8_r,temp_m2_1_8_i,temp_m2_3_6_r,temp_m2_3_6_i,temp_m2_3_8_r,temp_m2_3_8_i,`W2_real,`W2_imag,`W0_real,`W0_imag,`W2_real,`W2_imag);
butterfly butterfly22 (clk,temp_m2_1_6_r,temp_m2_1_6_i,temp_m2_1_8_r,temp_m2_1_8_i,temp_m2_3_6_r,temp_m2_3_6_i,temp_m2_3_8_r,temp_m2_3_8_i,temp_b2_1_6_r,temp_b2_1_6_i,temp_b2_1_8_r,temp_b2_1_8_i,temp_b2_3_6_r,temp_b2_3_6_i,temp_b2_3_8_r,temp_b2_3_8_i);
MULT MULT23 (clk,temp_b1_2_5_r,temp_b1_2_5_i,temp_b1_2_7_r,temp_b1_2_7_i,temp_b1_4_5_r,temp_b1_4_5_i,temp_b1_4_7_r,temp_b1_4_7_i,temp_m2_2_5_r,temp_m2_2_5_i,temp_m2_2_7_r,temp_m2_2_7_i,temp_m2_4_5_r,temp_m2_4_5_i,temp_m2_4_7_r,temp_m2_4_7_i,`W0_real,`W0_imag,`W2_real,`W2_imag,`W2_real,`W2_imag);
butterfly butterfly23 (clk,temp_m2_2_5_r,temp_m2_2_5_i,temp_m2_2_7_r,temp_m2_2_7_i,temp_m2_4_5_r,temp_m2_4_5_i,temp_m2_4_7_r,temp_m2_4_7_i,temp_b2_2_5_r,temp_b2_2_5_i,temp_b2_2_7_r,temp_b2_2_7_i,temp_b2_4_5_r,temp_b2_4_5_i,temp_b2_4_7_r,temp_b2_4_7_i);
MULT MULT24 (clk,temp_b1_2_6_r,temp_b1_2_6_i,temp_b1_2_8_r,temp_b1_2_8_i,temp_b1_4_6_r,temp_b1_4_6_i,temp_b1_4_8_r,temp_b1_4_8_i,temp_m2_2_6_r,temp_m2_2_6_i,temp_m2_2_8_r,temp_m2_2_8_i,temp_m2_4_6_r,temp_m2_4_6_i,temp_m2_4_8_r,temp_m2_4_8_i,`W2_real,`W2_imag,`W2_real,`W2_imag,`W4_real,`W4_imag);
butterfly butterfly24 (clk,temp_m2_2_6_r,temp_m2_2_6_i,temp_m2_2_8_r,temp_m2_2_8_i,temp_m2_4_6_r,temp_m2_4_6_i,temp_m2_4_8_r,temp_m2_4_8_i,temp_b2_2_6_r,temp_b2_2_6_i,temp_b2_2_8_r,temp_b2_2_8_i,temp_b2_4_6_r,temp_b2_4_6_i,temp_b2_4_8_r,temp_b2_4_8_i);
MULT MULT25 (clk,temp_b1_5_1_r,temp_b1_5_1_i,temp_b1_5_3_r,temp_b1_5_3_i,temp_b1_7_1_r,temp_b1_7_1_i,temp_b1_7_3_r,temp_b1_7_3_i,temp_m2_5_1_r,temp_m2_5_1_i,temp_m2_5_3_r,temp_m2_5_3_i,temp_m2_7_1_r,temp_m2_7_1_i,temp_m2_7_3_r,temp_m2_7_3_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly25 (clk,temp_m2_5_1_r,temp_m2_5_1_i,temp_m2_5_3_r,temp_m2_5_3_i,temp_m2_7_1_r,temp_m2_7_1_i,temp_m2_7_3_r,temp_m2_7_3_i,temp_b2_5_1_r,temp_b2_5_1_i,temp_b2_5_3_r,temp_b2_5_3_i,temp_b2_7_1_r,temp_b2_7_1_i,temp_b2_7_3_r,temp_b2_7_3_i);
MULT MULT26 (clk,temp_b1_5_2_r,temp_b1_5_2_i,temp_b1_5_4_r,temp_b1_5_4_i,temp_b1_7_2_r,temp_b1_7_2_i,temp_b1_7_4_r,temp_b1_7_4_i,temp_m2_5_2_r,temp_m2_5_2_i,temp_m2_5_4_r,temp_m2_5_4_i,temp_m2_7_2_r,temp_m2_7_2_i,temp_m2_7_4_r,temp_m2_7_4_i,`W2_real,`W2_imag,`W0_real,`W0_imag,`W2_real,`W2_imag);
butterfly butterfly26 (clk,temp_m2_5_2_r,temp_m2_5_2_i,temp_m2_5_4_r,temp_m2_5_4_i,temp_m2_7_2_r,temp_m2_7_2_i,temp_m2_7_4_r,temp_m2_7_4_i,temp_b2_5_2_r,temp_b2_5_2_i,temp_b2_5_4_r,temp_b2_5_4_i,temp_b2_7_2_r,temp_b2_7_2_i,temp_b2_7_4_r,temp_b2_7_4_i);
MULT MULT27 (clk,temp_b1_6_1_r,temp_b1_6_1_i,temp_b1_6_3_r,temp_b1_6_3_i,temp_b1_8_1_r,temp_b1_8_1_i,temp_b1_8_3_r,temp_b1_8_3_i,temp_m2_6_1_r,temp_m2_6_1_i,temp_m2_6_3_r,temp_m2_6_3_i,temp_m2_8_1_r,temp_m2_8_1_i,temp_m2_8_3_r,temp_m2_8_3_i,`W0_real,`W0_imag,`W2_real,`W2_imag,`W2_real,`W2_imag);
butterfly butterfly27 (clk,temp_m2_6_1_r,temp_m2_6_1_i,temp_m2_6_3_r,temp_m2_6_3_i,temp_m2_8_1_r,temp_m2_8_1_i,temp_m2_8_3_r,temp_m2_8_3_i,temp_b2_6_1_r,temp_b2_6_1_i,temp_b2_6_3_r,temp_b2_6_3_i,temp_b2_8_1_r,temp_b2_8_1_i,temp_b2_8_3_r,temp_b2_8_3_i);
MULT MULT28 (clk,temp_b1_6_2_r,temp_b1_6_2_i,temp_b1_6_4_r,temp_b1_6_4_i,temp_b1_8_2_r,temp_b1_8_2_i,temp_b1_8_4_r,temp_b1_8_4_i,temp_m2_6_2_r,temp_m2_6_2_i,temp_m2_6_4_r,temp_m2_6_4_i,temp_m2_8_2_r,temp_m2_8_2_i,temp_m2_8_4_r,temp_m2_8_4_i,`W2_real,`W2_imag,`W2_real,`W2_imag,`W4_real,`W4_imag);
butterfly butterfly28 (clk,temp_m2_6_2_r,temp_m2_6_2_i,temp_m2_6_4_r,temp_m2_6_4_i,temp_m2_8_2_r,temp_m2_8_2_i,temp_m2_8_4_r,temp_m2_8_4_i,temp_b2_6_2_r,temp_b2_6_2_i,temp_b2_6_4_r,temp_b2_6_4_i,temp_b2_8_2_r,temp_b2_8_2_i,temp_b2_8_4_r,temp_b2_8_4_i);
MULT MULT29 (clk,temp_b1_5_5_r,temp_b1_5_5_i,temp_b1_5_7_r,temp_b1_5_7_i,temp_b1_7_5_r,temp_b1_7_5_i,temp_b1_7_7_r,temp_b1_7_7_i,temp_m2_5_5_r,temp_m2_5_5_i,temp_m2_5_7_r,temp_m2_5_7_i,temp_m2_7_5_r,temp_m2_7_5_i,temp_m2_7_7_r,temp_m2_7_7_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly29 (clk,temp_m2_5_5_r,temp_m2_5_5_i,temp_m2_5_7_r,temp_m2_5_7_i,temp_m2_7_5_r,temp_m2_7_5_i,temp_m2_7_7_r,temp_m2_7_7_i,temp_b2_5_5_r,temp_b2_5_5_i,temp_b2_5_7_r,temp_b2_5_7_i,temp_b2_7_5_r,temp_b2_7_5_i,temp_b2_7_7_r,temp_b2_7_7_i);
MULT MULT30 (clk,temp_b1_5_6_r,temp_b1_5_6_i,temp_b1_5_8_r,temp_b1_5_8_i,temp_b1_7_6_r,temp_b1_7_6_i,temp_b1_7_8_r,temp_b1_7_8_i,temp_m2_5_6_r,temp_m2_5_6_i,temp_m2_5_8_r,temp_m2_5_8_i,temp_m2_7_6_r,temp_m2_7_6_i,temp_m2_7_8_r,temp_m2_7_8_i,`W2_real,`W2_imag,`W0_real,`W0_imag,`W2_real,`W2_imag);
butterfly butterfly30 (clk,temp_m2_5_6_r,temp_m2_5_6_i,temp_m2_5_8_r,temp_m2_5_8_i,temp_m2_7_6_r,temp_m2_7_6_i,temp_m2_7_8_r,temp_m2_7_8_i,temp_b2_5_6_r,temp_b2_5_6_i,temp_b2_5_8_r,temp_b2_5_8_i,temp_b2_7_6_r,temp_b2_7_6_i,temp_b2_7_8_r,temp_b2_7_8_i);
MULT MULT31 (clk,temp_b1_6_5_r,temp_b1_6_5_i,temp_b1_6_7_r,temp_b1_6_7_i,temp_b1_8_5_r,temp_b1_8_5_i,temp_b1_8_7_r,temp_b1_8_7_i,temp_m2_6_5_r,temp_m2_6_5_i,temp_m2_6_7_r,temp_m2_6_7_i,temp_m2_8_5_r,temp_m2_8_5_i,temp_m2_8_7_r,temp_m2_8_7_i,`W0_real,`W0_imag,`W2_real,`W2_imag,`W2_real,`W2_imag);
butterfly butterfly31 (clk,temp_m2_6_5_r,temp_m2_6_5_i,temp_m2_6_7_r,temp_m2_6_7_i,temp_m2_8_5_r,temp_m2_8_5_i,temp_m2_8_7_r,temp_m2_8_7_i,temp_b2_6_5_r,temp_b2_6_5_i,temp_b2_6_7_r,temp_b2_6_7_i,temp_b2_8_5_r,temp_b2_8_5_i,temp_b2_8_7_r,temp_b2_8_7_i);
MULT MULT32 (clk,temp_b1_6_6_r,temp_b1_6_6_i,temp_b1_6_8_r,temp_b1_6_8_i,temp_b1_8_6_r,temp_b1_8_6_i,temp_b1_8_8_r,temp_b1_8_8_i,temp_m2_6_6_r,temp_m2_6_6_i,temp_m2_6_8_r,temp_m2_6_8_i,temp_m2_8_6_r,temp_m2_8_6_i,temp_m2_8_8_r,temp_m2_8_8_i,`W2_real,`W2_imag,`W2_real,`W2_imag,`W4_real,`W4_imag);
butterfly butterfly32 (clk,temp_m2_6_6_r,temp_m2_6_6_i,temp_m2_6_8_r,temp_m2_6_8_i,temp_m2_8_6_r,temp_m2_8_6_i,temp_m2_8_8_r,temp_m2_8_8_i,temp_b2_6_6_r,temp_b2_6_6_i,temp_b2_6_8_r,temp_b2_6_8_i,temp_b2_8_6_r,temp_b2_8_6_i,temp_b2_8_8_r,temp_b2_8_8_i);
MULT MULT33 (clk,temp_b2_1_1_r,temp_b2_1_1_i,temp_b2_1_5_r,temp_b2_1_5_i,temp_b2_5_1_r,temp_b2_5_1_i,temp_b2_5_5_r,temp_b2_5_5_i,temp_m3_1_1_r,temp_m3_1_1_i,temp_m3_1_5_r,temp_m3_1_5_i,temp_m3_5_1_r,temp_m3_5_1_i,temp_m3_5_5_r,temp_m3_5_5_i,`W0_real,`W0_imag,`W0_real,`W0_imag,`W0_real,`W0_imag);
butterfly butterfly33 (clk,temp_m3_1_1_r,temp_m3_1_1_i,temp_m3_1_5_r,temp_m3_1_5_i,temp_m3_5_1_r,temp_m3_5_1_i,temp_m3_5_5_r,temp_m3_5_5_i,temp_b3_1_1_r,temp_b3_1_1_i,temp_b3_1_5_r,temp_b3_1_5_i,temp_b3_5_1_r,temp_b3_5_1_i,temp_b3_5_5_r,temp_b3_5_5_i);
MULT MULT34 (clk,temp_b2_1_2_r,temp_b2_1_2_i,temp_b2_1_6_r,temp_b2_1_6_i,temp_b2_5_2_r,temp_b2_5_2_i,temp_b2_5_6_r,temp_b2_5_6_i,temp_m3_1_2_r,temp_m3_1_2_i,temp_m3_1_6_r,temp_m3_1_6_i,temp_m3_5_2_r,temp_m3_5_2_i,temp_m3_5_6_r,temp_m3_5_6_i,`W1_real,`W1_imag,`W0_real,`W0_imag,`W1_real,`W1_imag);
butterfly butterfly34 (clk,temp_m3_1_2_r,temp_m3_1_2_i,temp_m3_1_6_r,temp_m3_1_6_i,temp_m3_5_2_r,temp_m3_5_2_i,temp_m3_5_6_r,temp_m3_5_6_i,temp_b3_1_2_r,temp_b3_1_2_i,temp_b3_1_6_r,temp_b3_1_6_i,temp_b3_5_2_r,temp_b3_5_2_i,temp_b3_5_6_r,temp_b3_5_6_i);
MULT MULT35 (clk,temp_b2_1_3_r,temp_b2_1_3_i,temp_b2_1_7_r,temp_b2_1_7_i,temp_b2_5_3_r,temp_b2_5_3_i,temp_b2_5_7_r,temp_b2_5_7_i,temp_m3_1_3_r,temp_m3_1_3_i,temp_m3_1_7_r,temp_m3_1_7_i,temp_m3_5_3_r,temp_m3_5_3_i,temp_m3_5_7_r,temp_m3_5_7_i,`W2_real,`W2_imag,`W0_real,`W0_imag,`W2_real,`W2_imag);
butterfly butterfly35 (clk,temp_m3_1_3_r,temp_m3_1_3_i,temp_m3_1_7_r,temp_m3_1_7_i,temp_m3_5_3_r,temp_m3_5_3_i,temp_m3_5_7_r,temp_m3_5_7_i,temp_b3_1_3_r,temp_b3_1_3_i,temp_b3_1_7_r,temp_b3_1_7_i,temp_b3_5_3_r,temp_b3_5_3_i,temp_b3_5_7_r,temp_b3_5_7_i);
MULT MULT36 (clk,temp_b2_1_4_r,temp_b2_1_4_i,temp_b2_1_8_r,temp_b2_1_8_i,temp_b2_5_4_r,temp_b2_5_4_i,temp_b2_5_8_r,temp_b2_5_8_i,temp_m3_1_4_r,temp_m3_1_4_i,temp_m3_1_8_r,temp_m3_1_8_i,temp_m3_5_4_r,temp_m3_5_4_i,temp_m3_5_8_r,temp_m3_5_8_i,`W3_real,`W3_imag,`W0_real,`W0_imag,`W3_real,`W3_imag);
butterfly butterfly36 (clk,temp_m3_1_4_r,temp_m3_1_4_i,temp_m3_1_8_r,temp_m3_1_8_i,temp_m3_5_4_r,temp_m3_5_4_i,temp_m3_5_8_r,temp_m3_5_8_i,temp_b3_1_4_r,temp_b3_1_4_i,temp_b3_1_8_r,temp_b3_1_8_i,temp_b3_5_4_r,temp_b3_5_4_i,temp_b3_5_8_r,temp_b3_5_8_i);
MULT MULT37 (clk,temp_b2_2_1_r,temp_b2_2_1_i,temp_b2_2_5_r,temp_b2_2_5_i,temp_b2_6_1_r,temp_b2_6_1_i,temp_b2_6_5_r,temp_b2_6_5_i,temp_m3_2_1_r,temp_m3_2_1_i,temp_m3_2_5_r,temp_m3_2_5_i,temp_m3_6_1_r,temp_m3_6_1_i,temp_m3_6_5_r,temp_m3_6_5_i,`W0_real,`W0_imag,`W1_real,`W1_imag,`W1_real,`W1_imag);
butterfly butterfly37 (clk,temp_m3_2_1_r,temp_m3_2_1_i,temp_m3_2_5_r,temp_m3_2_5_i,temp_m3_6_1_r,temp_m3_6_1_i,temp_m3_6_5_r,temp_m3_6_5_i,temp_b3_2_1_r,temp_b3_2_1_i,temp_b3_2_5_r,temp_b3_2_5_i,temp_b3_6_1_r,temp_b3_6_1_i,temp_b3_6_5_r,temp_b3_6_5_i);
MULT MULT38 (clk,temp_b2_2_2_r,temp_b2_2_2_i,temp_b2_2_6_r,temp_b2_2_6_i,temp_b2_6_2_r,temp_b2_6_2_i,temp_b2_6_6_r,temp_b2_6_6_i,temp_m3_2_2_r,temp_m3_2_2_i,temp_m3_2_6_r,temp_m3_2_6_i,temp_m3_6_2_r,temp_m3_6_2_i,temp_m3_6_6_r,temp_m3_6_6_i,`W1_real,`W1_imag,`W1_real,`W1_imag,`W2_real,`W2_imag);
butterfly butterfly38 (clk,temp_m3_2_2_r,temp_m3_2_2_i,temp_m3_2_6_r,temp_m3_2_6_i,temp_m3_6_2_r,temp_m3_6_2_i,temp_m3_6_6_r,temp_m3_6_6_i,temp_b3_2_2_r,temp_b3_2_2_i,temp_b3_2_6_r,temp_b3_2_6_i,temp_b3_6_2_r,temp_b3_6_2_i,temp_b3_6_6_r,temp_b3_6_6_i);
MULT MULT39 (clk,temp_b2_2_3_r,temp_b2_2_3_i,temp_b2_2_7_r,temp_b2_2_7_i,temp_b2_6_3_r,temp_b2_6_3_i,temp_b2_6_7_r,temp_b2_6_7_i,temp_m3_2_3_r,temp_m3_2_3_i,temp_m3_2_7_r,temp_m3_2_7_i,temp_m3_6_3_r,temp_m3_6_3_i,temp_m3_6_7_r,temp_m3_6_7_i,`W2_real,`W2_imag,`W1_real,`W1_imag,`W3_real,`W3_imag);
butterfly butterfly39 (clk,temp_m3_2_3_r,temp_m3_2_3_i,temp_m3_2_7_r,temp_m3_2_7_i,temp_m3_6_3_r,temp_m3_6_3_i,temp_m3_6_7_r,temp_m3_6_7_i,temp_b3_2_3_r,temp_b3_2_3_i,temp_b3_2_7_r,temp_b3_2_7_i,temp_b3_6_3_r,temp_b3_6_3_i,temp_b3_6_7_r,temp_b3_6_7_i);
MULT MULT40 (clk,temp_b2_2_4_r,temp_b2_2_4_i,temp_b2_2_8_r,temp_b2_2_8_i,temp_b2_6_4_r,temp_b2_6_4_i,temp_b2_6_8_r,temp_b2_6_8_i,temp_m3_2_4_r,temp_m3_2_4_i,temp_m3_2_8_r,temp_m3_2_8_i,temp_m3_6_4_r,temp_m3_6_4_i,temp_m3_6_8_r,temp_m3_6_8_i,`W3_real,`W3_imag,`W1_real,`W1_imag,`W4_real,`W4_imag);
butterfly butterfly40 (clk,temp_m3_2_4_r,temp_m3_2_4_i,temp_m3_2_8_r,temp_m3_2_8_i,temp_m3_6_4_r,temp_m3_6_4_i,temp_m3_6_8_r,temp_m3_6_8_i,temp_b3_2_4_r,temp_b3_2_4_i,temp_b3_2_8_r,temp_b3_2_8_i,temp_b3_6_4_r,temp_b3_6_4_i,temp_b3_6_8_r,temp_b3_6_8_i);
MULT MULT41 (clk,temp_b2_3_1_r,temp_b2_3_1_i,temp_b2_3_5_r,temp_b2_3_5_i,temp_b2_7_1_r,temp_b2_7_1_i,temp_b2_7_5_r,temp_b2_7_5_i,temp_m3_3_1_r,temp_m3_3_1_i,temp_m3_3_5_r,temp_m3_3_5_i,temp_m3_7_1_r,temp_m3_7_1_i,temp_m3_7_5_r,temp_m3_7_5_i,`W0_real,`W0_imag,`W2_real,`W2_imag,`W2_real,`W2_imag);
butterfly butterfly41 (clk,temp_m3_3_1_r,temp_m3_3_1_i,temp_m3_3_5_r,temp_m3_3_5_i,temp_m3_7_1_r,temp_m3_7_1_i,temp_m3_7_5_r,temp_m3_7_5_i,temp_b3_3_1_r,temp_b3_3_1_i,temp_b3_3_5_r,temp_b3_3_5_i,temp_b3_7_1_r,temp_b3_7_1_i,temp_b3_7_5_r,temp_b3_7_5_i);
MULT MULT42 (clk,temp_b2_3_2_r,temp_b2_3_2_i,temp_b2_3_6_r,temp_b2_3_6_i,temp_b2_7_2_r,temp_b2_7_2_i,temp_b2_7_6_r,temp_b2_7_6_i,temp_m3_3_2_r,temp_m3_3_2_i,temp_m3_3_6_r,temp_m3_3_6_i,temp_m3_7_2_r,temp_m3_7_2_i,temp_m3_7_6_r,temp_m3_7_6_i,`W1_real,`W1_imag,`W2_real,`W2_imag,`W3_real,`W3_imag);
butterfly butterfly42 (clk,temp_m3_3_2_r,temp_m3_3_2_i,temp_m3_3_6_r,temp_m3_3_6_i,temp_m3_7_2_r,temp_m3_7_2_i,temp_m3_7_6_r,temp_m3_7_6_i,temp_b3_3_2_r,temp_b3_3_2_i,temp_b3_3_6_r,temp_b3_3_6_i,temp_b3_7_2_r,temp_b3_7_2_i,temp_b3_7_6_r,temp_b3_7_6_i);
MULT MULT43 (clk,temp_b2_3_3_r,temp_b2_3_3_i,temp_b2_3_7_r,temp_b2_3_7_i,temp_b2_7_3_r,temp_b2_7_3_i,temp_b2_7_7_r,temp_b2_7_7_i,temp_m3_3_3_r,temp_m3_3_3_i,temp_m3_3_7_r,temp_m3_3_7_i,temp_m3_7_3_r,temp_m3_7_3_i,temp_m3_7_7_r,temp_m3_7_7_i,`W2_real,`W2_imag,`W2_real,`W2_imag,`W4_real,`W4_imag);
butterfly butterfly43 (clk,temp_m3_3_3_r,temp_m3_3_3_i,temp_m3_3_7_r,temp_m3_3_7_i,temp_m3_7_3_r,temp_m3_7_3_i,temp_m3_7_7_r,temp_m3_7_7_i,temp_b3_3_3_r,temp_b3_3_3_i,temp_b3_3_7_r,temp_b3_3_7_i,temp_b3_7_3_r,temp_b3_7_3_i,temp_b3_7_7_r,temp_b3_7_7_i);
MULT MULT44 (clk,temp_b2_3_4_r,temp_b2_3_4_i,temp_b2_3_8_r,temp_b2_3_8_i,temp_b2_7_4_r,temp_b2_7_4_i,temp_b2_7_8_r,temp_b2_7_8_i,temp_m3_3_4_r,temp_m3_3_4_i,temp_m3_3_8_r,temp_m3_3_8_i,temp_m3_7_4_r,temp_m3_7_4_i,temp_m3_7_8_r,temp_m3_7_8_i,`W3_real,`W3_imag,`W2_real,`W2_imag,`W5_real,`W5_imag);
butterfly butterfly44 (clk,temp_m3_3_4_r,temp_m3_3_4_i,temp_m3_3_8_r,temp_m3_3_8_i,temp_m3_7_4_r,temp_m3_7_4_i,temp_m3_7_8_r,temp_m3_7_8_i,temp_b3_3_4_r,temp_b3_3_4_i,temp_b3_3_8_r,temp_b3_3_8_i,temp_b3_7_4_r,temp_b3_7_4_i,temp_b3_7_8_r,temp_b3_7_8_i);
MULT MULT45 (clk,temp_b2_4_1_r,temp_b2_4_1_i,temp_b2_4_5_r,temp_b2_4_5_i,temp_b2_8_1_r,temp_b2_8_1_i,temp_b2_8_5_r,temp_b2_8_5_i,temp_m3_4_1_r,temp_m3_4_1_i,temp_m3_4_5_r,temp_m3_4_5_i,temp_m3_8_1_r,temp_m3_8_1_i,temp_m3_8_5_r,temp_m3_8_5_i,`W0_real,`W0_imag,`W3_real,`W3_imag,`W3_real,`W3_imag);
butterfly butterfly45 (clk,temp_m3_4_1_r,temp_m3_4_1_i,temp_m3_4_5_r,temp_m3_4_5_i,temp_m3_8_1_r,temp_m3_8_1_i,temp_m3_8_5_r,temp_m3_8_5_i,temp_b3_4_1_r,temp_b3_4_1_i,temp_b3_4_5_r,temp_b3_4_5_i,temp_b3_8_1_r,temp_b3_8_1_i,temp_b3_8_5_r,temp_b3_8_5_i);
MULT MULT46 (clk,temp_b2_4_2_r,temp_b2_4_2_i,temp_b2_4_6_r,temp_b2_4_6_i,temp_b2_8_2_r,temp_b2_8_2_i,temp_b2_8_6_r,temp_b2_8_6_i,temp_m3_4_2_r,temp_m3_4_2_i,temp_m3_4_6_r,temp_m3_4_6_i,temp_m3_8_2_r,temp_m3_8_2_i,temp_m3_8_6_r,temp_m3_8_6_i,`W1_real,`W1_imag,`W3_real,`W3_imag,`W4_real,`W4_imag);
butterfly butterfly46 (clk,temp_m3_4_2_r,temp_m3_4_2_i,temp_m3_4_6_r,temp_m3_4_6_i,temp_m3_8_2_r,temp_m3_8_2_i,temp_m3_8_6_r,temp_m3_8_6_i,temp_b3_4_2_r,temp_b3_4_2_i,temp_b3_4_6_r,temp_b3_4_6_i,temp_b3_8_2_r,temp_b3_8_2_i,temp_b3_8_6_r,temp_b3_8_6_i);
MULT MULT47 (clk,temp_b2_4_3_r,temp_b2_4_3_i,temp_b2_4_7_r,temp_b2_4_7_i,temp_b2_8_3_r,temp_b2_8_3_i,temp_b2_8_7_r,temp_b2_8_7_i,temp_m3_4_3_r,temp_m3_4_3_i,temp_m3_4_7_r,temp_m3_4_7_i,temp_m3_8_3_r,temp_m3_8_3_i,temp_m3_8_7_r,temp_m3_8_7_i,`W2_real,`W2_imag,`W3_real,`W3_imag,`W5_real,`W5_imag);
butterfly butterfly47 (clk,temp_m3_4_3_r,temp_m3_4_3_i,temp_m3_4_7_r,temp_m3_4_7_i,temp_m3_8_3_r,temp_m3_8_3_i,temp_m3_8_7_r,temp_m3_8_7_i,temp_b3_4_3_r,temp_b3_4_3_i,temp_b3_4_7_r,temp_b3_4_7_i,temp_b3_8_3_r,temp_b3_8_3_i,temp_b3_8_7_r,temp_b3_8_7_i);
MULT MULT48 (clk,temp_b2_4_4_r,temp_b2_4_4_i,temp_b2_4_8_r,temp_b2_4_8_i,temp_b2_8_4_r,temp_b2_8_4_i,temp_b2_8_8_r,temp_b2_8_8_i,temp_m3_4_4_r,temp_m3_4_4_i,temp_m3_4_8_r,temp_m3_4_8_i,temp_m3_8_4_r,temp_m3_8_4_i,temp_m3_8_8_r,temp_m3_8_8_i,`W3_real,`W3_imag,`W3_real,`W3_imag,`W6_real,`W6_imag);
butterfly butterfly48 (clk,temp_m3_4_4_r,temp_m3_4_4_i,temp_m3_4_8_r,temp_m3_4_8_i,temp_m3_8_4_r,temp_m3_8_4_i,temp_m3_8_8_r,temp_m3_8_8_i,temp_b3_4_4_r,temp_b3_4_4_i,temp_b3_4_8_r,temp_b3_4_8_i,temp_b3_8_4_r,temp_b3_8_4_i,temp_b3_8_8_r,temp_b3_8_8_i);

assign out_1_1_r = temp_b3_1_1_r;
assign out_1_1_i = temp_b3_1_1_i;
assign out_1_2_r = temp_b3_1_2_r;
assign out_1_2_i = temp_b3_1_2_i;
assign out_1_3_r = temp_b3_1_3_r;
assign out_1_3_i = temp_b3_1_3_i;
assign out_1_4_r = temp_b3_1_4_r;
assign out_1_4_i = temp_b3_1_4_i;
assign out_1_5_r = temp_b3_1_5_r;
assign out_1_5_i = temp_b3_1_5_i;
assign out_1_6_r = temp_b3_1_6_r;
assign out_1_6_i = temp_b3_1_6_i;
assign out_1_7_r = temp_b3_1_7_r;
assign out_1_7_i = temp_b3_1_7_i;
assign out_1_8_r = temp_b3_1_8_r;
assign out_1_8_i = temp_b3_1_8_i;
assign out_2_1_r = temp_b3_2_1_r;
assign out_2_1_i = temp_b3_2_1_i;
assign out_2_2_r = temp_b3_2_2_r;
assign out_2_2_i = temp_b3_2_2_i;
assign out_2_3_r = temp_b3_2_3_r;
assign out_2_3_i = temp_b3_2_3_i;
assign out_2_4_r = temp_b3_2_4_r;
assign out_2_4_i = temp_b3_2_4_i;
assign out_2_5_r = temp_b3_2_5_r;
assign out_2_5_i = temp_b3_2_5_i;
assign out_2_6_r = temp_b3_2_6_r;
assign out_2_6_i = temp_b3_2_6_i;
assign out_2_7_r = temp_b3_2_7_r;
assign out_2_7_i = temp_b3_2_7_i;
assign out_2_8_r = temp_b3_2_8_r;
assign out_2_8_i = temp_b3_2_8_i;
assign out_3_1_r = temp_b3_3_1_r;
assign out_3_1_i = temp_b3_3_1_i;
assign out_3_2_r = temp_b3_3_2_r;
assign out_3_2_i = temp_b3_3_2_i;
assign out_3_3_r = temp_b3_3_3_r;
assign out_3_3_i = temp_b3_3_3_i;
assign out_3_4_r = temp_b3_3_4_r;
assign out_3_4_i = temp_b3_3_4_i;
assign out_3_5_r = temp_b3_3_5_r;
assign out_3_5_i = temp_b3_3_5_i;
assign out_3_6_r = temp_b3_3_6_r;
assign out_3_6_i = temp_b3_3_6_i;
assign out_3_7_r = temp_b3_3_7_r;
assign out_3_7_i = temp_b3_3_7_i;
assign out_3_8_r = temp_b3_3_8_r;
assign out_3_8_i = temp_b3_3_8_i;
assign out_4_1_r = temp_b3_4_1_r;
assign out_4_1_i = temp_b3_4_1_i;
assign out_4_2_r = temp_b3_4_2_r;
assign out_4_2_i = temp_b3_4_2_i;
assign out_4_3_r = temp_b3_4_3_r;
assign out_4_3_i = temp_b3_4_3_i;
assign out_4_4_r = temp_b3_4_4_r;
assign out_4_4_i = temp_b3_4_4_i;
assign out_4_5_r = temp_b3_4_5_r;
assign out_4_5_i = temp_b3_4_5_i;
assign out_4_6_r = temp_b3_4_6_r;
assign out_4_6_i = temp_b3_4_6_i;
assign out_4_7_r = temp_b3_4_7_r;
assign out_4_7_i = temp_b3_4_7_i;
assign out_4_8_r = temp_b3_4_8_r;
assign out_4_8_i = temp_b3_4_8_i;
assign out_5_1_r = temp_b3_5_1_r;
assign out_5_1_i = temp_b3_5_1_i;
assign out_5_2_r = temp_b3_5_2_r;
assign out_5_2_i = temp_b3_5_2_i;
assign out_5_3_r = temp_b3_5_3_r;
assign out_5_3_i = temp_b3_5_3_i;
assign out_5_4_r = temp_b3_5_4_r;
assign out_5_4_i = temp_b3_5_4_i;
assign out_5_5_r = temp_b3_5_5_r;
assign out_5_5_i = temp_b3_5_5_i;
assign out_5_6_r = temp_b3_5_6_r;
assign out_5_6_i = temp_b3_5_6_i;
assign out_5_7_r = temp_b3_5_7_r;
assign out_5_7_i = temp_b3_5_7_i;
assign out_5_8_r = temp_b3_5_8_r;
assign out_5_8_i = temp_b3_5_8_i;
assign out_6_1_r = temp_b3_6_1_r;
assign out_6_1_i = temp_b3_6_1_i;
assign out_6_2_r = temp_b3_6_2_r;
assign out_6_2_i = temp_b3_6_2_i;
assign out_6_3_r = temp_b3_6_3_r;
assign out_6_3_i = temp_b3_6_3_i;
assign out_6_4_r = temp_b3_6_4_r;
assign out_6_4_i = temp_b3_6_4_i;
assign out_6_5_r = temp_b3_6_5_r;
assign out_6_5_i = temp_b3_6_5_i;
assign out_6_6_r = temp_b3_6_6_r;
assign out_6_6_i = temp_b3_6_6_i;
assign out_6_7_r = temp_b3_6_7_r;
assign out_6_7_i = temp_b3_6_7_i;
assign out_6_8_r = temp_b3_6_8_r;
assign out_6_8_i = temp_b3_6_8_i;
assign out_7_1_r = temp_b3_7_1_r;
assign out_7_1_i = temp_b3_7_1_i;
assign out_7_2_r = temp_b3_7_2_r;
assign out_7_2_i = temp_b3_7_2_i;
assign out_7_3_r = temp_b3_7_3_r;
assign out_7_3_i = temp_b3_7_3_i;
assign out_7_4_r = temp_b3_7_4_r;
assign out_7_4_i = temp_b3_7_4_i;
assign out_7_5_r = temp_b3_7_5_r;
assign out_7_5_i = temp_b3_7_5_i;
assign out_7_6_r = temp_b3_7_6_r;
assign out_7_6_i = temp_b3_7_6_i;
assign out_7_7_r = temp_b3_7_7_r;
assign out_7_7_i = temp_b3_7_7_i;
assign out_7_8_r = temp_b3_7_8_r;
assign out_7_8_i = temp_b3_7_8_i;
assign out_8_1_r = temp_b3_8_1_r;
assign out_8_1_i = temp_b3_8_1_i;
assign out_8_2_r = temp_b3_8_2_r;
assign out_8_2_i = temp_b3_8_2_i;
assign out_8_3_r = temp_b3_8_3_r;
assign out_8_3_i = temp_b3_8_3_i;
assign out_8_4_r = temp_b3_8_4_r;
assign out_8_4_i = temp_b3_8_4_i;
assign out_8_5_r = temp_b3_8_5_r;
assign out_8_5_i = temp_b3_8_5_i;
assign out_8_6_r = temp_b3_8_6_r;
assign out_8_6_i = temp_b3_8_6_i;
assign out_8_7_r = temp_b3_8_7_r;
assign out_8_7_i = temp_b3_8_7_i;
assign out_8_8_r = temp_b3_8_8_r;
assign out_8_8_i = temp_b3_8_8_i;



endmodule
